module top
#( parameter param51 = ((((8'ha7) >> {((8'hb4) ? (8'ha0) : (8'hac))}) ? (~(((8'h9e) ? (7'h40) : (8'ha5)) ? {(8'hbd)} : ((8'had) & (8'hbe)))) : ((((8'had) >>> (8'hb4)) ? (|(7'h40)) : ((8'hae) ? (8'hba) : (7'h41))) <= (((8'h9d) >= (8'hb8)) ? ((8'hb9) ? (8'ha8) : (8'hb2)) : (~^(8'ha7))))) <<< (((((8'ha9) && (7'h44)) | ((8'hbc) ? (8'h9e) : (8'ha6))) ? (~^(~|(8'ha7))) : (~^(!(8'h9e)))) & ((((8'hb1) ? (8'had) : (8'haf)) ? (~&(8'h9d)) : ((8'hbf) ~^ (8'ha0))) ? {{(8'hae)}, (~(8'hb0))} : (!(|(8'ha7))))))
, parameter param52 = ((({{param51, param51}} ? ((param51 ? param51 : param51) ? (7'h40) : (param51 ^ param51)) : {(param51 ? (8'ha3) : param51)}) | param51) ? param51 : (((param51 > param51) <= ((param51 ? param51 : param51) * param51)) && (((~^param51) && (|param51)) ? ((param51 ? param51 : (8'h9d)) ? ((8'hae) ? param51 : param51) : (^(8'hbd))) : ((~param51) > {param51})))) )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h251):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire3;
  input wire signed [(4'he):(1'h0)] wire2;
  input wire [(3'h5):(1'h0)] wire1;
  input wire signed [(4'hd):(1'h0)] wire0;
  wire signed [(4'hf):(1'h0)] wire50;
  wire signed [(3'h4):(1'h0)] wire49;
  reg [(4'hf):(1'h0)] reg48 = (1'h0);
  reg [(3'h7):(1'h0)] reg47 = (1'h0);
  reg [(2'h2):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg45 = (1'h0);
  reg [(4'h8):(1'h0)] reg44 = (1'h0);
  reg [(5'h10):(1'h0)] reg43 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar42 = (1'h0);
  reg [(5'h10):(1'h0)] reg41 = (1'h0);
  reg [(2'h2):(1'h0)] reg40 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar39 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar38 = (1'h0);
  wire [(4'hb):(1'h0)] wire37;
  wire signed [(4'h9):(1'h0)] wire36;
  wire signed [(5'h13):(1'h0)] wire35;
  wire signed [(4'hd):(1'h0)] wire34;
  wire signed [(5'h14):(1'h0)] wire33;
  reg signed [(5'h15):(1'h0)] reg32 = (1'h0);
  reg [(4'hf):(1'h0)] reg31 = (1'h0);
  reg [(3'h4):(1'h0)] reg30 = (1'h0);
  reg [(2'h3):(1'h0)] reg29 = (1'h0);
  reg [(4'hb):(1'h0)] reg28 = (1'h0);
  reg [(5'h13):(1'h0)] forvar27 = (1'h0);
  reg [(5'h13):(1'h0)] reg26 = (1'h0);
  reg [(4'hf):(1'h0)] reg25 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar24 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg22 = (1'h0);
  reg [(4'h9):(1'h0)] reg21 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg18 = (1'h0);
  reg [(4'hc):(1'h0)] forvar17 = (1'h0);
  reg [(5'h14):(1'h0)] reg16 = (1'h0);
  reg [(5'h12):(1'h0)] reg15 = (1'h0);
  reg [(2'h2):(1'h0)] forvar14 = (1'h0);
  wire [(5'h15):(1'h0)] wire13;
  wire [(4'h9):(1'h0)] wire12;
  reg [(5'h14):(1'h0)] reg11 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg10 = (1'h0);
  reg [(5'h10):(1'h0)] reg9 = (1'h0);
  reg [(3'h7):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar7 = (1'h0);
  reg [(4'hc):(1'h0)] reg6 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire5;
  wire [(4'h9):(1'h0)] wire4;
  assign y = {wire50,
                 wire49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 forvar42,
                 reg41,
                 reg40,
                 forvar39,
                 forvar38,
                 wire37,
                 wire36,
                 wire35,
                 wire34,
                 wire33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 forvar27,
                 reg26,
                 reg25,
                 forvar24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 forvar17,
                 reg16,
                 reg15,
                 forvar14,
                 wire13,
                 wire12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 forvar7,
                 reg6,
                 wire5,
                 wire4,
                 (1'h0)};
  assign wire4 = ($unsigned("Czv8L3zaGIg4x2zEPNBr") ?
                     wire0[(1'h0):(1'h0)] : $signed(wire2[(4'he):(1'h1)]));
  assign wire5 = $signed(("" << $unsigned({$unsigned(wire3),
                     wire2[(4'ha):(2'h3)]})));
  always
    @(posedge clk) begin
      reg6 = wire3;
      for (forvar7 = (1'h0); (forvar7 < (2'h3)); forvar7 = (forvar7 + (1'h1)))
        begin
          reg8 <= ($signed(reg6[(4'hc):(1'h1)]) ?
              ((8'had) * ($unsigned((~wire4)) != ("zPEoMXsk4ODoAyRslgO7" ?
                  "Zo3AOT" : $unsigned(wire4)))) : "TfEPHpU3esMhrdk");
          reg9 <= $signed($signed(reg8));
        end
      reg10 <= ((8'hbb) ? ("C" ~^ "") : forvar7);
      reg11 <= (8'hae);
    end
  assign wire12 = $signed("LOoZs8bfFCVV");
  assign wire13 = wire0[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      for (forvar14 = (1'h0); (forvar14 < (2'h3)); forvar14 = (forvar14 + (1'h1)))
        begin
          reg15 <= ((reg10 ?
              ({(wire5 ?
                      (8'hbb) : wire12)} & $signed(wire5)) : "PNMarhdCJxVd") < $unsigned(({reg11} ?
              (wire4[(3'h5):(2'h2)] == ((8'hbf) || wire12)) : wire13)));
          reg16 <= wire2;
          for (forvar17 = (1'h0); (forvar17 < (2'h3)); forvar17 = (forvar17 + (1'h1)))
            begin
              reg18 <= "2Fmbs";
              reg19 <= wire0;
            end
          reg20 <= ($unsigned($unsigned(((~^(8'hb2)) ?
                  $unsigned((8'hb1)) : $signed(reg10)))) ?
              {($signed(wire12) ?
                      $signed(reg6[(4'hb):(4'h8)]) : ((^~reg18) ?
                          "fdlqOLrkoudvAYVlQ" : $signed(wire1)))} : "P0Xbqay9zO6");
        end
      reg21 <= "JgW0cc5WJgxRLV6C";
      reg22 = "g1OaX9tnLQoQTv4";
      reg23 <= (!(8'hbc));
      for (forvar24 = (1'h0); (forvar24 < (3'h4)); forvar24 = (forvar24 + (1'h1)))
        begin
          reg25 <= $signed(("HB2HY5a" <<< "wf6Ar1Oaen3"));
          reg26 = {wire4};
        end
    end
  always
    @(posedge clk) begin
      for (forvar27 = (1'h0); (forvar27 < (2'h3)); forvar27 = (forvar27 + (1'h1)))
        begin
          reg28 = reg9[(4'h8):(1'h1)];
          reg29 <= (|(~^(-reg21)));
          reg30 <= wire13;
          reg31 <= $unsigned(($signed(wire3) << $unsigned((8'ha0))));
          reg32 <= (((wire0[(3'h5):(1'h0)] >>> ((^~wire4) < reg11)) ?
                  (wire13[(5'h12):(3'h5)] ?
                      reg21[(2'h2):(2'h2)] : $unsigned((wire5 ^~ reg6))) : {{reg22[(4'h9):(4'h8)]}}) ?
              (~^$signed((!((8'hb6) ?
                  wire5 : reg26)))) : {(~&$signed("sSRrTk"))});
        end
    end
  assign wire33 = $signed("Yk07WF7KSC1E3");
  assign wire34 = (($unsigned("OYOIzn0lS3ulkI2") ?
                      $unsigned({forvar14}) : "wess5DC4aUM") << wire5);
  assign wire35 = $unsigned((!$unsigned((8'hb3))));
  assign wire36 = {wire5};
  assign wire37 = (($signed($signed((|reg21))) && (-"G5Cnk3dvpzAiiI2mLcWP")) * (reg32 ?
                      ({$signed(reg16),
                          $signed((8'had))} < ($unsigned(forvar17) ?
                          $signed(forvar24) : (reg10 ?
                              reg25 : wire3))) : ("TPONpGhpfFCbEYv0PcS" ?
                          forvar14 : (8'hae))));
  always
    @(posedge clk) begin
      for (forvar38 = (1'h0); (forvar38 < (1'h1)); forvar38 = (forvar38 + (1'h1)))
        begin
          for (forvar39 = (1'h0); (forvar39 < (1'h0)); forvar39 = (forvar39 + (1'h1)))
            begin
              reg40 = ($signed(reg26) ? (!"G9FPR") : (!wire0[(4'h9):(3'h4)]));
            end
          reg41 = (forvar14[(1'h0):(1'h0)] ? "5Xx4aYtdhxACkWaJD" : "FNnd1O0V");
          for (forvar42 = (1'h0); (forvar42 < (3'h4)); forvar42 = (forvar42 + (1'h1)))
            begin
              reg43 <= reg28;
              reg44 <= (~|{reg6});
              reg45 <= (("" ?
                  "tRO1Rqku9iU" : ((reg31[(2'h3):(1'h1)] ?
                          (8'ha2) : $unsigned(reg22)) ?
                      $unsigned((wire2 ?
                          reg25 : reg9)) : {$unsigned(reg26)})) & $signed("OP6Jy"));
            end
          reg46 = $signed(("KWL" ?
              ("MfRIsTFAChr7JAd00ZW" + reg15) : $signed($signed(wire0[(3'h4):(3'h4)]))));
        end
      reg47 <= "shZhtLoIdrMyPPz0";
      reg48 <= {"gZZ",
          (forvar38 ? wire0[(1'h0):(1'h0)] : wire37[(4'hb):(3'h4)])};
    end
  assign wire49 = $signed((forvar27[(4'hf):(4'ha)] * (wire33 * {(wire12 + wire12),
                      ""})));
  assign wire50 = ((("FPvfxQeMDdaJfP3ru" <<< reg8[(3'h4):(1'h1)]) ~^ {wire49}) > wire0);
endmodule