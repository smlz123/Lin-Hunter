(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param283 = {{{({(8'hb9), (7'h43)} ? ((8'hb4) ? (8'h9f) : (8'hb5)) : ((8'ha6) ? (8'ha0) : (8'ha9))), (8'hbc)}, ((((7'h41) ? (7'h40) : (8'hba)) + ((8'hbd) || (8'hac))) ? (-((8'h9d) ? (8'ha0) : (8'h9c))) : ({(8'ha9), (8'hbe)} >>> {(7'h43)}))}, (|((^~((8'hb4) ? (8'ha9) : (8'h9f))) ? ((8'ha5) ? ((8'h9d) >>> (8'haf)) : ((8'had) >= (7'h42))) : (!((8'ha9) ? (8'haa) : (8'h9e)))))}
, parameter param284 = param283 )
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h3d9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire0;
  input wire [(4'ha):(1'h0)] wire1;
  input wire [(3'h6):(1'h0)] wire2;
  input wire [(4'hf):(1'h0)] wire3;
  reg [(3'h6):(1'h0)] reg4 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg6 = (1'h0);
  reg [(5'h15):(1'h0)] forvar7 = (1'h0);
  reg signed [(4'he):(1'h0)] reg8 = (1'h0);
  reg [(3'h5):(1'h0)] reg9 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg11 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg12 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg13 = (1'h0);
  reg [(5'h15):(1'h0)] reg14 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire15;
  wire signed [(3'h5):(1'h0)] wire16;
  reg signed [(4'hd):(1'h0)] reg17 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg18 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg19 = (1'h0);
  reg [(5'h14):(1'h0)] reg20 = (1'h0);
  reg [(4'hd):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg22 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg23 = (1'h0);
  reg [(5'h14):(1'h0)] reg24 = (1'h0);
  reg [(5'h11):(1'h0)] reg25 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg26 = (1'h0);
  reg [(5'h15):(1'h0)] reg27 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar28 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg29 = (1'h0);
  reg [(5'h10):(1'h0)] reg30 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg31 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire32;
  reg signed [(4'hf):(1'h0)] reg33 = (1'h0);
  reg [(5'h15):(1'h0)] reg34 = (1'h0);
  reg [(3'h7):(1'h0)] reg35 = (1'h0);
  wire [(5'h13):(1'h0)] wire107;
  reg [(5'h15):(1'h0)] reg109 = (1'h0);
  reg [(5'h12):(1'h0)] reg110 = (1'h0);
  reg signed [(4'he):(1'h0)] reg111 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar112 = (1'h0);
  reg [(5'h14):(1'h0)] forvar113 = (1'h0);
  reg [(5'h10):(1'h0)] reg114 = (1'h0);
  reg [(5'h12):(1'h0)] reg115 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg116 = (1'h0);
  reg [(5'h14):(1'h0)] reg117 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg118 = (1'h0);
  reg [(5'h14):(1'h0)] reg119 = (1'h0);
  reg signed [(4'he):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar121 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg122 = (1'h0);
  reg [(5'h10):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg124 = (1'h0);
  wire [(5'h13):(1'h0)] wire125;
  wire [(3'h4):(1'h0)] wire230;
  reg [(3'h7):(1'h0)] forvar232 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar233 = (1'h0);
  reg [(4'he):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg235 = (1'h0);
  reg [(4'ha):(1'h0)] reg236 = (1'h0);
  reg [(3'h7):(1'h0)] reg237 = (1'h0);
  reg [(5'h12):(1'h0)] forvar238 = (1'h0);
  reg [(5'h12):(1'h0)] forvar239 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg240 = (1'h0);
  reg [(5'h13):(1'h0)] reg241 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg242 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg243 = (1'h0);
  reg signed [(4'he):(1'h0)] reg244 = (1'h0);
  reg [(2'h3):(1'h0)] reg245 = (1'h0);
  reg [(3'h4):(1'h0)] reg246 = (1'h0);
  reg [(4'h8):(1'h0)] reg247 = (1'h0);
  reg [(4'ha):(1'h0)] reg248 = (1'h0);
  reg [(5'h14):(1'h0)] reg249 = (1'h0);
  reg [(4'hf):(1'h0)] forvar250 = (1'h0);
  reg [(3'h4):(1'h0)] reg251 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg252 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire253;
  wire signed [(5'h11):(1'h0)] wire281;
  assign y = {reg4,
                 forvar5,
                 reg6,
                 forvar7,
                 reg8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 wire15,
                 wire16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 forvar28,
                 reg29,
                 reg30,
                 reg31,
                 wire32,
                 reg33,
                 reg34,
                 reg35,
                 wire107,
                 reg109,
                 reg110,
                 reg111,
                 forvar112,
                 forvar113,
                 reg114,
                 reg115,
                 reg116,
                 reg117,
                 reg118,
                 reg119,
                 reg120,
                 forvar121,
                 reg122,
                 reg123,
                 reg124,
                 wire125,
                 wire230,
                 forvar232,
                 forvar233,
                 reg234,
                 reg235,
                 reg236,
                 reg237,
                 forvar238,
                 forvar239,
                 reg240,
                 reg241,
                 reg242,
                 reg243,
                 reg244,
                 reg245,
                 reg246,
                 reg247,
                 reg248,
                 reg249,
                 forvar250,
                 reg251,
                 reg252,
                 wire253,
                 wire281,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg4 = (!("tCi" ?
          $unsigned((((8'hb7) ?
              wire0 : wire1) - {wire1})) : $unsigned((~$unsigned(wire1)))));
      for (forvar5 = (1'h0); (forvar5 < (1'h1)); forvar5 = (forvar5 + (1'h1)))
        begin
          reg6 <= forvar5[(3'h7):(2'h2)];
        end
      for (forvar7 = (1'h0); (forvar7 < (1'h0)); forvar7 = (forvar7 + (1'h1)))
        begin
          reg8 = "w6RhC";
          reg9 = (forvar7 > ($unsigned((+(^wire3))) | $unsigned($signed("JteDHtn0Wic"))));
          reg10 <= wire0;
          reg11 = ($unsigned({reg9[(3'h4):(1'h0)],
              ($unsigned((8'ha2)) ?
                  wire2[(3'h6):(2'h3)] : $unsigned(reg6))}) << ($unsigned(reg9[(1'h0):(1'h0)]) < {(wire1[(3'h6):(2'h2)] ?
                  $unsigned(forvar7) : {wire1})}));
        end
    end
  always
    @(posedge clk) begin
      reg12 <= $signed(forvar5);
      reg13 <= reg11[(1'h1):(1'h1)];
      reg14 <= {(wire3[(4'hd):(4'hb)] && ({(~^reg12), {reg11, wire0}} ?
              $unsigned((forvar5 >>> forvar7)) : "MV5KF6")),
          reg6};
    end
  assign wire15 = "k61tlYg";
  assign wire16 = $signed((wire15 ?
                      (~&forvar7[(5'h12):(5'h10)]) : $unsigned(wire2[(3'h6):(3'h4)])));
  always
    @(posedge clk) begin
      reg17 = "u";
      reg18 = reg9[(2'h3):(2'h2)];
      reg19 <= (reg10[(4'he):(4'h9)] == reg12);
    end
  always
    @(posedge clk) begin
      reg20 <= ((8'h9d) ?
          "T33dFJbLNBECd2w" : ($signed(($unsigned(reg18) * (+reg18))) + reg18));
    end
  always
    @(posedge clk) begin
      reg21 <= (~|reg14[(3'h4):(3'h4)]);
      reg22 <= (~^"QsqBZ9m0pcUgi9wR9R");
      reg23 <= $unsigned({(reg17 * (reg21 && (~^reg21))), "qQcmi9"});
      reg24 <= (wire15[(5'h10):(3'h4)] ?
          ("P2C" ^~ ((-(reg13 * reg13)) ?
              (-(wire0 ? reg14 : (8'h9c))) : ((reg22 ? forvar5 : wire2) ?
                  (reg17 & reg21) : reg13))) : "IaaXEkx802T");
      reg25 = ("Q5tEQB9RzssCFVKiRzqv" ? reg18 : reg19[(4'hb):(3'h4)]);
    end
  always
    @(posedge clk) begin
      reg26 <= reg17;
      reg27 <= reg23;
      for (forvar28 = (1'h0); (forvar28 < (1'h1)); forvar28 = (forvar28 + (1'h1)))
        begin
          reg29 = ((|reg21[(3'h5):(1'h1)]) ?
              $signed(({"rgeZo"} ?
                  ((wire1 > (8'hb7)) > reg19) : "dSk1")) : (($signed($signed(reg17)) != "NF") || ("y7Xw" ?
                  (~|"4b5Eh") : (reg17[(4'hd):(1'h1)] <= {reg10}))));
        end
      reg30 = $signed({(wire16[(2'h2):(2'h2)] * "qok")});
      reg31 <= reg17;
    end
  assign wire32 = ((^~reg8[(4'he):(3'h4)]) ?
                      $unsigned((~|reg31[(3'h7):(3'h5)])) : $signed((((reg29 ^ wire1) < (reg22 != wire3)) & reg25)));
  always
    @(posedge clk) begin
      reg33 = ((^~(((wire16 < (8'ha3)) > $unsigned(reg10)) >>> $unsigned($unsigned((8'hb1))))) ^ reg4);
      reg34 <= reg17[(4'hc):(3'h6)];
      reg35 <= (($signed(reg17[(4'h9):(3'h4)]) > (($signed(reg29) ?
          reg23 : (reg21 ^~ reg4)) ^~ $unsigned(wire15[(5'h14):(4'h9)]))) >>> "FqnlmQeHlueesYfi1");
    end
  module36 modinst108 (wire107, clk, reg29, wire32, reg6, reg13);
  always
    @(posedge clk) begin
      reg109 = reg24;
      reg110 <= $signed(((8'h9c) ? reg19 : {(~(wire15 ? reg34 : reg25))}));
      reg111 = (reg17 - $unsigned((~&(|$signed(reg4)))));
      for (forvar112 = (1'h0); (forvar112 < (2'h2)); forvar112 = (forvar112 + (1'h1)))
        begin
          for (forvar113 = (1'h0); (forvar113 < (3'h4)); forvar113 = (forvar113 + (1'h1)))
            begin
              reg114 <= "BGZhoV";
              reg115 <= $unsigned(($unsigned($signed((reg14 || (8'hb3)))) * reg8));
              reg116 <= reg6;
              reg117 <= {$unsigned({reg19[(2'h3):(1'h1)]}), (^~wire1)};
            end
          reg118 = "p188W9UYx4VlEufvw";
          reg119 <= reg19[(3'h5):(2'h3)];
          reg120 <= ((reg13[(2'h3):(1'h1)] ?
              reg17[(4'h8):(4'h8)] : "6w") <= forvar5[(2'h2):(1'h1)]);
        end
    end
  always
    @(posedge clk) begin
      for (forvar121 = (1'h0); (forvar121 < (2'h3)); forvar121 = (forvar121 + (1'h1)))
        begin
          reg122 <= wire2[(1'h1):(1'h0)];
          reg123 = ((~($signed(reg116[(3'h7):(3'h7)]) ^ "oNpA0ZyALwtR4W1Dyp")) ?
              "lxi" : ($unsigned("kQ3SF") || $unsigned({$unsigned(wire15)})));
        end
      reg124 <= reg24;
    end
  assign wire125 = $signed("O");
  module126 modinst231 (wire230, clk, reg119, wire15, reg25, reg122);
  always
    @(posedge clk) begin
      for (forvar232 = (1'h0); (forvar232 < (2'h2)); forvar232 = (forvar232 + (1'h1)))
        begin
          for (forvar233 = (1'h0); (forvar233 < (1'h1)); forvar233 = (forvar233 + (1'h1)))
            begin
              reg234 = $signed(reg6);
            end
          reg235 <= $signed("8eu");
          reg236 <= (reg23 ?
              {(forvar121[(3'h5):(3'h5)] ?
                      $signed(reg29) : ((wire0 ^ forvar232) ~^ $unsigned(reg115))),
                  ((reg122 << (reg20 << reg111)) ^ (reg111 * (wire32 | reg34)))} : $unsigned(($unsigned("JHkMzG1Vn") ?
                  $unsigned($signed(wire230)) : $signed({(8'hac), wire230}))));
        end
      reg237 <= ($signed({$unsigned($unsigned((7'h44))), "vyJi"}) ?
          reg4[(2'h3):(2'h3)] : $signed({($signed(wire32) || (reg14 ?
                  wire0 : reg6)),
              ({reg27} ? $signed(reg13) : (reg109 & reg116))}));
      for (forvar238 = (1'h0); (forvar238 < (2'h2)); forvar238 = (forvar238 + (1'h1)))
        begin
          for (forvar239 = (1'h0); (forvar239 < (1'h0)); forvar239 = (forvar239 + (1'h1)))
            begin
              reg240 <= reg26[(4'ha):(4'ha)];
              reg241 <= ({forvar28, reg123} ?
                  ($unsigned((8'haa)) * ({"67shsyVR1PBv",
                      $signed(reg27)} >> reg12)) : "0GLgN6mqrIExD53CAK5");
              reg242 = (^~(7'h44));
              reg243 <= ($signed((reg18[(2'h2):(1'h0)] ?
                  {$signed((8'hb7))} : (7'h42))) & $signed((reg122[(3'h6):(2'h2)] ?
                  "EnSueWANB7M5aXhbXs6A" : ("ElvHIP8QStOYQD" && $unsigned((8'hab))))));
              reg244 <= $unsigned(wire230[(2'h3):(1'h1)]);
            end
          reg245 <= "3L8XHZFpFN";
        end
      reg246 <= $unsigned($unsigned("SP9HD"));
      reg247 <= (8'ha6);
    end
  always
    @(posedge clk) begin
      reg248 = forvar233[(3'h4):(2'h3)];
      reg249 <= ((~|reg119[(5'h13):(5'h13)]) ?
          "pKWNG0Jds4PKk7L" : reg237[(3'h5):(3'h4)]);
    end
  always
    @(posedge clk) begin
      for (forvar250 = (1'h0); (forvar250 < (2'h3)); forvar250 = (forvar250 + (1'h1)))
        begin
          reg251 <= $signed("5mw");
        end
      reg252 = $unsigned($signed((^~$signed($unsigned(reg12)))));
    end
  assign wire253 = (("aQycM" ?
                       "HeXd1RSOFZs0r" : reg237[(1'h1):(1'h0)]) != reg27[(1'h0):(1'h0)]);
  module254 modinst282 (wire281, clk, reg29, wire3, reg33, reg123, forvar121);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module254
#( parameter param280 = (({((~^(8'hb7)) ^ ((8'hb5) ? (8'hb7) : (7'h40)))} ? ((((8'had) < (8'hba)) >= (^(8'hb4))) ? ((8'hb0) <<< (~^(8'hbc))) : (-((8'haa) >> (8'hbd)))) : (((~^(8'hb2)) ? {(8'hb6)} : {(8'hb5)}) ? (|(~&(8'hbc))) : (((8'hb2) * (8'ha5)) >>> (~&(8'hb5))))) ~^ ((~^((&(8'ha0)) >= ((8'h9e) ? (8'ha7) : (8'hbd)))) || {(~|((8'ha5) | (8'hb3))), {((8'ha7) ~^ (8'hbd)), ((8'ha7) >> (7'h42))}})) )
(y, clk, wire259, wire258, wire257, wire256, wire255);
  output wire [(32'hee):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire259;
  input wire signed [(4'hb):(1'h0)] wire258;
  input wire signed [(4'hf):(1'h0)] wire257;
  input wire [(3'h6):(1'h0)] wire256;
  input wire [(5'h12):(1'h0)] wire255;
  wire [(4'h8):(1'h0)] wire279;
  reg [(5'h10):(1'h0)] reg278 = (1'h0);
  reg [(4'h9):(1'h0)] reg277 = (1'h0);
  reg [(4'hc):(1'h0)] reg276 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire275;
  reg signed [(3'h7):(1'h0)] reg274 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg273 = (1'h0);
  reg signed [(4'he):(1'h0)] reg272 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg271 = (1'h0);
  reg [(3'h5):(1'h0)] reg270 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg269 = (1'h0);
  reg [(4'hf):(1'h0)] forvar268 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg267 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg266 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg265 = (1'h0);
  reg [(5'h11):(1'h0)] reg264 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar263 = (1'h0);
  reg [(3'h4):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar260 = (1'h0);
  assign y = {wire279,
                 reg278,
                 reg277,
                 reg276,
                 wire275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 forvar268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 forvar263,
                 reg262,
                 reg261,
                 forvar260,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar260 = (1'h0); (forvar260 < (2'h2)); forvar260 = (forvar260 + (1'h1)))
        begin
          reg261 = ("NUQXostL4" ?
              (+(((wire256 >>> wire259) << (wire255 && forvar260)) >> $signed($unsigned(wire257)))) : (^wire259));
          reg262 <= $unsigned($signed($signed(wire258[(2'h3):(1'h0)])));
          for (forvar263 = (1'h0); (forvar263 < (2'h3)); forvar263 = (forvar263 + (1'h1)))
            begin
              reg264 <= ($signed("Z") == $signed((reg262[(2'h3):(1'h0)] ?
                  (~&(wire258 <<< forvar260)) : $unsigned((~^reg261)))));
              reg265 = wire259;
            end
        end
      reg266 = "6lYDXJd9WMQ4";
      reg267 <= ("Hn7tYV3Nuk0DN" >> (~&$unsigned("O3")));
    end
  always
    @(posedge clk) begin
      for (forvar268 = (1'h0); (forvar268 < (2'h3)); forvar268 = (forvar268 + (1'h1)))
        begin
          reg269 <= ($signed($signed((((7'h41) ? reg265 : reg266) ?
                  $unsigned(reg264) : $unsigned(reg265)))) ?
              reg266[(4'hc):(4'ha)] : wire259[(4'hd):(2'h3)]);
          reg270 <= "Wo0";
          reg271 <= $unsigned(wire256[(1'h0):(1'h0)]);
          reg272 <= ($unsigned({$signed("olx")}) && ((reg264 ?
                  reg266[(3'h6):(3'h4)] : forvar263[(2'h2):(2'h2)]) ?
              {($signed(wire259) ? "LQ9qatN9wABprwtyc" : reg270),
                  {(forvar263 ? forvar268 : reg266),
                      {reg267,
                          (7'h43)}}} : $signed(($signed(wire255) && reg266))));
        end
    end
  always
    @(posedge clk) begin
      reg273 <= ($signed(($unsigned((-wire257)) ?
          "bYJU5t6ZRl6z" : {(reg264 < wire255),
              $unsigned((8'hbe))})) >= forvar268);
      reg274 <= "kQIAwal";
    end
  assign wire275 = $unsigned($signed($signed(reg261[(3'h4):(1'h0)])));
  always
    @(posedge clk) begin
      reg276 <= ("KMUkOLOtS" < wire275[(3'h7):(3'h5)]);
      reg277 = "Lprd2pg";
      reg278 = "A6eG9xiPq8";
    end
  assign wire279 = $unsigned((((^(wire255 <<< reg274)) ^ ((reg266 ?
                           reg264 : reg266) ^ $signed(forvar263))) ?
                       "IJ" : $signed({(8'hbe)})));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module126  (y, clk, wire127, wire128, wire129, wire130);
  output wire [(32'h230):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire127;
  input wire signed [(3'h4):(1'h0)] wire128;
  input wire [(5'h11):(1'h0)] wire129;
  input wire signed [(5'h10):(1'h0)] wire130;
  reg [(2'h2):(1'h0)] reg229 = (1'h0);
  reg [(3'h6):(1'h0)] reg228 = (1'h0);
  reg [(5'h15):(1'h0)] forvar227 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg226 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg224 = (1'h0);
  reg [(5'h12):(1'h0)] reg223 = (1'h0);
  reg [(4'h9):(1'h0)] reg222 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg220 = (1'h0);
  reg [(5'h11):(1'h0)] reg219 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg218 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar217 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg216 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg215 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg214 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg213 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg212 = (1'h0);
  reg [(4'hb):(1'h0)] reg211 = (1'h0);
  reg [(3'h5):(1'h0)] forvar210 = (1'h0);
  reg [(5'h14):(1'h0)] forvar209 = (1'h0);
  wire [(3'h6):(1'h0)] wire208;
  reg signed [(4'hd):(1'h0)] reg207 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg206 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire205;
  wire [(2'h2):(1'h0)] wire204;
  reg [(3'h4):(1'h0)] reg203 = (1'h0);
  reg [(4'hc):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg201 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg131 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar132 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg134 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg135 = (1'h0);
  reg [(3'h5):(1'h0)] reg136 = (1'h0);
  reg [(5'h13):(1'h0)] reg137 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg138 = (1'h0);
  wire [(5'h11):(1'h0)] wire139;
  reg [(5'h14):(1'h0)] reg140 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar141 = (1'h0);
  reg [(5'h15):(1'h0)] reg142 = (1'h0);
  reg [(3'h5):(1'h0)] reg143 = (1'h0);
  reg [(2'h3):(1'h0)] reg144 = (1'h0);
  reg [(4'h8):(1'h0)] reg145 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg146 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire147;
  reg [(4'h8):(1'h0)] reg148 = (1'h0);
  reg [(4'he):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg150 = (1'h0);
  reg [(4'h9):(1'h0)] reg151 = (1'h0);
  reg [(5'h10):(1'h0)] reg152 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg153 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire199;
  assign y = {reg229,
                 reg228,
                 forvar227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 forvar217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 forvar210,
                 forvar209,
                 wire208,
                 reg207,
                 reg206,
                 wire205,
                 wire204,
                 reg203,
                 reg202,
                 reg201,
                 reg131,
                 forvar132,
                 reg133,
                 reg134,
                 reg135,
                 reg136,
                 reg137,
                 reg138,
                 wire139,
                 reg140,
                 forvar141,
                 reg142,
                 reg143,
                 reg144,
                 reg145,
                 reg146,
                 wire147,
                 reg148,
                 reg149,
                 reg150,
                 reg151,
                 reg152,
                 reg153,
                 wire199,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg131 <= "uu";
    end
  always
    @(posedge clk) begin
      for (forvar132 = (1'h0); (forvar132 < (1'h1)); forvar132 = (forvar132 + (1'h1)))
        begin
          reg133 <= $signed(($signed(wire130) ?
              (~|("z91" ? (&wire127) : (forvar132 >= (8'hae)))) : "EiZJF"));
          reg134 <= {$signed((!((~(8'hb0)) ?
                  ((8'ha9) >>> wire130) : "HElt4g4lkszK8kV"))),
              "BFpD0"};
          reg135 <= reg134[(3'h6):(3'h6)];
          reg136 <= wire130;
          reg137 <= "DeQ6JxCx9sop4ePpXCS1";
        end
      reg138 <= (($unsigned({(&(8'h9c)), {wire129}}) > "xhm7fzpI9a") ?
          ($unsigned(((8'hb6) << wire129[(4'ha):(3'h5)])) >>> reg137[(1'h0):(1'h0)]) : $unsigned(((wire128 > "5Kqu") < reg137)));
    end
  assign wire139 = wire130;
  always
    @(posedge clk) begin
      reg140 <= $signed(($unsigned({$unsigned(reg135),
          $signed(wire127)}) >= {$signed((forvar132 ? reg131 : wire128)),
          "44UD4M8ca43"}));
      for (forvar141 = (1'h0); (forvar141 < (2'h2)); forvar141 = (forvar141 + (1'h1)))
        begin
          reg142 <= "P5";
          reg143 = ((~^{"ei5NwLW2m"}) ? reg135[(2'h3):(1'h0)] : "Dh");
        end
    end
  always
    @(posedge clk) begin
      reg144 <= "pgONbp8eQ3";
    end
  always
    @(posedge clk) begin
      reg145 <= (reg142[(5'h11):(3'h6)] ?
          $unsigned((reg142 ?
              reg133 : ((reg143 + reg135) ?
                  $signed((8'hbf)) : wire129))) : ((("XBW5gIHVhnRfln" & $signed(wire130)) | $unsigned($signed((8'h9d)))) ?
              (wire130[(4'he):(4'hb)] ?
                  "uSQgb4r3rnXpqXU" : "4v") : (wire129[(1'h0):(1'h0)] ^ (reg131[(3'h5):(2'h2)] ?
                  $unsigned(reg134) : (~&wire130)))));
      reg146 = $signed($unsigned(reg131));
    end
  assign wire147 = reg137[(4'he):(4'hb)];
  always
    @(posedge clk) begin
      reg148 = reg144;
      reg149 = {wire147[(3'h5):(2'h3)]};
      reg150 <= (~^((~^reg145[(1'h0):(1'h0)]) != ({"huC3tM",
              (wire129 ? reg138 : forvar132)} ?
          {((8'ha1) ? wire128 : reg142)} : {(wire129 ? wire128 : forvar141),
              reg144})));
    end
  always
    @(posedge clk) begin
      reg151 <= $unsigned((forvar141[(3'h4):(1'h1)] ?
          ((wire127 + wire147[(1'h1):(1'h1)]) >>> $unsigned("yUZOLTh")) : "Ax"));
    end
  always
    @(posedge clk) begin
      reg152 <= reg133[(3'h4):(3'h4)];
      reg153 = reg146;
    end
  module154 modinst200 (.wire157(reg142), .wire156(reg134), .wire155(reg138), .wire159(reg140), .clk(clk), .y(wire199), .wire158(wire147));
  always
    @(posedge clk) begin
      reg201 <= ((8'ha7) ? (~|"") : wire128[(2'h2):(2'h2)]);
      reg202 <= "JH";
    end
  always
    @(posedge clk) begin
      reg203 <= "MblQ661tQa1LKRQ";
    end
  assign wire204 = "sxHbGkQKOhB7e3Y";
  assign wire205 = "HKI8B0bzf6xmf8p5xpr";
  always
    @(posedge clk) begin
      reg206 <= reg201[(4'hb):(3'h4)];
      reg207 <= ($unsigned((+"qqVAl")) >= wire139);
    end
  assign wire208 = $signed(wire130);
  always
    @(posedge clk) begin
      for (forvar209 = (1'h0); (forvar209 < (1'h1)); forvar209 = (forvar209 + (1'h1)))
        begin
          for (forvar210 = (1'h0); (forvar210 < (3'h4)); forvar210 = (forvar210 + (1'h1)))
            begin
              reg211 <= wire199[(2'h2):(2'h2)];
              reg212 <= {reg153[(4'ha):(2'h3)]};
              reg213 <= ((({(&reg144), (forvar132 ? reg138 : reg212)} ?
                  (^~(reg137 >> (8'haa))) : wire147) + $unsigned("A")) ^ forvar132[(3'h4):(1'h1)]);
              reg214 <= "De";
            end
          reg215 <= $signed(reg131[(3'h4):(1'h0)]);
          reg216 <= "ZKL";
        end
      for (forvar217 = (1'h0); (forvar217 < (1'h1)); forvar217 = (forvar217 + (1'h1)))
        begin
          reg218 <= ({forvar210[(3'h5):(2'h2)],
              reg151} * $unsigned($signed((8'hbb))));
          reg219 <= (("ixIqc03KcvvQk" ^~ reg146[(1'h0):(1'h0)]) < (-$signed((^~"IvswQ6hPa7KzTT"))));
        end
      reg220 <= wire204;
      reg221 <= ("LqVWYfOYevlNS" ? reg145 : wire204);
      reg222 <= {((|{$signed(wire147),
              (forvar217 ?
                  (8'h9d) : reg151)}) <<< $signed((+(reg143 && reg218))))};
    end
  always
    @(posedge clk) begin
      reg223 = $signed("");
      reg224 <= "6wwGwvFnMU99JeEwQVbZ";
      reg225 <= wire127;
      reg226 = {(~&(|reg134[(4'h9):(3'h7)]))};
    end
  always
    @(posedge clk) begin
      for (forvar227 = (1'h0); (forvar227 < (1'h1)); forvar227 = (forvar227 + (1'h1)))
        begin
          reg228 <= (($signed({"YpKgn"}) ? $signed((+wire208)) : forvar227) ?
              $signed(forvar227) : (|(-$unsigned((-reg138)))));
          reg229 <= ("" ? $signed({wire129[(2'h2):(1'h1)]}) : forvar217);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module36
#(parameter param106 = (8'hab))
(y, clk, wire40, wire39, wire38, wire37);
  output wire [(32'h305):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire40;
  input wire signed [(4'hb):(1'h0)] wire39;
  input wire [(5'h11):(1'h0)] wire38;
  input wire signed [(3'h4):(1'h0)] wire37;
  reg signed [(3'h5):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg103 = (1'h0);
  reg [(4'hb):(1'h0)] reg102 = (1'h0);
  wire [(5'h13):(1'h0)] wire101;
  wire [(4'he):(1'h0)] wire100;
  wire [(4'ha):(1'h0)] wire99;
  wire [(4'h8):(1'h0)] wire98;
  reg [(3'h4):(1'h0)] reg97 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg96 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar95 = (1'h0);
  reg [(3'h7):(1'h0)] reg94 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg93 = (1'h0);
  reg [(5'h15):(1'h0)] reg92 = (1'h0);
  reg [(3'h4):(1'h0)] reg91 = (1'h0);
  reg [(3'h4):(1'h0)] reg90 = (1'h0);
  reg [(3'h6):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar88 = (1'h0);
  reg [(5'h13):(1'h0)] reg87 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar86 = (1'h0);
  reg [(5'h15):(1'h0)] reg85 = (1'h0);
  reg [(4'he):(1'h0)] reg84 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg83 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg82 = (1'h0);
  reg [(5'h14):(1'h0)] reg81 = (1'h0);
  reg [(5'h14):(1'h0)] reg80 = (1'h0);
  reg [(4'h8):(1'h0)] forvar79 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg78 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg77 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg76 = (1'h0);
  reg [(3'h7):(1'h0)] reg75 = (1'h0);
  reg [(3'h6):(1'h0)] reg74 = (1'h0);
  reg [(5'h11):(1'h0)] reg73 = (1'h0);
  reg [(3'h5):(1'h0)] reg72 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg71 = (1'h0);
  reg [(5'h11):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg69 = (1'h0);
  reg [(2'h3):(1'h0)] reg68 = (1'h0);
  reg [(5'h13):(1'h0)] reg67 = (1'h0);
  reg [(5'h12):(1'h0)] forvar66 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg65 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg64 = (1'h0);
  reg [(4'ha):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg62 = (1'h0);
  reg [(4'he):(1'h0)] reg61 = (1'h0);
  reg [(2'h3):(1'h0)] reg60 = (1'h0);
  reg [(5'h13):(1'h0)] reg59 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg57 = (1'h0);
  reg [(4'h9):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg55 = (1'h0);
  reg [(4'hf):(1'h0)] reg54 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg53 = (1'h0);
  reg [(2'h2):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg51 = (1'h0);
  reg [(5'h15):(1'h0)] reg50 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar49 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar48 = (1'h0);
  wire [(2'h3):(1'h0)] wire47;
  wire [(5'h13):(1'h0)] wire46;
  wire signed [(4'hd):(1'h0)] wire45;
  reg [(4'hb):(1'h0)] reg44 = (1'h0);
  reg [(3'h7):(1'h0)] reg43 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg41 = (1'h0);
  assign y = {reg105,
                 reg104,
                 reg103,
                 reg102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 reg97,
                 reg96,
                 forvar95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 forvar88,
                 reg87,
                 forvar86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 forvar79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 forvar66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 forvar49,
                 forvar48,
                 wire47,
                 wire46,
                 wire45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg41 = (~&((wire37[(2'h3):(2'h3)] ?
          wire38 : $signed($unsigned((8'hbe)))) <<< $signed((8'hb5))));
      reg42 = wire37[(2'h3):(1'h0)];
      reg43 <= "";
      reg44 <= ("p6x2T0M7FWD" < "d");
    end
  assign wire45 = "8JY2";
  assign wire46 = (^~"RHLI");
  assign wire47 = reg41;
  always
    @(posedge clk) begin
      for (forvar48 = (1'h0); (forvar48 < (2'h2)); forvar48 = (forvar48 + (1'h1)))
        begin
          for (forvar49 = (1'h0); (forvar49 < (1'h1)); forvar49 = (forvar49 + (1'h1)))
            begin
              reg50 = wire47;
              reg51 <= wire37;
              reg52 <= ((forvar49 ?
                  reg42[(5'h12):(2'h2)] : wire37) * wire39[(4'ha):(3'h6)]);
              reg53 <= $signed(wire46[(4'hd):(1'h0)]);
              reg54 = ("5v" ? wire37 : $unsigned(wire38[(1'h0):(1'h0)]));
            end
          reg55 <= {wire46[(4'h9):(3'h7)]};
          reg56 <= ((reg52[(1'h0):(1'h0)] ?
              reg43[(3'h7):(1'h0)] : $unsigned("ine4MAIIa4ipsXs")) >> wire38[(5'h11):(4'he)]);
          reg57 = reg54;
          reg58 <= ((+(-("3hPWSyOm4thzc0Bv" ?
              $signed(wire37) : $unsigned(forvar48)))) ~^ ($unsigned(reg41[(1'h0):(1'h0)]) ^~ $signed(reg41[(2'h3):(1'h0)])));
        end
      reg59 <= $unsigned($unsigned(reg54));
      reg60 <= (("0ZZaLLN6E3rcIH6" ?
          (!"ZkRudq8bc9F") : reg57[(4'h8):(3'h6)]) >> (reg59[(4'hd):(3'h7)] ?
          reg59[(3'h6):(3'h5)] : $unsigned(reg57)));
      reg61 <= "";
      reg62 <= reg54[(4'h8):(3'h7)];
    end
  always
    @(posedge clk) begin
      reg63 <= ((wire40 ?
          {($unsigned((8'hb0)) >> $signed(reg55)),
              (|{wire37})} : reg61) > reg56);
      reg64 <= (+$unsigned($signed((reg59[(4'hf):(4'he)] ?
          (~reg44) : (~&(7'h44))))));
      reg65 <= "CP8wza1eFDNMoh5";
    end
  always
    @(posedge clk) begin
      for (forvar66 = (1'h0); (forvar66 < (2'h2)); forvar66 = (forvar66 + (1'h1)))
        begin
          reg67 = $signed((&reg42[(4'he):(4'ha)]));
          if ("KY15t18O")
            begin
              reg68 <= wire40[(3'h5):(3'h5)];
              reg69 = {reg68,
                  ((+($signed(reg50) ?
                      $unsigned(reg68) : $unsigned(reg53))) ^ (wire38[(5'h11):(4'hf)] - ($signed((7'h44)) <= $signed(reg53))))};
              reg70 <= (~^reg69);
              reg71 <= $signed(reg52);
              reg72 <= reg51;
            end
          else
            begin
              reg68 <= (({(((8'hb6) ? forvar48 : wire39) ?
                      ((8'h9d) ?
                          reg62 : reg58) : (!(8'ha3)))} != (+(^~$unsigned((8'hb3))))) > reg68);
              reg69 <= "";
              reg70 <= (wire38[(2'h3):(1'h0)] ?
                  wire38[(3'h4):(3'h4)] : {($signed(reg41) ?
                          $unsigned($signed(reg72)) : ("zEEw6kkO" ?
                              (reg65 ? reg71 : reg42) : (reg67 ?
                                  wire40 : wire39)))});
              reg71 <= {(~^wire38)};
            end
          reg73 <= ("O0" >> "npXaoMz97MOZd");
          if (wire37)
            begin
              reg74 = reg67[(4'hb):(2'h3)];
              reg75 <= (+reg41);
              reg76 = $signed({reg42, $signed((~^{reg54}))});
            end
          else
            begin
              reg74 <= "ti4ige0K";
              reg75 <= ("HkY3bpq1elb5JE" ~^ $signed($unsigned(((reg52 ?
                      (8'hb8) : reg42) ?
                  wire38 : $unsigned(reg58)))));
              reg76 <= (8'h9c);
              reg77 <= "doSV";
            end
        end
      reg78 <= "8";
    end
  always
    @(posedge clk) begin
      for (forvar79 = (1'h0); (forvar79 < (2'h2)); forvar79 = (forvar79 + (1'h1)))
        begin
          reg80 <= {("" ?
                  ({"w"} ?
                      (wire45 > wire45) : reg54[(3'h4):(2'h3)]) : $unsigned(($signed(reg56) && "Tuq5M6Xn"))),
              (reg54 << wire39[(3'h6):(1'h0)])};
        end
      reg81 <= "B";
      reg82 <= (^~reg76[(2'h3):(2'h2)]);
      reg83 <= $unsigned((wire46 ?
          ($signed(reg43[(1'h1):(1'h1)]) == wire45) : ("o9alUv7Jitx" ?
              reg65 : "Cl4AHo21ugg0y84Oba9")));
      reg84 = $signed("NDi1");
    end
  always
    @(posedge clk) begin
      reg85 <= "BUhVucQW7";
      for (forvar86 = (1'h0); (forvar86 < (1'h1)); forvar86 = (forvar86 + (1'h1)))
        begin
          reg87 = ((~^(!$signed((reg65 - reg76)))) ?
              forvar48[(2'h3):(2'h2)] : ({$unsigned((forvar49 > reg50))} < $signed("gzSeeEgKC")));
          for (forvar88 = (1'h0); (forvar88 < (2'h3)); forvar88 = (forvar88 + (1'h1)))
            begin
              reg89 <= (8'hb3);
            end
          reg90 = $unsigned((+"HbHUMGmZcoWwWff"));
          if ($signed((reg89[(3'h5):(2'h3)] ?
              (+((reg63 ? reg58 : reg78) >> {forvar66,
                  reg62})) : "DogZwnaGIqxKCkErJCM")))
            begin
              reg91 <= "cpxL";
              reg92 = wire45;
            end
          else
            begin
              reg91 <= "QwFHaA";
              reg92 = ((forvar49[(3'h4):(1'h0)] ?
                      (reg92[(5'h11):(2'h3)] << {{(7'h40),
                              forvar49}}) : "NkR9IkT") ?
                  $signed({({reg82, reg57} ?
                          (reg92 ?
                              wire46 : reg55) : $signed((8'hb2)))}) : reg77);
            end
          reg93 <= (reg74 ^~ {reg81[(5'h14):(5'h11)]});
        end
      reg94 <= forvar66[(5'h12):(1'h0)];
      for (forvar95 = (1'h0); (forvar95 < (1'h0)); forvar95 = (forvar95 + (1'h1)))
        begin
          reg96 <= (reg64[(1'h0):(1'h0)] >> reg93);
        end
    end
  always
    @(posedge clk) begin
      reg97 <= $unsigned(reg89);
    end
  assign wire98 = ($unsigned((~reg67[(2'h2):(1'h0)])) ^~ reg59);
  assign wire99 = "PECx6Zb";
  assign wire100 = reg82[(4'ha):(4'ha)];
  assign wire101 = wire40;
  always
    @(posedge clk) begin
      reg102 <= (^~wire40[(3'h5):(2'h3)]);
      reg103 <= ((!(reg81[(4'ha):(1'h0)] <= reg72)) && $unsigned({reg43,
          wire101[(4'hf):(4'he)]}));
      reg104 <= ((!reg75) == "k4PuM79MDet70Pcbk");
      reg105 <= ((8'ha2) ?
          {($signed(reg71) <= ((~^wire45) ?
                  $unsigned(wire46) : "U9hr4KqcU8Pem7llc8"))} : wire47);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module154
#( parameter param197 = ((&((((8'hbd) * (7'h40)) ? (!(8'h9f)) : {(7'h42)}) ? (((8'haf) << (8'hb6)) ? ((8'h9f) * (8'ha2)) : ((7'h40) ? (8'hb3) : (8'hae))) : (-{(8'hb0)}))) ? {(~&{((8'hac) ? (8'hb1) : (8'hb4)), ((8'hb2) ? (8'hb4) : (8'h9c))}), ((((8'hb8) ? (8'ha0) : (8'hb2)) ? ((8'h9d) <<< (8'ha9)) : (!(8'hb7))) > (~{(8'hbd), (8'ha7)}))} : ((~&{((8'hb7) ? (8'ha1) : (8'ha7))}) | (^(((7'h42) ? (7'h42) : (8'haa)) >> ((8'hb8) ? (8'hb4) : (7'h42))))))
, parameter param198 = param197 )
(y, clk, wire159, wire158, wire157, wire156, wire155);
  output wire [(32'h190):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire159;
  input wire [(5'h13):(1'h0)] wire158;
  input wire signed [(5'h15):(1'h0)] wire157;
  input wire [(5'h14):(1'h0)] wire156;
  input wire signed [(3'h7):(1'h0)] wire155;
  reg [(4'h9):(1'h0)] reg196 = (1'h0);
  reg [(5'h11):(1'h0)] reg195 = (1'h0);
  reg [(3'h7):(1'h0)] reg194 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg192 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg191 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg190 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar189 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg188 = (1'h0);
  reg [(4'hf):(1'h0)] reg187 = (1'h0);
  reg [(4'hb):(1'h0)] reg186 = (1'h0);
  reg [(5'h12):(1'h0)] reg185 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire184;
  reg [(4'he):(1'h0)] reg183 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire182;
  reg [(4'hb):(1'h0)] reg181 = (1'h0);
  reg [(3'h6):(1'h0)] reg180 = (1'h0);
  reg [(4'he):(1'h0)] reg179 = (1'h0);
  reg [(4'hb):(1'h0)] reg178 = (1'h0);
  reg [(3'h6):(1'h0)] reg177 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg176 = (1'h0);
  reg [(4'ha):(1'h0)] reg175 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg174 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg173 = (1'h0);
  reg [(5'h10):(1'h0)] forvar172 = (1'h0);
  reg [(4'hd):(1'h0)] reg171 = (1'h0);
  reg [(2'h2):(1'h0)] reg170 = (1'h0);
  reg [(3'h7):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg166 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg164 = (1'h0);
  reg [(2'h3):(1'h0)] reg163 = (1'h0);
  reg [(3'h4):(1'h0)] forvar162 = (1'h0);
  reg [(5'h12):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar160 = (1'h0);
  assign y = {reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 forvar189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 wire184,
                 reg183,
                 wire182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 forvar172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 forvar162,
                 reg161,
                 forvar160,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar160 = (1'h0); (forvar160 < (1'h0)); forvar160 = (forvar160 + (1'h1)))
        begin
          reg161 <= $signed((-wire155));
          for (forvar162 = (1'h0); (forvar162 < (2'h3)); forvar162 = (forvar162 + (1'h1)))
            begin
              reg163 = (8'hbf);
              reg164 <= ((8'hb1) << ($signed(wire157) ?
                  (~^reg161[(2'h2):(1'h1)]) : (!(-(~wire156)))));
              reg165 <= forvar160;
              reg166 <= (reg165[(2'h3):(1'h1)] ?
                  (reg163 && (8'ha9)) : "UYLTNMtq1OaLWsLZ5");
              reg167 <= $signed("W1e");
            end
          reg168 <= (((|{{reg165}, (&forvar162)}) ?
                  ((8'hbf) || {$signed(wire156)}) : wire158[(5'h10):(2'h2)]) ?
              wire155 : $unsigned(($signed("qTvEWsCzd53FagpvqdZ") ?
                  $unsigned((~(8'hb9))) : wire156)));
          reg169 <= (+reg167[(3'h4):(1'h0)]);
        end
      reg170 <= {(wire157 != reg163[(2'h2):(1'h0)])};
      reg171 <= "N4xSiMnYM3p5GV0779NF";
    end
  always
    @(posedge clk) begin
      for (forvar172 = (1'h0); (forvar172 < (3'h4)); forvar172 = (forvar172 + (1'h1)))
        begin
          reg173 <= wire156;
          reg174 <= (((^~$signed("9tZKYAbp")) + $signed(($unsigned(wire158) ?
                  $signed(reg167) : wire156))) ?
              ((wire155[(3'h4):(3'h4)] & {{reg168, reg161},
                  wire155}) >>> (((reg163 ? reg171 : reg165) ?
                  $unsigned(reg169) : "blTxRPeTrgS0W20KF") ^~ ($signed((8'hb4)) ?
                  (reg170 >> (7'h40)) : $signed(reg173)))) : wire159);
          reg175 <= ((($unsigned("yApKgt") >>> reg174) ?
              (("tOZlzg6ztAvnfu6dxZ" <= wire155) ?
                  ({wire159,
                      reg165} < (reg161 ~^ (8'hb4))) : {reg170[(1'h1):(1'h1)]}) : (~{reg170[(1'h0):(1'h0)]})) <<< reg170[(2'h2):(1'h1)]);
        end
    end
  always
    @(posedge clk) begin
      reg176 = reg163[(1'h1):(1'h1)];
      reg177 <= (-(("mYEiyRgsGiaL" ^ {"rhEdnrEq7KsWLim7w", $signed(reg164)}) ?
          wire155 : forvar162[(1'h0):(1'h0)]));
      reg178 <= (~^($unsigned(reg176) * {$unsigned(wire159[(3'h5):(1'h1)])}));
    end
  always
    @(posedge clk) begin
      reg179 <= {wire156[(4'hf):(4'he)], reg165};
    end
  always
    @(posedge clk) begin
      reg180 <= ((reg166 ?
          wire157 : reg177[(3'h6):(1'h0)]) || wire159[(3'h5):(1'h0)]);
      reg181 <= (~^($unsigned((&"evObcgdMxd6F")) <<< $signed(($signed((8'hb4)) ?
          (|(8'hb1)) : "NDCq"))));
    end
  assign wire182 = wire156[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg183 <= "h";
    end
  assign wire184 = $signed(($unsigned(((~|wire182) ?
                       (reg167 || wire182) : "")) ^ reg183[(3'h4):(1'h0)]));
  always
    @(posedge clk) begin
      reg185 <= {{$unsigned((|(^~(8'hb7))))}};
      reg186 <= (wire159[(1'h0):(1'h0)] ?
          (reg173[(2'h2):(1'h0)] != $signed(reg168)) : $signed(wire184));
      reg187 <= "yu8TRAT2qsxrnK11K";
      reg188 <= ({$signed("xuFRYHRV")} ?
          $unsigned((+(wire184 ?
              (&reg180) : reg168[(3'h7):(3'h7)]))) : (("sIf2x6oeJuNcOVsx" >>> (((8'hb4) ?
                  wire156 : reg179) < "4dnk")) ?
              (forvar160 ?
                  (reg165[(3'h6):(1'h0)] ?
                      ((8'h9c) ?
                          wire184 : (8'ha7)) : $unsigned(wire156)) : $signed((reg164 - wire156))) : reg174));
    end
  always
    @(posedge clk) begin
      for (forvar189 = (1'h0); (forvar189 < (1'h1)); forvar189 = (forvar189 + (1'h1)))
        begin
          reg190 <= wire182;
          reg191 = (~&$signed($signed(((reg178 ~^ wire182) ?
              (reg186 | reg177) : reg173[(2'h3):(1'h0)]))));
        end
    end
  always
    @(posedge clk) begin
      reg192 <= reg176[(2'h3):(1'h1)];
      reg193 <= "Ut07XNXFwuZ";
      reg194 <= (!(($signed("IP") + {{reg191, reg183},
          reg170}) << ($unsigned($unsigned(forvar172)) ?
          (~^{reg178}) : reg164[(1'h1):(1'h0)])));
      reg195 <= ($signed("VNwCPXWCI4") ?
          (-(reg161[(2'h2):(1'h1)] < reg169[(2'h3):(2'h3)])) : ($signed(wire157) * ((8'hb4) != reg186)));
      reg196 <= reg176;
    end
endmodule