(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param1001 = (~{(~|({(8'ha9)} <<< (^~(8'ha0)))), ((((8'haf) - (8'hbe)) ? {(8'hb1)} : (-(8'ha8))) ? {(~^(8'hbe))} : (~&{(8'hab)}))}) )
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h205):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire0;
  input wire [(5'h14):(1'h0)] wire1;
  input wire [(5'h10):(1'h0)] wire2;
  input wire [(5'h14):(1'h0)] wire3;
  input wire [(2'h3):(1'h0)] wire4;
  wire [(4'h9):(1'h0)] wire1000;
  wire signed [(5'h15):(1'h0)] wire5;
  wire signed [(5'h13):(1'h0)] wire6;
  wire [(5'h14):(1'h0)] wire961;
  wire signed [(2'h3):(1'h0)] wire963;
  reg signed [(5'h15):(1'h0)] reg964 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire965;
  wire [(5'h12):(1'h0)] wire966;
  wire signed [(3'h7):(1'h0)] wire967;
  wire signed [(4'h8):(1'h0)] wire968;
  wire signed [(5'h15):(1'h0)] wire969;
  wire [(4'hb):(1'h0)] wire970;
  wire signed [(5'h15):(1'h0)] wire972;
  wire signed [(4'hd):(1'h0)] wire974;
  wire signed [(5'h11):(1'h0)] wire975;
  wire [(5'h10):(1'h0)] wire976;
  wire signed [(2'h2):(1'h0)] wire977;
  reg signed [(4'h9):(1'h0)] reg978 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg979 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg980 = (1'h0);
  reg [(4'hb):(1'h0)] reg981 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg982 = (1'h0);
  reg [(4'ha):(1'h0)] reg983 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg984 = (1'h0);
  reg [(5'h13):(1'h0)] reg985 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg986 = (1'h0);
  reg [(4'he):(1'h0)] reg987 = (1'h0);
  reg [(5'h15):(1'h0)] reg988 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg989 = (1'h0);
  reg [(3'h7):(1'h0)] reg990 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg991 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg992 = (1'h0);
  reg [(5'h10):(1'h0)] reg993 = (1'h0);
  reg [(5'h10):(1'h0)] reg994 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg995 = (1'h0);
  reg [(5'h12):(1'h0)] reg996 = (1'h0);
  wire signed [(4'he):(1'h0)] wire997;
  wire signed [(4'hf):(1'h0)] wire998;
  assign y = {wire1000,
                 wire5,
                 wire6,
                 wire961,
                 wire963,
                 reg964,
                 wire965,
                 wire966,
                 wire967,
                 wire968,
                 wire969,
                 wire970,
                 wire972,
                 wire974,
                 wire975,
                 wire976,
                 wire977,
                 reg978,
                 reg979,
                 reg980,
                 reg981,
                 reg982,
                 reg983,
                 reg984,
                 reg985,
                 reg986,
                 reg987,
                 reg988,
                 reg989,
                 reg990,
                 reg991,
                 reg992,
                 reg993,
                 reg994,
                 reg995,
                 reg996,
                 wire997,
                 wire998,
                 (1'h0)};
  assign wire5 = (|wire2[(1'h1):(1'h1)]);
  assign wire6 = (wire4[(2'h2):(2'h2)] >> wire3);
  module7 modinst962 (wire961, clk, wire1, wire3, wire5, wire0);
  assign wire963 = $unsigned((wire5 >= $unsigned(((wire961 ?
                       wire6 : wire2) * (wire6 - wire4)))));
  always
    @(posedge clk) begin
      reg964 <= wire6;
    end
  assign wire965 = ((-wire6) << ((wire6 > $signed($signed(wire3))) ?
                       wire6 : wire0[(5'h12):(5'h10)]));
  assign wire966 = {(~|wire965[(2'h3):(2'h2)])};
  assign wire967 = ($signed(wire961) ?
                       (!$unsigned($signed($signed((8'h9f))))) : (~^wire3[(4'hf):(4'hd)]));
  assign wire968 = wire965;
  assign wire969 = ({({(wire967 <= (8'hbf))} ?
                           wire2[(3'h6):(2'h2)] : $unsigned((wire5 ?
                               wire0 : (8'h9f))))} == (|$signed(($unsigned(wire968) ?
                       wire961[(5'h10):(4'hf)] : (wire1 ? wire2 : wire2)))));
  module12 modinst971 (wire970, clk, wire3, wire0, reg964, wire965);
  module239 modinst973 (wire972, clk, wire5, wire970, reg964, wire961);
  assign wire974 = ((+(((wire966 ? wire967 : wire972) > wire1) ?
                       wire968 : (^wire3[(3'h5):(3'h4)]))) & $signed((~&(^~{wire0}))));
  assign wire975 = wire972[(3'h5):(2'h2)];
  assign wire976 = ({($unsigned($unsigned(wire1)) != $unsigned(reg964[(4'h8):(2'h3)])),
                           $unsigned($signed({(8'haa)}))} ?
                       $unsigned(reg964) : {wire2[(4'hd):(4'ha)],
                           reg964[(5'h15):(4'hd)]});
  assign wire977 = {$unsigned((wire1 ? (8'ha8) : $unsigned($signed(wire972))))};
  always
    @(posedge clk) begin
      if ($unsigned((~^(wire965[(3'h7):(3'h5)] ? $unsigned(wire2) : wire974))))
        begin
          reg978 <= (8'ha3);
          reg979 <= wire3;
        end
      else
        begin
          if ($signed(wire965[(2'h2):(2'h2)]))
            begin
              reg978 <= wire968;
              reg979 <= reg964;
              reg980 <= wire1;
              reg981 <= $signed(reg978[(4'h8):(3'h6)]);
              reg982 <= $unsigned({(((^wire963) ^ (reg964 ? wire4 : reg981)) ?
                      {wire6} : {(reg981 + wire977), wire5}),
                  (~^((reg980 ? wire975 : wire4) ?
                      wire974[(1'h0):(1'h0)] : wire6))});
            end
          else
            begin
              reg978 <= wire968;
              reg979 <= $signed($unsigned(((wire5[(3'h7):(3'h7)] ?
                  (wire1 ? reg964 : reg978) : (wire965 ?
                      (8'hae) : (7'h43))) * (~|(+wire5)))));
            end
          reg983 <= $unsigned(((^~$unsigned({reg964,
              wire966})) && $signed((8'hb3))));
          reg984 <= wire0;
          if ((((+wire1) - wire967) ?
              $unsigned($unsigned($unsigned((reg964 ^~ reg983)))) : (~$signed(wire966))))
            begin
              reg985 <= $signed({(-{wire977[(2'h2):(1'h0)], (^wire968)})});
              reg986 <= wire976;
              reg987 <= wire967[(1'h0):(1'h0)];
            end
          else
            begin
              reg985 <= $unsigned((~&reg984));
            end
        end
      if ($unsigned($unsigned(wire976)))
        begin
          if (wire2)
            begin
              reg988 <= ($unsigned(((~^$signed(wire961)) && ((wire966 ?
                          wire1 : wire970) ?
                      ((8'hb8) ? reg983 : wire5) : wire961))) ?
                  $unsigned($unsigned($unsigned((wire977 ?
                      reg984 : wire963)))) : $unsigned(wire0[(4'hf):(2'h3)]));
              reg989 <= $signed({reg982[(4'he):(4'h8)], wire0});
            end
          else
            begin
              reg988 <= $unsigned(wire963[(1'h0):(1'h0)]);
              reg989 <= (~&((+{reg982}) ?
                  $unsigned(((wire961 != wire974) + $unsigned(wire963))) : wire972));
              reg990 <= (~|wire961);
            end
          if (wire1)
            begin
              reg991 <= wire3;
              reg992 <= $signed((-wire970[(3'h4):(2'h3)]));
              reg993 <= reg983[(2'h3):(1'h0)];
            end
          else
            begin
              reg991 <= wire968;
              reg992 <= $signed({$unsigned((~$unsigned((8'hbb))))});
              reg993 <= {$signed(wire963),
                  (($signed((reg989 >= wire5)) ?
                      wire4 : wire967) * (((reg980 <= reg988) <<< $signed(reg989)) >> {$unsigned(reg978)}))};
              reg994 <= $signed(wire961);
            end
          reg995 <= $unsigned(((((~^wire5) >= $signed(reg991)) || reg980) ?
              reg986 : $signed({$unsigned((8'h9c)), (~^wire961)})));
        end
      else
        begin
          reg988 <= (wire4[(2'h3):(1'h1)] || (wire970 >= (reg978[(1'h0):(1'h0)] ?
              {$signed((8'hb3)),
                  {(8'hab), (8'haf)}} : $unsigned((wire968 < wire3)))));
          reg989 <= $unsigned(reg985);
          reg990 <= (~&$signed((+((wire5 ?
              wire4 : reg981) >= reg989[(1'h1):(1'h0)]))));
        end
      reg996 <= (8'hb4);
    end
  assign wire997 = {{(wire968 & (+((8'hb3) ? reg980 : reg988)))},
                       {$signed(((wire969 ^ reg980) ?
                               wire967 : $signed(reg987))),
                           {{reg995, (~&reg995)}}}};
  module190 modinst999 (.clk(clk), .wire195(wire961), .wire193(reg995), .wire191(reg996), .y(wire998), .wire194(reg994), .wire192(wire6));
  assign wire1000 = wire5;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module7  (y, clk, wire11, wire10, wire9, wire8);
  output wire [(32'hb1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire11;
  input wire signed [(5'h14):(1'h0)] wire10;
  input wire signed [(5'h15):(1'h0)] wire9;
  input wire signed [(5'h15):(1'h0)] wire8;
  wire [(3'h5):(1'h0)] wire960;
  wire signed [(3'h7):(1'h0)] wire959;
  wire [(4'h9):(1'h0)] wire958;
  wire signed [(5'h11):(1'h0)] wire957;
  wire signed [(3'h5):(1'h0)] wire956;
  wire signed [(5'h12):(1'h0)] wire955;
  wire signed [(5'h12):(1'h0)] wire953;
  wire signed [(3'h4):(1'h0)] wire952;
  wire signed [(2'h2):(1'h0)] wire951;
  wire signed [(4'hd):(1'h0)] wire950;
  wire [(5'h14):(1'h0)] wire949;
  wire [(4'h9):(1'h0)] wire948;
  wire [(3'h5):(1'h0)] wire947;
  wire [(4'ha):(1'h0)] wire946;
  wire [(5'h15):(1'h0)] wire945;
  wire signed [(4'hd):(1'h0)] wire943;
  assign y = {wire960,
                 wire959,
                 wire958,
                 wire957,
                 wire956,
                 wire955,
                 wire953,
                 wire952,
                 wire951,
                 wire950,
                 wire949,
                 wire948,
                 wire947,
                 wire946,
                 wire945,
                 wire943,
                 (1'h0)};
  module12 modinst944 (wire943, clk, wire10, wire11, wire8, wire9);
  assign wire945 = ((wire11[(2'h2):(1'h0)] ~^ (wire943[(3'h5):(2'h3)] ?
                       $signed((wire10 & wire8)) : ((wire8 ? (8'h9c) : wire8) ?
                           $signed(wire943) : $signed((8'ha7))))) == ({(~|$signed(wire8)),
                           $unsigned({wire9, wire9})} ?
                       (~^$signed(wire10)) : (~^$unsigned(wire11[(4'hf):(4'ha)]))));
  assign wire946 = wire943;
  assign wire947 = ($unsigned(($signed($signed((7'h42))) ?
                           wire946 : (~^$signed((8'hbc))))) ?
                       ((8'ha0) ?
                           (((wire946 ? wire943 : wire943) * {(8'hac),
                               wire11}) <<< (wire9 < {wire945,
                               wire946})) : $signed(wire946[(3'h4):(1'h0)])) : ((-(~|(wire946 ~^ wire8))) ?
                           wire943[(2'h3):(2'h2)] : $unsigned(($signed(wire943) & {wire10}))));
  assign wire948 = wire11;
  assign wire949 = $unsigned($signed(($signed($signed((8'ha9))) == {(wire948 ?
                           wire943 : wire10),
                       $unsigned(wire946)})));
  assign wire950 = (!(((+wire948[(3'h5):(2'h3)]) ?
                           ($unsigned(wire8) ?
                               (8'hbe) : (~^wire949)) : wire949[(3'h7):(2'h3)]) ?
                       {$unsigned($signed(wire945))} : {$unsigned((~&wire946)),
                           (wire948 - (!wire10))}));
  assign wire951 = wire943[(4'ha):(4'ha)];
  assign wire952 = $unsigned(((wire950[(4'ha):(2'h3)] ?
                       $signed((wire10 ?
                           (8'hbc) : wire947)) : $unsigned((+(8'ha6)))) | wire946));
  module479 modinst954 (.y(wire953), .wire481(wire949), .wire482(wire945), .clk(clk), .wire480(wire946), .wire483(wire948));
  assign wire955 = (wire10[(5'h13):(5'h13)] | wire10);
  assign wire956 = (~&((8'hb9) ? $unsigned(wire943[(3'h4):(2'h3)]) : (8'hb7)));
  assign wire957 = wire947[(3'h5):(1'h0)];
  assign wire958 = (~^(wire11[(3'h6):(1'h1)] != (~^($unsigned(wire953) ?
                       {(8'ha2), wire8} : ((7'h43) <= wire950)))));
  assign wire959 = wire950[(4'hd):(1'h1)];
  assign wire960 = (^~wire950);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module12
#( parameter param941 = {(-(!{{(8'hbf)}, ((8'ha9) ? (8'ha6) : (7'h43))}))}
, parameter param942 = (8'h9c) )
(y, clk, wire13, wire14, wire15, wire16);
  output wire [(32'h1d3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire13;
  input wire [(5'h14):(1'h0)] wire14;
  input wire [(5'h15):(1'h0)] wire15;
  input wire signed [(3'h7):(1'h0)] wire16;
  wire signed [(4'ha):(1'h0)] wire940;
  wire [(4'hb):(1'h0)] wire939;
  reg signed [(5'h13):(1'h0)] reg938 = (1'h0);
  reg [(4'hf):(1'h0)] reg937 = (1'h0);
  reg [(4'h8):(1'h0)] reg936 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg935 = (1'h0);
  reg [(2'h2):(1'h0)] reg934 = (1'h0);
  reg [(4'he):(1'h0)] reg933 = (1'h0);
  reg [(4'hb):(1'h0)] reg932 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg931 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg930 = (1'h0);
  reg [(4'hf):(1'h0)] reg929 = (1'h0);
  reg [(5'h13):(1'h0)] reg928 = (1'h0);
  reg [(4'hf):(1'h0)] reg927 = (1'h0);
  reg [(4'hd):(1'h0)] reg926 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg925 = (1'h0);
  reg [(3'h4):(1'h0)] reg924 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg923 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg922 = (1'h0);
  reg [(4'hc):(1'h0)] reg921 = (1'h0);
  wire [(4'hd):(1'h0)] wire920;
  wire signed [(4'hd):(1'h0)] wire919;
  wire [(4'he):(1'h0)] wire918;
  wire [(5'h14):(1'h0)] wire917;
  wire signed [(3'h5):(1'h0)] wire916;
  wire [(5'h12):(1'h0)] wire17;
  wire signed [(5'h15):(1'h0)] wire18;
  wire signed [(5'h12):(1'h0)] wire19;
  wire [(5'h12):(1'h0)] wire20;
  wire signed [(4'hf):(1'h0)] wire413;
  wire signed [(4'hf):(1'h0)] wire640;
  wire signed [(5'h13):(1'h0)] wire642;
  wire signed [(5'h15):(1'h0)] wire643;
  wire signed [(5'h12):(1'h0)] wire644;
  wire [(2'h3):(1'h0)] wire645;
  wire signed [(4'h9):(1'h0)] wire688;
  wire [(3'h7):(1'h0)] wire690;
  wire [(2'h2):(1'h0)] wire914;
  assign y = {wire940,
                 wire939,
                 reg938,
                 reg937,
                 reg936,
                 reg935,
                 reg934,
                 reg933,
                 reg932,
                 reg931,
                 reg930,
                 reg929,
                 reg928,
                 reg927,
                 reg926,
                 reg925,
                 reg924,
                 reg923,
                 reg922,
                 reg921,
                 wire920,
                 wire919,
                 wire918,
                 wire917,
                 wire916,
                 wire17,
                 wire18,
                 wire19,
                 wire20,
                 wire413,
                 wire640,
                 wire642,
                 wire643,
                 wire644,
                 wire645,
                 wire688,
                 wire690,
                 wire914,
                 (1'h0)};
  assign wire17 = $signed(($signed(($signed((8'hbf)) == {wire14})) ~^ $signed((~|{wire16,
                      (8'h9c)}))));
  assign wire18 = wire15;
  assign wire19 = $unsigned($signed(($unsigned((wire17 ~^ wire13)) ^ (7'h44))));
  assign wire20 = $unsigned(((wire15[(5'h15):(4'h8)] ^~ (|$unsigned(wire13))) ?
                      wire16 : $signed((~(wire19 >> wire14)))));
  module21 modinst414 (wire413, clk, wire20, wire14, wire18, wire19);
  module415 modinst641 (.y(wire640), .wire419(wire13), .wire418(wire18), .wire416(wire19), .wire417(wire14), .clk(clk));
  assign wire642 = ({($unsigned($unsigned((8'hb7))) ?
                           wire640[(1'h0):(1'h0)] : wire17[(5'h12):(3'h4)]),
                       (^wire14[(4'hd):(4'hc)])} << wire413);
  assign wire643 = $unsigned($signed(($signed((8'hb8)) ?
                       (~|$unsigned(wire19)) : ({(8'ha0), wire14} ?
                           (wire15 ? wire19 : wire20) : (wire640 <= wire17)))));
  assign wire644 = $unsigned($unsigned($unsigned((wire642 >>> (&(8'ha7))))));
  assign wire645 = ($unsigned((($unsigned(wire17) ?
                           {wire13} : (wire642 != wire642)) ^ $signed((^wire16)))) ?
                       wire14[(5'h12):(5'h12)] : ((~$unsigned((wire15 | wire19))) | wire640));
  module646 modinst689 (wire688, clk, wire644, wire642, wire643, wire13);
  assign wire690 = wire688;
  module691 modinst915 (.wire695(wire644), .clk(clk), .wire694(wire15), .wire696(wire643), .wire693(wire13), .y(wire914), .wire692(wire642));
  assign wire916 = (wire18 && (+$signed((wire15[(2'h2):(1'h0)] | $signed(wire642)))));
  assign wire917 = ((~&wire16) ~^ $unsigned({$unsigned((wire15 && (8'h9d))),
                       ((^(8'h9f)) ? ((8'hb7) | wire18) : $signed(wire688))}));
  assign wire918 = ($unsigned((wire19 ?
                       wire640[(2'h3):(1'h1)] : wire413[(4'h9):(4'h8)])) << {(~(8'hb3))});
  assign wire919 = $signed($unsigned($signed((8'ha1))));
  assign wire920 = wire20;
  always
    @(posedge clk) begin
      if (wire918[(4'hd):(2'h2)])
        begin
          if (wire413)
            begin
              reg921 <= $signed(wire413[(2'h3):(2'h3)]);
              reg922 <= $unsigned((((-(wire16 ^~ wire920)) ?
                      wire690[(3'h7):(3'h6)] : (^~$unsigned(wire15))) ?
                  (8'h9c) : wire916));
              reg923 <= wire916;
              reg924 <= (^~(~^(^~wire16)));
              reg925 <= (~|$signed((reg923[(3'h4):(2'h3)] < {{wire413}})));
            end
          else
            begin
              reg921 <= wire413[(4'hc):(3'h7)];
              reg922 <= (^wire20);
            end
        end
      else
        begin
          if (reg921[(3'h7):(2'h2)])
            begin
              reg921 <= $unsigned($signed(wire644[(4'hf):(2'h2)]));
              reg922 <= ($signed(wire917) && $unsigned(reg921[(1'h1):(1'h0)]));
              reg923 <= reg925;
            end
          else
            begin
              reg921 <= {((-$unsigned(wire17)) == (^~(|{wire640}))),
                  {($signed(wire644) - {reg924,
                          (wire917 ? wire645 : wire413)})}};
              reg922 <= ((~^wire688) ?
                  wire18[(4'hf):(4'he)] : $unsigned((($signed(wire688) + (reg923 ?
                          wire642 : wire644)) ?
                      wire914 : (((8'ha8) & wire20) & reg922[(2'h2):(2'h2)]))));
              reg923 <= wire14;
              reg924 <= (~((|((wire919 <<< (8'ha6)) ^~ (~&wire645))) ~^ reg923));
            end
          reg925 <= ($signed($signed(((&reg924) >>> $signed(wire17)))) ?
              (!((wire16[(3'h7):(1'h1)] ? (~|(8'hb1)) : ((8'ha1) >> wire914)) ?
                  wire13 : ((wire14 ? reg923 : wire19) ?
                      $unsigned(wire917) : {wire919}))) : reg925);
          if ($unsigned(wire20[(3'h6):(1'h0)]))
            begin
              reg926 <= ($signed(({(|wire20), ((7'h40) ? (8'h9f) : wire14)} ?
                  (7'h43) : $signed($unsigned(reg925)))) ^~ (((((8'ha9) ?
                          wire919 : wire14) ?
                      wire919[(4'hb):(4'hb)] : {wire20, reg925}) ?
                  reg921[(4'hb):(3'h4)] : ((wire918 ?
                      wire13 : wire16) && (&(8'ha6)))) > ({wire690[(2'h2):(2'h2)]} <= wire642)));
              reg927 <= $unsigned(((((~|wire643) || (~^(8'ha1))) ?
                  $signed(((7'h42) ? reg922 : wire690)) : ($signed(wire643) ?
                      $signed(wire688) : ((8'hbe) ?
                          wire919 : (8'h9d)))) <<< $signed((wire16 ?
                  (wire916 ? wire16 : wire15) : wire17))));
              reg928 <= ({$unsigned({$signed((8'hb1)), ((8'ha6) & reg923)}),
                  ($signed(reg923) ?
                      ((&wire644) ~^ wire14[(3'h4):(1'h0)]) : wire918)} >= $unsigned((|(reg926[(2'h3):(1'h0)] >> (~&reg921)))));
              reg929 <= $signed((~|$signed(wire690[(1'h0):(1'h0)])));
              reg930 <= (~&(^~wire413));
            end
          else
            begin
              reg926 <= ((!(!wire643[(3'h5):(2'h2)])) >>> $unsigned(wire13[(4'h9):(2'h2)]));
              reg927 <= ((reg921[(4'h9):(4'h8)] + wire643) ?
                  wire918[(1'h0):(1'h0)] : (~{$signed(wire914),
                      (^$signed(wire16))}));
              reg928 <= ((8'h9f) <= wire920[(4'hc):(3'h5)]);
              reg929 <= reg922[(4'ha):(3'h4)];
            end
          reg931 <= {($signed((((8'ha9) ?
                      (8'haf) : wire690) >>> $signed(wire642))) ?
                  {wire20[(4'hb):(3'h6)]} : $unsigned($signed(wire919[(2'h2):(1'h1)]))),
              {(&$signed((wire914 ? (8'h9e) : wire17)))}};
          if (wire413[(4'he):(4'hb)])
            begin
              reg932 <= ((~(&$signed((reg925 == wire640)))) <<< ({{wire643,
                          $signed(wire13)}} ?
                  ((&$signed(wire644)) ?
                      reg922[(4'ha):(3'h7)] : $unsigned($signed(wire914))) : (|(((7'h42) ?
                          wire20 : wire413) ?
                      $unsigned(wire917) : (wire688 << reg923)))));
              reg933 <= ((+wire14[(1'h1):(1'h1)]) ?
                  reg932[(4'h8):(3'h5)] : ($unsigned(($signed(wire14) ?
                      (+wire14) : (wire17 != (8'ha0)))) <= (-(^~$signed(reg927)))));
              reg934 <= wire918;
              reg935 <= ({(($unsigned(reg924) << reg924[(1'h0):(1'h0)]) ?
                          $signed($signed(wire918)) : $signed((|reg929)))} ?
                  wire15[(5'h15):(4'ha)] : (wire914[(1'h1):(1'h0)] ?
                      $unsigned(wire16[(3'h5):(2'h2)]) : (reg930 ?
                          $unsigned($unsigned(wire640)) : reg933[(1'h1):(1'h0)])));
              reg936 <= $unsigned({$unsigned(($unsigned(reg929) <<< $signed(wire917))),
                  ($signed({wire917}) - reg929)});
            end
          else
            begin
              reg932 <= wire640;
              reg933 <= wire920;
              reg934 <= ($signed((reg921[(4'h9):(2'h3)] ?
                  wire916[(3'h4):(2'h2)] : $signed($unsigned(wire15)))) || wire14[(4'ha):(3'h6)]);
              reg935 <= ($unsigned($signed((reg935[(2'h3):(2'h2)] > ((8'hbf) >>> reg930)))) ?
                  ($unsigned((!(&(8'hab)))) - $unsigned((reg933[(4'h8):(3'h5)] ?
                      (reg922 ?
                          reg923 : reg935) : reg923))) : ({$unsigned(reg922),
                      reg927[(4'h9):(3'h7)]} <<< $signed(($unsigned((7'h41)) == wire13[(3'h7):(3'h6)]))));
              reg936 <= wire17[(2'h2):(1'h0)];
            end
        end
      reg937 <= (|reg926[(1'h0):(1'h0)]);
      reg938 <= $signed((wire918 ?
          {(wire918 - ((8'hb9) - reg922)),
              wire916[(1'h0):(1'h0)]} : {$signed($signed(wire643)),
              ({reg929} ? wire15 : $signed(reg935))}));
    end
  assign wire939 = (((!(8'hb2)) <<< ($unsigned(reg938[(3'h4):(2'h2)]) ~^ (-reg930[(1'h1):(1'h1)]))) != ({(&wire645[(2'h3):(1'h0)]),
                       $signed($unsigned(wire642))} >>> (~$signed((wire644 ?
                       (8'h9f) : (7'h40))))));
  assign wire940 = $unsigned((~|$unsigned(((wire14 || wire645) ?
                       (~^wire17) : {wire939}))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module691
#(parameter param913 = {(8'hb6)})
(y, clk, wire696, wire695, wire694, wire693, wire692);
  output wire [(32'h1d5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire696;
  input wire [(5'h12):(1'h0)] wire695;
  input wire [(4'hd):(1'h0)] wire694;
  input wire signed [(2'h2):(1'h0)] wire693;
  input wire signed [(5'h11):(1'h0)] wire692;
  reg signed [(4'ha):(1'h0)] reg912 = (1'h0);
  reg [(4'hb):(1'h0)] reg911 = (1'h0);
  reg [(3'h5):(1'h0)] reg910 = (1'h0);
  reg [(4'hf):(1'h0)] reg909 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg908 = (1'h0);
  reg [(4'hd):(1'h0)] reg907 = (1'h0);
  reg signed [(4'he):(1'h0)] reg906 = (1'h0);
  reg [(5'h15):(1'h0)] reg905 = (1'h0);
  reg [(4'h9):(1'h0)] reg904 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg903 = (1'h0);
  reg [(4'hb):(1'h0)] reg902 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg901 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg900 = (1'h0);
  reg [(5'h11):(1'h0)] reg899 = (1'h0);
  reg signed [(4'he):(1'h0)] reg898 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg897 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg896 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg895 = (1'h0);
  reg [(4'ha):(1'h0)] reg894 = (1'h0);
  reg [(4'h8):(1'h0)] reg893 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg892 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg891 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg890 = (1'h0);
  reg signed [(4'he):(1'h0)] reg889 = (1'h0);
  reg [(4'hc):(1'h0)] reg888 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg887 = (1'h0);
  reg [(4'ha):(1'h0)] reg886 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire885;
  wire signed [(4'he):(1'h0)] wire884;
  wire signed [(3'h5):(1'h0)] wire883;
  wire signed [(4'hc):(1'h0)] wire882;
  wire [(4'h8):(1'h0)] wire880;
  wire [(4'hc):(1'h0)] wire870;
  wire signed [(4'h8):(1'h0)] wire868;
  wire [(5'h13):(1'h0)] wire700;
  wire [(5'h13):(1'h0)] wire699;
  wire [(2'h2):(1'h0)] wire698;
  wire [(5'h14):(1'h0)] wire697;
  assign y = {reg912,
                 reg911,
                 reg910,
                 reg909,
                 reg908,
                 reg907,
                 reg906,
                 reg905,
                 reg904,
                 reg903,
                 reg902,
                 reg901,
                 reg900,
                 reg899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 reg893,
                 reg892,
                 reg891,
                 reg890,
                 reg889,
                 reg888,
                 reg887,
                 reg886,
                 wire885,
                 wire884,
                 wire883,
                 wire882,
                 wire880,
                 wire870,
                 wire868,
                 wire700,
                 wire699,
                 wire698,
                 wire697,
                 (1'h0)};
  assign wire697 = {wire696[(5'h14):(4'hd)],
                       ($unsigned((!wire693)) >= ($signed(((8'hba) ?
                               wire695 : wire693)) ?
                           wire692 : ((wire692 ?
                               wire696 : wire694) | ((8'ha8) >> wire693))))};
  assign wire698 = (&{({wire692} <= wire693),
                       ((~&$signed((8'ha1))) ?
                           $signed({wire697}) : ((~^wire693) ^~ wire695))});
  assign wire699 = $unsigned(({(8'hb8), wire697} ?
                       wire694[(3'h5):(1'h1)] : $signed(($unsigned((8'hba)) ?
                           (-wire697) : (wire697 != wire693)))));
  assign wire700 = $unsigned((wire695 >= wire696[(4'h8):(2'h3)]));
  module701 modinst869 (.wire703(wire697), .wire702(wire696), .clk(clk), .wire704(wire700), .wire705(wire692), .y(wire868));
  assign wire870 = {$unsigned($unsigned((~^$signed(wire699)))),
                       ($signed((!wire698)) ?
                           {$unsigned((&wire696)), wire868} : wire699)};
  module871 modinst881 (.clk(clk), .wire874(wire696), .y(wire880), .wire875(wire700), .wire872(wire695), .wire873(wire870));
  assign wire882 = ((wire699 ?
                       (!(|{wire868,
                           wire696})) : (($signed(wire699) << $unsigned(wire696)) ?
                           $signed((wire694 != (8'hb1))) : $unsigned(wire693[(1'h1):(1'h1)]))) & $unsigned($unsigned((-wire698[(1'h1):(1'h1)]))));
  assign wire883 = (wire870 && $signed(wire698));
  assign wire884 = {{wire698[(1'h0):(1'h0)]}};
  assign wire885 = wire698;
  always
    @(posedge clk) begin
      reg886 <= $signed((^~(wire695[(5'h10):(4'hd)] ?
          $unsigned((wire698 ^~ wire693)) : ({wire695, wire885} ?
              $signed(wire697) : $unsigned((8'hb2))))));
      if ({($signed((wire880 ? $unsigned(wire692) : wire698)) ?
              $unsigned($unsigned((wire699 ?
                  (8'hb4) : wire697))) : $signed((^wire695))),
          $signed((-wire882[(4'h9):(3'h4)]))})
        begin
          if (wire693[(1'h0):(1'h0)])
            begin
              reg887 <= ($unsigned(((!{wire695}) ?
                  ($unsigned(wire882) >> $unsigned(reg886)) : wire695[(4'hc):(2'h3)])) <= $signed($signed((-(|wire884)))));
              reg888 <= $unsigned((+wire700));
              reg889 <= ($signed(wire882[(4'h8):(1'h0)]) >>> $signed({$unsigned(wire697[(3'h7):(1'h0)]),
                  wire883[(3'h5):(3'h4)]}));
              reg890 <= reg889;
              reg891 <= wire880[(1'h1):(1'h1)];
            end
          else
            begin
              reg887 <= $unsigned(((|((&(8'hac)) ?
                      (8'h9f) : $unsigned(wire883))) ?
                  (~wire696[(3'h5):(3'h5)]) : ($signed($signed(wire880)) ?
                      (-(+reg887)) : wire693)));
              reg888 <= wire885;
              reg889 <= ((|({(&reg887)} ^ ((reg890 & wire883) ?
                  (wire880 ?
                      (8'hb9) : reg889) : $unsigned(wire700)))) ~^ $unsigned((|{$unsigned(wire692)})));
            end
          reg892 <= $unsigned($unsigned(wire880[(1'h1):(1'h0)]));
          reg893 <= $unsigned(wire697);
          if ($unsigned($unsigned((~&reg886))))
            begin
              reg894 <= wire698;
            end
          else
            begin
              reg894 <= (($signed((wire883[(2'h2):(2'h2)] << reg887)) ?
                      $unsigned($signed((wire700 - wire697))) : wire692[(2'h2):(1'h1)]) ?
                  $signed((|wire698)) : (~|{(wire870[(1'h0):(1'h0)] << (8'ha9)),
                      (reg894[(3'h5):(3'h5)] ?
                          reg887[(3'h4):(1'h0)] : {reg887})}));
              reg895 <= (!((-$signed($unsigned(reg891))) <<< {((wire696 ?
                          wire885 : wire880) ?
                      (wire883 ? (8'hae) : wire868) : reg893[(2'h3):(1'h1)])}));
              reg896 <= (reg895[(4'ha):(4'h9)] ?
                  (|wire699) : reg892[(2'h3):(2'h3)]);
              reg897 <= (|$unsigned($signed($signed($unsigned(wire884)))));
            end
          if (reg894[(1'h1):(1'h1)])
            begin
              reg898 <= $signed(wire698[(2'h2):(1'h0)]);
              reg899 <= reg888[(2'h2):(1'h0)];
              reg900 <= $unsigned((8'hbd));
              reg901 <= ($signed(reg894) ?
                  (8'hb4) : (~^$signed($unsigned(((8'hb9) == wire880)))));
              reg902 <= (reg889[(4'hc):(1'h0)] ? $unsigned((8'ha3)) : wire692);
            end
          else
            begin
              reg898 <= $signed(((~^reg902) > reg901));
              reg899 <= wire884;
              reg900 <= wire697[(3'h6):(1'h0)];
              reg901 <= (~wire883[(1'h1):(1'h1)]);
              reg902 <= (wire883 <= wire699[(3'h5):(3'h5)]);
            end
        end
      else
        begin
          reg887 <= ($unsigned($unsigned(((reg890 ~^ reg902) ?
                  {wire699} : $unsigned(wire697)))) ?
              $unsigned(reg890) : reg891[(2'h2):(1'h1)]);
          reg888 <= wire885;
          reg889 <= (|$unsigned($unsigned((~(wire693 >= wire693)))));
          reg890 <= (7'h40);
        end
      if ((wire693[(1'h1):(1'h0)] ?
          $signed({reg901}) : (reg886 ^~ $unsigned(wire692))))
        begin
          if (reg895)
            begin
              reg903 <= (~|{(wire882 * ({wire695} || wire870[(4'h8):(4'h8)]))});
              reg904 <= (($signed({reg902, (8'haf)}) ? reg889 : wire883) ?
                  wire700[(2'h2):(1'h0)] : ($signed($unsigned(((8'hae) ?
                      reg898 : wire695))) && (8'hb7)));
              reg905 <= wire883;
            end
          else
            begin
              reg903 <= (!((8'hae) == $signed($unsigned((wire868 ?
                  (8'hba) : reg896)))));
              reg904 <= $unsigned((($signed(reg904) && (|{wire692})) ?
                  {{$signed(reg895)}} : (~|((reg900 ~^ (8'hbc)) | wire698[(1'h0):(1'h0)]))));
              reg905 <= ((reg904 ?
                  ((wire870 ? (7'h43) : $signed(wire883)) ?
                      $signed(((8'hb0) ? wire692 : reg896)) : {reg903,
                          wire870[(4'hb):(3'h6)]}) : reg905[(5'h15):(5'h14)]) != wire883[(3'h4):(1'h1)]);
              reg906 <= $unsigned(reg900);
            end
          reg907 <= (wire882 ?
              (^~$signed($signed((reg899 ?
                  (8'hb1) : (8'hab))))) : ({reg903[(1'h1):(1'h1)],
                      ($signed(wire698) & (wire870 ? reg892 : (8'ha2)))} ?
                  ((reg903 ? $unsigned(wire882) : (+wire695)) ?
                      $unsigned({reg906}) : (&reg901)) : ((8'hba) <= (8'hbd))));
        end
      else
        begin
          reg903 <= (~^(~$unsigned(($unsigned(reg890) >> (wire694 ?
              wire884 : reg896)))));
          if ((wire697 ?
              $signed({$signed((&wire694))}) : (reg896 ?
                  $unsigned({(8'hbc),
                      (reg894 && reg896)}) : (^~{$unsigned((8'hab)),
                      $unsigned(wire698)}))))
            begin
              reg904 <= $unsigned(($unsigned((reg893 ?
                      $signed(reg887) : {wire884, wire884})) ?
                  reg903 : $unsigned($signed((wire884 >= reg896)))));
              reg905 <= $unsigned($unsigned(reg896));
              reg906 <= (reg904[(3'h5):(2'h3)] ?
                  {$unsigned($unsigned(wire699))} : $unsigned({$signed($unsigned((7'h40))),
                      wire882[(4'ha):(1'h1)]}));
              reg907 <= ($signed(wire692) <= $signed($unsigned($unsigned({reg907}))));
              reg908 <= $signed($signed(reg906));
            end
          else
            begin
              reg904 <= {$unsigned({reg903}),
                  $signed($unsigned($unsigned(reg889[(3'h5):(2'h2)])))};
              reg905 <= reg897;
              reg906 <= (^{{reg886[(3'h5):(2'h3)]},
                  {$signed(reg888[(3'h5):(1'h0)]),
                      (reg890[(3'h4):(1'h1)] ?
                          {(8'hbc), wire700} : $signed(reg905))}});
              reg907 <= wire882[(1'h0):(1'h0)];
              reg908 <= $unsigned((-(((~wire697) == (wire693 && reg890)) ?
                  ((8'hae) ^~ (reg899 == reg892)) : ((wire884 <<< wire883) && $signed(reg902)))));
            end
          if ((8'hb9))
            begin
              reg909 <= (~$signed($signed({reg900[(5'h11):(4'he)],
                  $unsigned(wire698)})));
              reg910 <= wire880;
            end
          else
            begin
              reg909 <= reg894[(1'h0):(1'h0)];
              reg910 <= {((((reg888 < reg902) >>> $signed(wire700)) ?
                      reg898[(4'hc):(2'h2)] : ((wire695 != wire693) | (+(8'hb1)))) - $signed($unsigned(reg888)))};
              reg911 <= {{{{{reg898}},
                          (reg902[(4'h8):(3'h5)] ~^ $unsigned(reg908))}}};
            end
          reg912 <= ($signed(((-$signed((8'hac))) ?
                  (&$signed(reg898)) : (^(^wire883)))) ?
              reg910[(1'h1):(1'h1)] : wire884[(4'h8):(3'h5)]);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module646
#( parameter param686 = {((^(((8'hb3) * (8'hb7)) ? ((8'h9e) >>> (8'hb3)) : (8'h9e))) <<< ((-((8'ha6) ^ (8'hab))) != {((8'hb4) << (8'ha3))}))}
, parameter param687 = param686 )
(y, clk, wire650, wire649, wire648, wire647);
  output wire [(32'h110):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire650;
  input wire [(5'h13):(1'h0)] wire649;
  input wire [(4'hb):(1'h0)] wire648;
  input wire signed [(4'h9):(1'h0)] wire647;
  wire [(3'h4):(1'h0)] wire685;
  wire [(4'hc):(1'h0)] wire684;
  reg [(5'h10):(1'h0)] reg683 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg682 = (1'h0);
  reg [(4'h9):(1'h0)] reg681 = (1'h0);
  reg [(4'h9):(1'h0)] reg680 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg679 = (1'h0);
  reg [(5'h10):(1'h0)] reg678 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire677;
  wire [(3'h7):(1'h0)] wire676;
  wire signed [(3'h7):(1'h0)] wire674;
  reg [(5'h14):(1'h0)] reg662 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg661 = (1'h0);
  reg [(5'h13):(1'h0)] reg660 = (1'h0);
  reg [(4'h9):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg658 = (1'h0);
  reg [(4'he):(1'h0)] reg657 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg656 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg655 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg654 = (1'h0);
  reg [(5'h12):(1'h0)] reg653 = (1'h0);
  wire [(4'hb):(1'h0)] wire652;
  wire [(3'h5):(1'h0)] wire651;
  assign y = {wire685,
                 wire684,
                 reg683,
                 reg682,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 wire677,
                 wire676,
                 wire674,
                 reg662,
                 reg661,
                 reg660,
                 reg659,
                 reg658,
                 reg657,
                 reg656,
                 reg655,
                 reg654,
                 reg653,
                 wire652,
                 wire651,
                 (1'h0)};
  assign wire651 = $signed({wire647, wire650});
  assign wire652 = ((((-{wire650}) ^~ wire651[(2'h3):(2'h3)]) ?
                       wire649[(5'h11):(4'hc)] : ($signed((wire650 ^ wire649)) ?
                           ((wire648 >>> wire648) - {wire650,
                               wire651}) : wire648[(2'h3):(1'h0)])) == wire649);
  always
    @(posedge clk) begin
      if (wire649[(3'h7):(3'h7)])
        begin
          reg653 <= wire651[(1'h0):(1'h0)];
          if ($unsigned($unsigned((((~reg653) ^ (~|wire648)) & $signed((wire650 >> (8'ha8)))))))
            begin
              reg654 <= (($signed({reg653[(1'h0):(1'h0)]}) ^ wire649) >>> (|(^wire651)));
              reg655 <= ((&wire649[(5'h11):(2'h3)]) ^~ ($signed(((^wire647) > wire650)) ?
                  wire650[(1'h1):(1'h0)] : {wire648[(1'h0):(1'h0)], wire648}));
            end
          else
            begin
              reg654 <= (wire651 ?
                  (~{wire647[(2'h3):(2'h2)]}) : (&(wire649 ?
                      wire652 : ($signed(reg653) ?
                          (wire649 ? wire650 : wire651) : $signed(wire650)))));
              reg655 <= (~|reg653);
              reg656 <= $unsigned($signed((^~$unsigned(reg654))));
              reg657 <= (wire651 ?
                  $unsigned(reg653) : ((~|$unsigned(reg655)) && (reg653 < $signed($unsigned((8'hbb))))));
            end
          reg658 <= reg656;
          if (reg655)
            begin
              reg659 <= wire648;
              reg660 <= (^$unsigned((7'h43)));
              reg661 <= (&$signed((^wire652[(4'ha):(4'h9)])));
            end
          else
            begin
              reg659 <= ((wire648[(1'h0):(1'h0)] >>> (~&(~|reg656))) | (^~wire652));
              reg660 <= ($unsigned(wire648) ?
                  wire650 : (reg653 ?
                      $unsigned($signed(reg656[(2'h2):(1'h1)])) : ({(reg661 ?
                                  reg653 : reg656)} ?
                          (reg659[(2'h3):(2'h3)] ^~ (wire647 ?
                              wire651 : reg657)) : (wire650 || (reg656 | reg660)))));
              reg661 <= ({(~^wire652),
                  ({$unsigned(reg660)} ?
                      $unsigned($signed((8'ha8))) : $signed(((8'hb5) ~^ wire648)))} <= (!(|{reg658,
                  $signed(wire648)})));
            end
          reg662 <= wire648;
        end
      else
        begin
          reg653 <= $signed((~|reg658[(4'ha):(3'h6)]));
          reg654 <= wire651[(3'h5):(1'h0)];
          if ((($unsigned(reg655[(3'h5):(1'h1)]) ?
                  (~^(8'ha2)) : (!({(8'h9c), (8'ha5)} != $signed(reg654)))) ?
              {wire647,
                  $unsigned($unsigned(reg656[(5'h11):(3'h7)]))} : $signed(wire649)))
            begin
              reg655 <= $signed(reg659);
              reg656 <= $unsigned(reg660[(4'ha):(3'h7)]);
            end
          else
            begin
              reg655 <= $signed($unsigned(wire651[(2'h2):(2'h2)]));
            end
          reg657 <= $unsigned((~^(wire647[(3'h4):(1'h0)] || (&(!wire651)))));
          reg658 <= $signed(reg659[(3'h5):(2'h2)]);
        end
    end
  module663 modinst675 (.wire666(wire652), .y(wire674), .clk(clk), .wire665(wire647), .wire667(reg656), .wire664(reg660));
  assign wire676 = $unsigned(((reg657 ?
                           $unsigned(reg657) : (reg654 ?
                               wire648[(3'h4):(1'h0)] : wire651)) ?
                       wire652[(3'h7):(3'h7)] : (reg661[(2'h2):(1'h0)] <= $signed(wire650[(1'h0):(1'h0)]))));
  assign wire677 = reg662;
  always
    @(posedge clk) begin
      if ((+$unsigned((((wire677 ?
          reg658 : reg656) > wire650) * $unsigned(wire650[(1'h1):(1'h1)])))))
        begin
          reg678 <= (reg662 ?
              reg653[(5'h10):(4'hb)] : (($signed((reg653 * wire651)) ^ (-reg659)) ?
                  wire648[(4'h9):(4'h9)] : (((~|reg656) ?
                      $unsigned(wire676) : (reg656 <<< reg658)) | (reg655 ^~ $signed(wire650)))));
          reg679 <= reg662;
          if ((($unsigned($unsigned((8'hb9))) ?
                  $unsigned($unsigned($signed(reg659))) : ((~|$unsigned(reg653)) ?
                      wire649 : (wire650[(1'h0):(1'h0)] || $unsigned(wire652)))) ?
              ($signed(($unsigned(wire651) ? reg660 : (^reg659))) ?
                  $unsigned(((~^(8'ha2)) ?
                      reg658 : $unsigned(reg659))) : $signed(reg654[(1'h1):(1'h1)])) : $signed(wire651)))
            begin
              reg680 <= (8'hae);
              reg681 <= reg656;
              reg682 <= reg656[(2'h3):(1'h0)];
            end
          else
            begin
              reg680 <= reg681;
              reg681 <= $signed((+($unsigned($unsigned(wire648)) ?
                  wire649[(4'hb):(3'h4)] : (wire651[(1'h0):(1'h0)] ?
                      reg655[(3'h5):(1'h1)] : (|reg680)))));
            end
        end
      else
        begin
          reg678 <= ((+(~&{reg655})) ?
              {(|wire651[(1'h1):(1'h1)]), wire677} : ({{((8'hb0) << wire647),
                          ((8'hb7) >> reg679)},
                      $unsigned((reg678 || reg659))} ?
                  (reg680[(1'h1):(1'h1)] < wire647[(2'h3):(1'h0)]) : ((~^$unsigned(wire677)) + $unsigned(reg661[(1'h0):(1'h0)]))));
        end
      reg683 <= $signed($signed($signed((+((8'hb5) ? (7'h44) : wire652)))));
    end
  assign wire684 = ((reg660 ?
                           (reg657 ^ (wire650[(2'h2):(2'h2)] ^ (reg653 ?
                               (8'hb5) : wire651))) : {{$unsigned((8'h9f))}}) ?
                       $unsigned(reg659[(4'h8):(3'h6)]) : $signed(reg658));
  assign wire685 = $signed((~&(({wire650} >>> $signed(wire649)) ?
                       wire650[(2'h2):(2'h2)] : $unsigned((reg657 > reg680)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module415  (y, clk, wire419, wire418, wire417, wire416);
  output wire [(32'h107):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire419;
  input wire signed [(5'h14):(1'h0)] wire418;
  input wire [(4'hd):(1'h0)] wire417;
  input wire signed [(4'hd):(1'h0)] wire416;
  reg [(4'h8):(1'h0)] reg639 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg638 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg637 = (1'h0);
  reg [(3'h6):(1'h0)] reg636 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg635 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg634 = (1'h0);
  reg [(5'h14):(1'h0)] reg633 = (1'h0);
  reg [(4'he):(1'h0)] reg632 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg631 = (1'h0);
  reg [(5'h13):(1'h0)] reg630 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg629 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg628 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg627 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg626 = (1'h0);
  reg [(4'h9):(1'h0)] reg625 = (1'h0);
  reg [(5'h14):(1'h0)] reg624 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg623 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg622 = (1'h0);
  reg [(2'h3):(1'h0)] reg621 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire620;
  wire signed [(4'ha):(1'h0)] wire619;
  wire [(5'h13):(1'h0)] wire618;
  wire [(4'h9):(1'h0)] wire617;
  wire signed [(3'h7):(1'h0)] wire616;
  wire [(4'h8):(1'h0)] wire614;
  assign y = {reg639,
                 reg638,
                 reg637,
                 reg636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 reg621,
                 wire620,
                 wire619,
                 wire618,
                 wire617,
                 wire616,
                 wire614,
                 (1'h0)};
  module420 modinst615 (.wire421((8'hbb)), .wire425(wire419), .clk(clk), .y(wire614), .wire423(wire418), .wire422(wire416), .wire424(wire417));
  assign wire616 = (($signed($unsigned(wire419)) ?
                       $unsigned((^~wire614)) : wire416[(3'h5):(3'h5)]) & wire419);
  assign wire617 = ($signed($unsigned(wire419)) ?
                       (-wire416[(4'hd):(1'h1)]) : (!$unsigned(wire416[(1'h1):(1'h0)])));
  assign wire618 = ($unsigned($signed(((^wire418) ?
                           {wire616, wire614} : {wire417, (8'ha8)}))) ?
                       ($signed(wire418) * $signed($unsigned($signed(wire614)))) : (|($signed($unsigned((8'ha9))) ?
                           $signed($unsigned(wire419)) : ($unsigned(wire616) ?
                               $unsigned(wire614) : (+wire614)))));
  assign wire619 = wire417[(3'h5):(1'h1)];
  assign wire620 = wire619;
  always
    @(posedge clk) begin
      reg621 <= (|$signed(wire620));
      reg622 <= ((~&(wire417[(3'h7):(2'h2)] | ($unsigned(wire416) ?
              (wire617 | reg621) : wire616[(2'h2):(1'h0)]))) ?
          {((+$unsigned(wire616)) ?
                  wire417[(4'hb):(4'h9)] : wire416[(3'h7):(3'h7)]),
              $unsigned(wire417)} : $signed(wire620[(1'h0):(1'h0)]));
      if ((((reg622 - ((wire619 ? reg622 : wire418) <= $signed(wire417))) ?
              wire416 : $unsigned((reg622 ?
                  ((8'hbc) ? wire416 : wire418) : (wire416 || wire416)))) ?
          ($unsigned(($unsigned(wire620) != wire418)) > (reg621 & ({wire618,
                  wire620} ?
              $unsigned((8'hba)) : wire620))) : (8'hb9)))
        begin
          if (wire619[(2'h2):(2'h2)])
            begin
              reg623 <= (+(-{(wire620[(1'h1):(1'h0)] ?
                      reg621 : wire418[(4'hd):(3'h6)]),
                  $signed(wire614[(3'h4):(1'h1)])}));
              reg624 <= $unsigned(((wire620 << ({(8'haa), reg623} > (wire618 ?
                  reg621 : wire618))) > $unsigned($signed($signed(wire418)))));
              reg625 <= $unsigned(reg621);
              reg626 <= wire418;
              reg627 <= $unsigned(((^~wire614[(1'h1):(1'h1)]) ?
                  $unsigned(wire614[(3'h4):(1'h0)]) : $unsigned({(wire620 <<< reg622)})));
            end
          else
            begin
              reg623 <= $signed($signed({(|((8'ha3) ? wire616 : reg622))}));
              reg624 <= (~|(reg626[(2'h2):(1'h0)] < reg622[(1'h1):(1'h1)]));
            end
          reg628 <= wire620[(3'h5):(1'h1)];
          if ((~^(~wire419[(5'h11):(1'h0)])))
            begin
              reg629 <= (8'h9f);
              reg630 <= $signed((|(|{$signed((8'ha4))})));
              reg631 <= (~$unsigned((~^(~|{wire418}))));
              reg632 <= {(-(^~$signed((~^(8'ha7))))),
                  ((wire419[(4'h8):(2'h3)] << wire417[(4'hd):(1'h1)]) >>> wire419[(3'h4):(2'h3)])};
            end
          else
            begin
              reg629 <= $unsigned($signed(($unsigned((^wire416)) ?
                  (8'hae) : reg624[(2'h2):(1'h1)])));
              reg630 <= (((^(wire618 < $signed(reg621))) ?
                      wire418 : $unsigned($unsigned($unsigned(reg624)))) ?
                  reg627[(2'h2):(1'h0)] : (~($unsigned(reg632[(4'h8):(3'h5)]) ?
                      reg621[(1'h1):(1'h0)] : reg622)));
            end
          reg633 <= ($unsigned((&$signed($unsigned(reg627)))) <= reg632[(1'h1):(1'h0)]);
          if (((8'hbe) || ((($signed(wire614) * (-reg623)) ?
                  reg628[(1'h1):(1'h0)] : $unsigned((~&wire618))) ?
              wire619 : (~($unsigned(reg632) || {reg627})))))
            begin
              reg634 <= (~&(!reg622));
              reg635 <= {wire618[(5'h12):(1'h0)]};
              reg636 <= $unsigned(($unsigned($unsigned((reg631 ?
                  reg623 : reg621))) > (((8'h9c) ?
                  wire616[(3'h7):(1'h1)] : reg624[(4'hf):(4'hd)]) == $signed((^~wire416)))));
              reg637 <= ($signed($signed({(wire618 ? reg634 : reg628),
                  (reg636 || (8'hb3))})) >> $unsigned(wire616[(3'h7):(3'h6)]));
            end
          else
            begin
              reg634 <= reg633[(5'h10):(4'hf)];
              reg635 <= (-$signed($unsigned(wire417[(4'hb):(4'h9)])));
            end
        end
      else
        begin
          reg623 <= ($signed((8'hb4)) ? (8'hab) : reg627);
          reg624 <= ($signed({$unsigned((reg630 ? reg626 : reg630))}) ?
              ((reg625[(1'h1):(1'h0)] < (((8'hab) >>> reg621) & (wire617 >> reg628))) < ((~$unsigned(wire616)) ?
                  $signed($signed(wire617)) : $unsigned((&reg627)))) : ({reg632[(4'h9):(2'h3)],
                  $unsigned((reg626 ?
                      (7'h43) : reg629))} + {$signed((&wire416)),
                  ($signed(reg637) | $unsigned((8'ha0)))}));
          if ((reg631[(2'h3):(2'h2)] << $signed($unsigned(((+reg627) && (wire614 >= wire616))))))
            begin
              reg625 <= wire616;
              reg626 <= wire416;
              reg627 <= reg636;
            end
          else
            begin
              reg625 <= $signed($unsigned(wire619[(1'h0):(1'h0)]));
              reg626 <= ((^~(~|(^$unsigned(reg627)))) ?
                  $signed($signed($unsigned((reg621 ?
                      wire616 : reg627)))) : (reg632[(2'h2):(2'h2)] ?
                      ((~^{reg621}) >> $unsigned((|wire418))) : $signed($unsigned((~^(7'h44))))));
            end
        end
      reg638 <= $signed(($signed($unsigned((~&wire416))) > (|((reg625 ?
          wire620 : reg630) >>> (wire419 <<< (8'hac))))));
      reg639 <= {$unsigned($signed($unsigned(reg625[(2'h3):(1'h0)]))),
          {wire417[(1'h0):(1'h0)],
              ($signed($unsigned(wire614)) ~^ wire416[(1'h0):(1'h0)])}};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module21  (y, clk, wire25, wire24, wire23, wire22);
  output wire [(32'h102):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire25;
  input wire [(5'h13):(1'h0)] wire24;
  input wire signed [(5'h14):(1'h0)] wire23;
  input wire signed [(4'hc):(1'h0)] wire22;
  wire [(5'h15):(1'h0)] wire412;
  wire [(3'h5):(1'h0)] wire411;
  wire [(3'h6):(1'h0)] wire410;
  wire [(5'h10):(1'h0)] wire409;
  wire signed [(4'hd):(1'h0)] wire408;
  wire signed [(4'hf):(1'h0)] wire407;
  wire signed [(4'hc):(1'h0)] wire323;
  wire [(5'h14):(1'h0)] wire189;
  wire signed [(2'h2):(1'h0)] wire187;
  wire signed [(4'h9):(1'h0)] wire28;
  wire signed [(5'h11):(1'h0)] wire27;
  wire [(5'h13):(1'h0)] wire26;
  wire [(4'hd):(1'h0)] wire325;
  wire signed [(3'h5):(1'h0)] wire326;
  wire [(4'h8):(1'h0)] wire327;
  wire [(4'hb):(1'h0)] wire328;
  wire [(5'h15):(1'h0)] wire329;
  wire signed [(5'h15):(1'h0)] wire330;
  wire signed [(5'h10):(1'h0)] wire331;
  wire signed [(3'h7):(1'h0)] wire405;
  assign y = {wire412,
                 wire411,
                 wire410,
                 wire409,
                 wire408,
                 wire407,
                 wire323,
                 wire189,
                 wire187,
                 wire28,
                 wire27,
                 wire26,
                 wire325,
                 wire326,
                 wire327,
                 wire328,
                 wire329,
                 wire330,
                 wire331,
                 wire405,
                 (1'h0)};
  assign wire26 = wire25;
  assign wire27 = wire25;
  assign wire28 = $unsigned(($signed(wire24) ~^ wire27));
  module29 modinst188 (.wire32(wire23), .wire30(wire27), .clk(clk), .wire33(wire26), .wire31(wire24), .y(wire187));
  assign wire189 = (((8'hbc) >>> $signed(wire23)) || wire28[(3'h4):(1'h1)]);
  module190 modinst324 (wire323, clk, wire23, wire27, wire189, wire26, wire22);
  assign wire325 = $signed((~^(wire187 ? wire323 : (~wire189[(4'h9):(3'h5)]))));
  assign wire326 = ((((8'ha1) ? wire25 : $unsigned((wire189 != wire24))) ?
                           (+(~&((8'ha0) >> wire27))) : wire26[(3'h7):(2'h2)]) ?
                       wire23 : $signed(((~(|wire28)) ?
                           $signed({wire187,
                               (8'hbc)}) : (!wire26[(4'he):(1'h0)]))));
  assign wire327 = ($unsigned($unsigned(wire187[(1'h0):(1'h0)])) ^~ $unsigned($signed((wire25 ?
                       (wire22 ~^ (8'had)) : $signed((8'ha9))))));
  assign wire328 = {wire22};
  assign wire329 = ($unsigned($unsigned({$signed(wire189),
                       (^~wire27)})) > wire28[(3'h5):(1'h0)]);
  assign wire330 = wire328;
  assign wire331 = {{(wire28[(3'h4):(1'h0)] ?
                               $unsigned(wire326[(2'h2):(2'h2)]) : wire323[(3'h7):(3'h5)])},
                       wire28[(4'h9):(2'h3)]};
  module332 modinst406 (wire405, clk, wire27, wire331, wire28, wire189, wire329);
  assign wire407 = (wire325[(3'h4):(1'h1)] ?
                       wire189 : (|($unsigned((wire187 ? wire187 : wire326)) ?
                           wire27[(1'h0):(1'h0)] : ((wire28 ?
                                   wire26 : (8'hae)) ?
                               $unsigned(wire23) : $signed((8'ha2))))));
  assign wire408 = ((wire24 || wire331[(3'h4):(2'h3)]) ~^ wire25);
  assign wire409 = $signed($unsigned($unsigned((wire326[(2'h3):(2'h2)] >= wire327))));
  assign wire410 = $signed($signed(wire331));
  assign wire411 = {wire323,
                       ({$signed($signed(wire410)), wire22} != (((~&wire24) ?
                               wire330 : (-wire326)) ?
                           (wire330[(4'h9):(4'h8)] ~^ wire28) : $signed({wire331,
                               wire410})))};
  assign wire412 = {$signed($unsigned(($signed(wire328) > {(8'hbf), wire23}))),
                       $signed(($unsigned((|wire323)) != {$signed(wire22),
                           $signed((8'ha6))}))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module332  (y, clk, wire337, wire336, wire335, wire334, wire333);
  output wire [(32'hfe):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire337;
  input wire [(3'h6):(1'h0)] wire336;
  input wire signed [(4'h9):(1'h0)] wire335;
  input wire [(3'h7):(1'h0)] wire334;
  input wire [(5'h15):(1'h0)] wire333;
  reg [(3'h4):(1'h0)] reg404 = (1'h0);
  reg [(2'h3):(1'h0)] reg403 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg402 = (1'h0);
  reg [(5'h10):(1'h0)] reg401 = (1'h0);
  reg [(4'hd):(1'h0)] reg400 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg399 = (1'h0);
  reg [(3'h6):(1'h0)] reg398 = (1'h0);
  reg [(4'hf):(1'h0)] reg397 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg396 = (1'h0);
  reg signed [(4'he):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg394 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg393 = (1'h0);
  reg [(5'h10):(1'h0)] reg392 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire391;
  wire signed [(2'h3):(1'h0)] wire390;
  wire [(4'h8):(1'h0)] wire388;
  wire [(5'h12):(1'h0)] wire345;
  wire [(4'hc):(1'h0)] wire344;
  wire signed [(5'h11):(1'h0)] wire343;
  wire [(4'ha):(1'h0)] wire342;
  wire [(3'h5):(1'h0)] wire341;
  wire signed [(4'he):(1'h0)] wire340;
  wire [(2'h2):(1'h0)] wire339;
  wire [(5'h12):(1'h0)] wire338;
  assign y = {reg404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 wire391,
                 wire390,
                 wire388,
                 wire345,
                 wire344,
                 wire343,
                 wire342,
                 wire341,
                 wire340,
                 wire339,
                 wire338,
                 (1'h0)};
  assign wire338 = {(^~$signed((wire333 ^ (^~wire334))))};
  assign wire339 = (((wire333[(4'h8):(4'h8)] != wire333) ?
                           wire337 : (((wire333 | wire335) ?
                                   wire333[(5'h10):(5'h10)] : wire338[(3'h7):(3'h7)]) ?
                               (|(8'hb8)) : ((wire337 ?
                                   wire338 : wire335) ^~ wire337))) ?
                       {$unsigned(($signed((8'hbe)) + $signed(wire336)))} : (wire338 <= ($unsigned((wire335 ?
                           wire333 : wire333)) != wire337)));
  assign wire340 = wire336[(3'h5):(1'h0)];
  assign wire341 = (wire336 != (wire334 || {{(wire339 ? wire338 : (8'hb4))},
                       wire334}));
  assign wire342 = (7'h41);
  assign wire343 = $signed(wire336[(3'h6):(2'h2)]);
  assign wire344 = ($unsigned((~^(~&(wire335 ?
                       wire340 : wire341)))) << wire339);
  assign wire345 = ($unsigned(wire339) ?
                       $unsigned($unsigned(((wire341 > wire337) < {(8'h9d),
                           wire333}))) : (wire344 ?
                           $signed((-wire339[(2'h2):(1'h0)])) : ((&(~(8'haa))) ?
                               wire340[(1'h1):(1'h0)] : (wire338 ?
                                   $unsigned(wire337) : (-wire333)))));
  module346 modinst389 (.y(wire388), .clk(clk), .wire347(wire333), .wire350(wire345), .wire349(wire342), .wire348(wire338));
  assign wire390 = (($unsigned(($unsigned(wire334) ?
                           $unsigned(wire388) : (+wire388))) << $signed(wire334[(3'h4):(1'h0)])) ?
                       wire334[(3'h7):(3'h6)] : $unsigned($signed((wire343 ?
                           (wire334 ? wire339 : wire333) : (~wire339)))));
  assign wire391 = ($signed((((wire340 << wire342) ?
                           (wire334 ? wire345 : wire339) : (~&wire337)) ?
                       wire388[(2'h3):(1'h0)] : $unsigned(wire339))) & ((((wire339 >> wire337) ?
                           {wire333,
                               wire335} : (wire345 & wire388)) ^~ (wire390 ?
                           {(8'hba), wire340} : (wire388 * wire334))) ?
                       wire338 : ({(&wire340)} ?
                           (wire343 ?
                               (-wire338) : wire339) : (wire333 & wire345[(4'hd):(1'h1)]))));
  always
    @(posedge clk) begin
      if ($signed({wire388[(3'h7):(3'h4)],
          $signed((+(wire388 ? wire390 : wire336)))}))
        begin
          reg392 <= ((({{wire343}} ?
                  wire337 : $unsigned((wire342 || wire344))) ?
              ($signed(wire390) ?
                  wire338[(4'hb):(1'h0)] : ((&wire391) >> $unsigned(wire340))) : wire338[(5'h10):(4'hf)]) < {$unsigned($signed($unsigned(wire334))),
              $unsigned((+wire339))});
        end
      else
        begin
          if (wire344[(3'h6):(2'h2)])
            begin
              reg392 <= wire342;
            end
          else
            begin
              reg392 <= (+(wire335[(4'h8):(2'h2)] ?
                  ($unsigned($signed(wire339)) * ($unsigned(wire333) ?
                      $signed(wire336) : {wire341})) : {$unsigned((~&wire391))}));
              reg393 <= (~^reg392);
              reg394 <= $unsigned({$signed(((wire338 ?
                      wire345 : (7'h43)) >>> (8'hba)))});
              reg395 <= ($unsigned((($unsigned(wire340) ?
                  {(8'hbb)} : $unsigned(wire345)) >= {(8'hb7),
                  (wire342 ? reg392 : wire388)})) || wire342);
              reg396 <= (wire340 + ((wire344 < wire338) && (~|$unsigned(wire342))));
            end
        end
      reg397 <= reg392[(1'h1):(1'h1)];
      reg398 <= (wire337[(3'h5):(2'h2)] && (8'hbb));
      if ((-(($signed(wire388) ?
          reg395 : wire343[(2'h2):(2'h2)]) >>> {(~|{(8'ha4)})})))
        begin
          reg399 <= (^$unsigned((~&$unsigned((-wire340)))));
          reg400 <= (wire390 && wire343[(2'h2):(2'h2)]);
          reg401 <= wire337[(4'h8):(1'h1)];
          reg402 <= wire390[(1'h1):(1'h1)];
          reg403 <= (wire335 ?
              $signed(($signed((reg398 != reg393)) >= wire339)) : $unsigned((~|((8'ha4) || (wire340 ?
                  wire342 : wire343)))));
        end
      else
        begin
          reg399 <= $unsigned(reg392[(2'h2):(2'h2)]);
          reg400 <= ((~^($signed((~|wire345)) ?
              {reg396} : reg402)) ^~ reg396[(1'h1):(1'h0)]);
        end
      reg404 <= reg392[(3'h5):(1'h1)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module190  (y, clk, wire195, wire194, wire193, wire192, wire191);
  output wire [(32'h26f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire195;
  input wire signed [(4'h9):(1'h0)] wire194;
  input wire signed [(5'h14):(1'h0)] wire193;
  input wire signed [(5'h13):(1'h0)] wire192;
  input wire [(4'hc):(1'h0)] wire191;
  wire signed [(3'h7):(1'h0)] wire322;
  wire [(5'h12):(1'h0)] wire321;
  wire [(3'h6):(1'h0)] wire320;
  wire [(5'h13):(1'h0)] wire319;
  wire [(4'ha):(1'h0)] wire317;
  wire [(5'h12):(1'h0)] wire238;
  reg signed [(5'h12):(1'h0)] reg237 = (1'h0);
  reg [(4'hc):(1'h0)] reg236 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg235 = (1'h0);
  reg [(4'hf):(1'h0)] reg234 = (1'h0);
  reg [(4'hb):(1'h0)] reg233 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg232 = (1'h0);
  reg [(4'hb):(1'h0)] reg231 = (1'h0);
  reg [(3'h6):(1'h0)] reg230 = (1'h0);
  reg [(3'h7):(1'h0)] reg229 = (1'h0);
  reg [(5'h12):(1'h0)] reg228 = (1'h0);
  wire [(4'h9):(1'h0)] wire227;
  wire signed [(5'h15):(1'h0)] wire226;
  reg signed [(4'h8):(1'h0)] reg225 = (1'h0);
  wire signed [(4'he):(1'h0)] wire224;
  wire [(4'h8):(1'h0)] wire223;
  wire signed [(2'h3):(1'h0)] wire222;
  wire signed [(4'hf):(1'h0)] wire221;
  wire [(4'h9):(1'h0)] wire220;
  reg [(5'h11):(1'h0)] reg219 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg218 = (1'h0);
  reg [(4'he):(1'h0)] reg217 = (1'h0);
  reg [(5'h10):(1'h0)] reg216 = (1'h0);
  reg [(5'h15):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg214 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg213 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg212 = (1'h0);
  reg [(2'h3):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg210 = (1'h0);
  reg [(4'h8):(1'h0)] reg209 = (1'h0);
  reg [(4'ha):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg207 = (1'h0);
  reg [(4'h8):(1'h0)] reg206 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg205 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg204 = (1'h0);
  reg [(4'hf):(1'h0)] reg203 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire202;
  wire [(5'h15):(1'h0)] wire201;
  wire signed [(4'hc):(1'h0)] wire200;
  wire [(4'h8):(1'h0)] wire199;
  wire [(4'ha):(1'h0)] wire198;
  wire signed [(5'h15):(1'h0)] wire197;
  wire signed [(5'h15):(1'h0)] wire196;
  assign y = {wire322,
                 wire321,
                 wire320,
                 wire319,
                 wire317,
                 wire238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 wire227,
                 wire226,
                 reg225,
                 wire224,
                 wire223,
                 wire222,
                 wire221,
                 wire220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 wire202,
                 wire201,
                 wire200,
                 wire199,
                 wire198,
                 wire197,
                 wire196,
                 (1'h0)};
  assign wire196 = (^~wire194[(4'h8):(3'h5)]);
  assign wire197 = {$unsigned($signed((+wire196[(4'hb):(3'h4)]))),
                       (wire196[(4'hb):(4'ha)] ?
                           ((+{wire196, (7'h43)}) ?
                               (~$unsigned((8'ha6))) : (|wire192[(2'h2):(1'h0)])) : wire193)};
  assign wire198 = wire192;
  assign wire199 = $signed(wire191[(4'ha):(4'ha)]);
  assign wire200 = (wire195[(4'hb):(2'h3)] ?
                       ($unsigned((wire191[(2'h2):(2'h2)] ?
                           ((8'haf) >>> wire195) : (+wire194))) * (~^(wire194[(3'h6):(1'h0)] ?
                           $unsigned(wire197) : (~(8'ha4))))) : {wire192,
                           {$unsigned({wire196})}});
  assign wire201 = (~|(8'hb6));
  assign wire202 = (8'hb0);
  always
    @(posedge clk) begin
      reg203 <= $signed((-{((+wire194) || (8'hb2)),
          ({wire193, wire196} << {wire199, (8'hb7)})}));
      reg204 <= wire196[(5'h14):(3'h5)];
      reg205 <= (|$signed(wire195));
      reg206 <= wire198;
      if (((wire198[(3'h6):(2'h3)] ?
          $unsigned(reg206[(3'h5):(3'h4)]) : wire195) >>> $unsigned(wire196[(3'h5):(3'h5)])))
        begin
          reg207 <= $signed(((|wire192) | $unsigned((-wire198))));
          if ($signed($unsigned($signed(wire192))))
            begin
              reg208 <= (($signed(($unsigned(wire192) ?
                  (reg203 ? wire202 : reg203) : {wire193,
                      reg206})) * wire197[(3'h5):(1'h0)]) << (~|$signed($signed((wire193 + reg207)))));
              reg209 <= $unsigned(reg208);
              reg210 <= wire198[(2'h2):(2'h2)];
            end
          else
            begin
              reg208 <= reg209[(1'h0):(1'h0)];
              reg209 <= (((~^$unsigned(reg205[(4'h8):(3'h5)])) < (((wire202 ?
                          wire200 : wire194) ?
                      (~^wire195) : (wire196 == reg207)) ?
                  wire199 : ($signed(wire195) == (reg203 > wire194)))) << ({reg206,
                  $signed(((8'ha9) ? wire197 : wire194))} ~^ $signed((8'hac))));
              reg210 <= {($unsigned(reg208[(3'h6):(3'h4)]) == wire192[(4'hc):(4'h8)])};
              reg211 <= wire191[(3'h6):(2'h2)];
              reg212 <= ((8'hb6) ~^ (^~(~|wire191[(4'h8):(2'h2)])));
            end
          reg213 <= ((reg207[(1'h1):(1'h1)] >= $unsigned(reg211)) ?
              {(wire196[(1'h1):(1'h0)] ^~ $signed(((8'haf) ?
                      (8'hac) : wire195)))} : reg203[(4'ha):(3'h4)]);
          reg214 <= (-$unsigned($unsigned(reg207[(5'h10):(2'h2)])));
          reg215 <= ($unsigned($signed({(8'hbe)})) ?
              wire199[(3'h6):(2'h3)] : $signed((($signed(reg203) + {wire202,
                      (8'ha4)}) ?
                  reg207[(3'h5):(3'h5)] : $unsigned(wire196[(3'h4):(1'h1)]))));
        end
      else
        begin
          if (wire191[(4'h9):(1'h1)])
            begin
              reg207 <= reg207;
              reg208 <= wire201[(3'h5):(2'h3)];
              reg209 <= {$unsigned($signed(({reg207} ~^ reg211))),
                  $unsigned((reg206[(3'h4):(2'h2)] ?
                      wire194[(2'h3):(2'h3)] : $signed(reg203[(3'h5):(1'h0)])))};
              reg210 <= ((-((!(~&wire193)) ? reg204[(1'h1):(1'h0)] : (8'h9f))) ?
                  ((+(wire194 ?
                      (~^wire202) : (wire196 ?
                          (7'h40) : wire201))) == (($signed(wire192) ?
                      wire192[(4'ha):(4'h9)] : (wire201 ^ wire202)) && ((wire196 ?
                          (8'ha1) : wire201) ?
                      $unsigned(wire198) : (reg209 ?
                          reg212 : reg212)))) : (~|$unsigned(($signed(reg208) ?
                      (~&reg211) : $unsigned((8'hac))))));
              reg211 <= reg214[(5'h12):(1'h1)];
            end
          else
            begin
              reg207 <= ($signed({wire195[(4'hf):(4'he)]}) ^ reg213[(4'hd):(3'h4)]);
              reg208 <= reg210[(3'h7):(1'h1)];
              reg209 <= (-($signed(((~^reg209) < reg209[(2'h3):(1'h1)])) ^~ ($unsigned((|(7'h40))) ?
                  $signed({wire191}) : wire201[(4'hc):(2'h3)])));
            end
          reg212 <= {({$unsigned($unsigned(wire198)),
                  reg210[(3'h4):(1'h1)]} * wire195),
              $unsigned((-reg212))};
          if ((~|{reg207[(3'h4):(1'h1)], reg207[(4'hf):(4'he)]}))
            begin
              reg213 <= $unsigned(reg212[(3'h4):(2'h2)]);
              reg214 <= $signed($unsigned(((~&(wire195 ? (8'haa) : wire196)) ?
                  (wire195[(4'h8):(3'h7)] && $signed(wire195)) : ($unsigned(wire193) != wire200[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg213 <= (reg209 <= wire199[(3'h7):(2'h3)]);
              reg214 <= ($unsigned($signed((&(-wire197)))) >= wire195[(4'h9):(3'h6)]);
            end
          if (reg213[(3'h4):(1'h0)])
            begin
              reg215 <= ($unsigned({$signed((reg213 + reg206)),
                  reg203[(3'h7):(3'h5)]}) > ({$signed(((8'hb1) ?
                          reg215 : reg213)),
                      reg211} ?
                  (wire194[(4'h9):(2'h3)] ^ ({reg205} ?
                      (wire200 ^ reg214) : ((8'haa) | reg213))) : $unsigned((^~(reg209 ?
                      wire194 : wire197)))));
              reg216 <= $unsigned($unsigned($signed(reg205[(4'h8):(1'h1)])));
              reg217 <= (((-(~&reg209)) ?
                      $unsigned({$signed(wire192)}) : reg214) ?
                  wire201[(4'hd):(3'h4)] : (~&($unsigned(((8'ha2) ^ reg215)) ?
                      $unsigned((wire192 == reg213)) : ((wire199 >= reg209) ?
                          wire199 : (wire194 + reg207)))));
              reg218 <= wire202;
            end
          else
            begin
              reg215 <= reg208[(2'h2):(1'h1)];
              reg216 <= (~|reg207[(3'h4):(2'h3)]);
            end
          reg219 <= (((8'h9d) + (~|{(reg213 ?
                  reg215 : reg216)})) ~^ wire198[(2'h2):(2'h2)]);
        end
    end
  assign wire220 = ({(($unsigned(wire199) ?
                           (!reg206) : ((8'hba) ?
                               wire195 : reg210)) ~^ wire195),
                       $unsigned(($signed(wire196) ?
                           reg212[(1'h1):(1'h1)] : (reg214 ^ reg214)))} <<< {$signed($unsigned((8'hae))),
                       (reg216 ? {((8'h9f) ? reg209 : (8'h9e))} : reg213)});
  assign wire221 = reg208[(3'h7):(3'h7)];
  assign wire222 = $signed($unsigned((($signed(wire220) > {wire195}) ?
                       $unsigned(reg207) : reg211)));
  assign wire223 = (~(~^(~&wire195[(4'h9):(3'h6)])));
  assign wire224 = ($unsigned($unsigned($signed((-reg205)))) << (!$signed((8'ha1))));
  always
    @(posedge clk) begin
      reg225 <= ((reg206 != $unsigned((^(wire222 || reg217)))) ?
          $unsigned(wire222[(2'h3):(2'h3)]) : reg209[(4'h8):(3'h7)]);
    end
  assign wire226 = $signed((&wire194));
  assign wire227 = {{$unsigned(($unsigned(reg209) >>> $signed(reg212)))},
                       {$signed({(reg225 ? reg208 : reg208)})}};
  always
    @(posedge clk) begin
      if ((~{{((reg206 >> wire197) ? (~wire194) : (reg209 * reg209))}}))
        begin
          if ($unsigned((reg218 ?
              $signed($unsigned((+reg207))) : (((reg205 | wire224) ?
                  $signed((8'ha6)) : wire220) ^ $unsigned($signed(wire223))))))
            begin
              reg228 <= (!(8'hac));
              reg229 <= reg225[(3'h4):(2'h2)];
              reg230 <= wire202;
              reg231 <= $unsigned(((($unsigned(wire194) <<< (+wire201)) ?
                      $signed($signed(wire226)) : $signed($signed(reg203))) ?
                  $signed((reg204[(2'h2):(1'h1)] < (reg229 ^ (8'hb4)))) : ($signed($unsigned((8'hb2))) ?
                      ((~|reg217) || $signed(reg204)) : (-{(8'h9e),
                          wire223}))));
              reg232 <= ((reg210[(4'h9):(1'h0)] ?
                  $signed($signed($signed((8'hab)))) : $unsigned(((~reg212) ?
                      $unsigned(reg208) : {wire220}))) * (wire223 ?
                  (reg231[(3'h6):(2'h3)] << wire198) : {reg229}));
            end
          else
            begin
              reg228 <= (&reg214);
              reg229 <= ({((~&(wire227 ?
                          wire220 : reg231)) ~^ reg206[(4'h8):(2'h3)]),
                      wire192} ?
                  (~&($unsigned(((8'hae) ?
                      wire199 : wire197)) ~^ {(reg214 >> reg209)})) : ({($signed(wire196) <= reg229),
                      ((~reg228) ?
                          $signed(reg204) : $unsigned(reg203))} | (reg205[(3'h6):(3'h6)] ~^ ((reg230 ?
                          reg231 : wire226) ?
                      {(7'h42)} : (reg217 <<< (8'hb5))))));
            end
          reg233 <= wire220[(4'h8):(3'h5)];
        end
      else
        begin
          if ((|($unsigned((+$signed(reg233))) ?
              wire199 : (~$signed($signed(reg211))))))
            begin
              reg228 <= wire221[(4'hd):(4'hd)];
              reg229 <= ((wire195[(4'ha):(4'ha)] <= $signed((wire227[(3'h7):(3'h7)] >> $unsigned((8'ha7))))) ?
                  $unsigned({$unsigned(reg207),
                      ((-wire223) ?
                          (~wire196) : (wire198 ?
                              wire221 : reg217))}) : $signed({(8'ha5),
                      {$signed(wire227)}}));
              reg230 <= $signed(($unsigned(reg206[(3'h7):(3'h5)]) ?
                  (|(~wire198[(1'h1):(1'h1)])) : (^~$unsigned($signed(reg213)))));
            end
          else
            begin
              reg228 <= $signed($unsigned($signed($signed((reg215 ?
                  reg203 : wire201)))));
              reg229 <= ((((~&$unsigned(wire201)) ?
                      ($signed(wire227) + wire194[(3'h6):(1'h1)]) : wire222[(2'h2):(1'h1)]) >= (wire199[(1'h1):(1'h0)] >> $unsigned(reg217[(4'h9):(4'h8)]))) ?
                  wire226 : wire196[(3'h6):(2'h2)]);
              reg230 <= ($unsigned({reg225}) ?
                  ($unsigned(({reg218} & (wire226 ?
                      reg211 : wire199))) | $signed($signed((wire227 ?
                      wire226 : wire200)))) : wire200[(4'hc):(3'h4)]);
              reg231 <= ($unsigned({(((8'ha5) ^~ (8'hab)) ?
                      (reg218 ?
                          wire198 : reg210) : (wire197 << wire221))}) >> {(~(((8'ha2) ?
                      wire192 : reg207) + wire198))});
              reg232 <= reg225;
            end
          if ($signed($unsigned($unsigned(wire195))))
            begin
              reg233 <= reg232[(4'hf):(3'h5)];
              reg234 <= $signed(((~|$signed(reg207[(4'hc):(3'h6)])) != {($unsigned(reg212) * wire197),
                  reg211[(1'h1):(1'h0)]}));
            end
          else
            begin
              reg233 <= $unsigned($signed(({(wire222 && (8'ha2)),
                  (wire201 ? reg209 : reg203)} || reg210[(1'h1):(1'h1)])));
              reg234 <= (((reg228 << ((~^wire197) && $unsigned(wire220))) ?
                      $signed($signed($unsigned((8'ha0)))) : $signed(((~|reg219) ?
                          (wire220 ? reg234 : reg232) : $unsigned(reg229)))) ?
                  ((^~{reg210[(5'h10):(1'h0)]}) ~^ (7'h41)) : reg218[(2'h2):(2'h2)]);
              reg235 <= (({((wire223 ?
                          reg230 : reg208) * reg211[(2'h2):(1'h0)]),
                      {(wire227 ? wire192 : wire201), $unsigned(reg219)}} ?
                  ($signed($signed(wire226)) ?
                      {reg216, {wire191}} : (wire196 >= (reg229 ?
                          reg207 : (8'hb0)))) : ($signed(((8'hae) ?
                      wire194 : reg203)) ~^ (reg229 ?
                      (wire195 ?
                          wire197 : (8'ha5)) : $unsigned(wire224)))) ~^ ({(reg218 ?
                          (reg203 >> wire201) : reg204[(3'h4):(1'h0)]),
                      $signed((reg233 - wire223))} ?
                  (8'h9c) : (~|{$signed((8'hbe)), (wire199 <= reg234)})));
              reg236 <= reg218;
            end
          reg237 <= $signed(wire196);
        end
    end
  assign wire238 = wire191[(3'h4):(2'h2)];
  module239 modinst318 (.wire241(reg233), .wire243(wire193), .y(wire317), .wire242(wire224), .clk(clk), .wire240(wire202));
  assign wire319 = {$signed(((((8'hb6) ? wire226 : reg229) ?
                               wire238[(4'ha):(3'h4)] : (wire226 ?
                                   wire193 : wire193)) ?
                           $signed(reg216) : (((8'haa) ?
                               reg215 : reg234) * $unsigned(wire222))))};
  assign wire320 = wire226[(4'hf):(1'h0)];
  assign wire321 = ($unsigned(($unsigned((8'hab)) * ($unsigned((7'h41)) == $signed(reg234)))) ?
                       $signed(reg206[(3'h6):(3'h4)]) : (~wire193[(3'h5):(3'h5)]));
  assign wire322 = $unsigned((!reg219));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module29
#( parameter param186 = ((((((8'hac) | (8'ha9)) * (8'hbc)) << (^~((8'ha7) ? (7'h40) : (8'hb4)))) & (8'ha2)) - (^~{(((8'ha3) | (8'h9d)) <<< ((8'h9d) << (8'hbe)))})) )
(y, clk, wire33, wire32, wire31, wire30);
  output wire [(32'h78):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire33;
  input wire [(5'h14):(1'h0)] wire32;
  input wire [(5'h13):(1'h0)] wire31;
  input wire signed [(5'h10):(1'h0)] wire30;
  wire signed [(5'h10):(1'h0)] wire185;
  wire signed [(4'hf):(1'h0)] wire184;
  wire [(4'hb):(1'h0)] wire183;
  wire [(5'h15):(1'h0)] wire182;
  wire signed [(4'ha):(1'h0)] wire125;
  wire signed [(2'h2):(1'h0)] wire75;
  wire signed [(3'h4):(1'h0)] wire74;
  wire signed [(4'hb):(1'h0)] wire72;
  wire [(5'h15):(1'h0)] wire34;
  wire signed [(4'h8):(1'h0)] wire180;
  assign y = {wire185,
                 wire184,
                 wire183,
                 wire182,
                 wire125,
                 wire75,
                 wire74,
                 wire72,
                 wire34,
                 wire180,
                 (1'h0)};
  assign wire34 = $signed(({(wire33 - (wire33 >= (8'ha2)))} ?
                      wire30[(2'h2):(1'h1)] : ((^~(wire32 || wire33)) ?
                          wire33 : $signed(((8'ha2) ^ (8'haa))))));
  module35 modinst73 (wire72, clk, wire32, wire30, wire33, wire31);
  assign wire74 = (8'hb0);
  assign wire75 = wire34;
  module76 modinst126 (wire125, clk, wire31, wire30, wire74, wire32, wire72);
  module127 modinst181 (.y(wire180), .wire132(wire30), .wire128(wire32), .wire130(wire34), .wire131(wire31), .clk(clk), .wire129(wire33));
  assign wire182 = (wire125 >> $signed($unsigned($signed(wire75[(2'h2):(1'h1)]))));
  assign wire183 = {$unsigned(wire72)};
  assign wire184 = $signed({wire72[(2'h3):(2'h3)]});
  assign wire185 = wire183;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module127
#( parameter param178 = (|((((8'hb4) >>> (~(8'hbd))) ? {((8'hbf) ? (8'ha0) : (7'h40))} : (((8'ha3) <= (8'hb2)) ? ((7'h40) ? (8'haf) : (8'hab)) : {(8'hb6), (8'hba)})) ~^ {(((7'h41) <= (8'ha2)) ? (~|(8'ha6)) : (|(8'hb5))), (((8'hae) * (8'hba)) ? ((8'h9d) >> (8'hb5)) : {(8'ha2)})}))
, parameter param179 = {param178, ((~(~{(8'ha7), param178})) >= {((param178 ? param178 : param178) ? param178 : ((8'ha3) ? param178 : (8'ha6))), param178})} )
(y, clk, wire132, wire131, wire130, wire129, wire128);
  output wire [(32'h1fe):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire132;
  input wire signed [(5'h12):(1'h0)] wire131;
  input wire [(5'h15):(1'h0)] wire130;
  input wire signed [(3'h6):(1'h0)] wire129;
  input wire [(5'h12):(1'h0)] wire128;
  wire [(3'h4):(1'h0)] wire177;
  reg [(2'h3):(1'h0)] reg176 = (1'h0);
  reg [(2'h3):(1'h0)] reg175 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg174 = (1'h0);
  reg [(5'h10):(1'h0)] reg173 = (1'h0);
  reg [(5'h15):(1'h0)] reg172 = (1'h0);
  reg [(2'h2):(1'h0)] reg171 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg170 = (1'h0);
  reg [(4'h9):(1'h0)] reg169 = (1'h0);
  reg [(2'h3):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg167 = (1'h0);
  reg [(4'he):(1'h0)] reg166 = (1'h0);
  reg [(5'h15):(1'h0)] reg165 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg164 = (1'h0);
  reg [(3'h5):(1'h0)] reg163 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg162 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg161 = (1'h0);
  reg [(2'h3):(1'h0)] reg160 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg159 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg158 = (1'h0);
  reg [(3'h7):(1'h0)] reg157 = (1'h0);
  reg [(5'h15):(1'h0)] reg156 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg155 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg154 = (1'h0);
  reg [(3'h7):(1'h0)] reg153 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg152 = (1'h0);
  reg [(4'hd):(1'h0)] reg151 = (1'h0);
  reg [(4'h8):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg148 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg146 = (1'h0);
  reg [(4'hc):(1'h0)] reg145 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg143 = (1'h0);
  reg [(5'h15):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg141 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg140 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg139 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg138 = (1'h0);
  reg [(3'h5):(1'h0)] reg137 = (1'h0);
  wire [(5'h14):(1'h0)] wire136;
  wire [(4'hb):(1'h0)] wire135;
  wire [(4'h9):(1'h0)] wire134;
  wire [(4'h9):(1'h0)] wire133;
  assign y = {wire177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 wire136,
                 wire135,
                 wire134,
                 wire133,
                 (1'h0)};
  assign wire133 = ($unsigned((wire132[(3'h7):(1'h0)] == $unsigned(wire130))) && $signed($signed(wire129)));
  assign wire134 = (wire130[(5'h12):(3'h6)] ?
                       (wire132 ? wire130 : wire130) : wire131);
  assign wire135 = (($unsigned($signed((~&wire134))) >>> wire131[(1'h1):(1'h1)]) ?
                       {wire133[(3'h4):(2'h2)],
                           (((wire132 > wire131) ?
                                   (wire129 ?
                                       wire132 : (8'hb1)) : (wire134 & wire134)) ?
                               wire134[(3'h5):(3'h4)] : {wire132,
                                   $signed((8'hbb))})} : wire128[(2'h3):(2'h2)]);
  assign wire136 = $signed(wire133);
  always
    @(posedge clk) begin
      if (wire136[(5'h14):(4'he)])
        begin
          if ((($signed(wire135[(1'h1):(1'h0)]) - $signed($unsigned((~&wire134)))) ?
              $signed($signed(wire136[(3'h7):(3'h5)])) : {$unsigned(($unsigned((8'had)) >= (wire129 ?
                      wire136 : (8'h9c))))}))
            begin
              reg137 <= ((^((+(7'h42)) ~^ ({wire135} ?
                      (^~wire133) : (wire130 < wire133)))) ?
                  $signed(wire135[(3'h4):(2'h3)]) : $unsigned(wire130));
              reg138 <= {$signed({(8'ha1)})};
            end
          else
            begin
              reg137 <= $unsigned(wire135[(3'h4):(2'h3)]);
              reg138 <= {$signed(wire136), wire128};
            end
          reg139 <= wire135;
        end
      else
        begin
          if ((~^((^~$unsigned({wire133})) + $unsigned(wire130))))
            begin
              reg137 <= (~$unsigned($unsigned(($unsigned(wire135) ?
                  $signed(wire136) : (!wire134)))));
              reg138 <= (wire134 != wire129);
            end
          else
            begin
              reg137 <= (~|$unsigned(wire135[(3'h7):(3'h6)]));
              reg138 <= (wire132[(4'he):(1'h1)] != ((wire134[(2'h2):(1'h0)] & $signed(wire132[(3'h5):(2'h2)])) <<< wire133[(4'h9):(4'h8)]));
              reg139 <= ((8'hbb) | ((reg138[(3'h4):(1'h1)] > wire128[(4'hd):(4'hd)]) ?
                  $unsigned(((~^wire130) >>> wire128[(5'h10):(4'ha)])) : (wire128 ?
                      wire136[(4'hc):(3'h6)] : $signed($unsigned(wire132)))));
              reg140 <= $signed($unsigned(wire133));
              reg141 <= (~&(8'had));
            end
        end
      if (reg140)
        begin
          reg142 <= wire135;
          reg143 <= (~&reg142[(3'h7):(3'h4)]);
        end
      else
        begin
          reg142 <= reg140[(3'h4):(1'h0)];
          reg143 <= {$signed(reg142)};
          reg144 <= (reg142 << {wire130,
              $signed(((wire133 && (8'hab)) >= (wire130 ? reg141 : wire136)))});
          if (((^($signed((wire129 ? (8'hbd) : reg142)) ?
              $signed((wire132 >= wire136)) : {$unsigned(wire134),
                  reg140[(4'he):(4'h9)]})) * ((wire133 ?
                  ({wire134} ?
                      wire133 : (~|reg144)) : (|(wire136 ~^ wire129))) ?
              (~&wire135) : (!((reg138 ?
                  (8'hba) : reg139) >> (reg138 >> reg142))))))
            begin
              reg145 <= ($signed({($unsigned(wire128) ?
                      reg141[(1'h1):(1'h1)] : reg144),
                  (-$unsigned(reg140))}) > ($signed(((&wire134) <= (wire132 >> wire136))) <<< $unsigned(((reg143 ~^ wire133) <<< (-wire129)))));
              reg146 <= (($unsigned($signed({wire135})) ?
                  $signed((reg143 ?
                      wire132 : {(8'hb7),
                          (8'ha9)})) : (+(^$unsigned(wire131)))) << reg137);
            end
          else
            begin
              reg145 <= $unsigned(wire128[(4'hf):(4'ha)]);
              reg146 <= wire128[(2'h2):(1'h1)];
              reg147 <= wire136[(4'he):(3'h4)];
              reg148 <= $signed($signed(($unsigned({wire128}) && $unsigned((wire130 ?
                  reg140 : reg147)))));
              reg149 <= reg147[(3'h5):(2'h2)];
            end
          reg150 <= wire132;
        end
      reg151 <= reg146;
    end
  always
    @(posedge clk) begin
      reg152 <= ((+$unsigned((reg141[(2'h2):(1'h0)] > (wire132 <<< wire131)))) == reg141[(3'h5):(1'h1)]);
      reg153 <= ($unsigned(wire136[(2'h2):(1'h1)]) == (~|reg141));
      if ($unsigned($unsigned(($signed((wire133 ? reg150 : reg139)) ?
          $signed(reg153) : reg147))))
        begin
          reg154 <= (((^~(~$signed(wire133))) ?
                  {wire129} : reg140[(2'h3):(2'h3)]) ?
              (reg138 * $signed((^~$signed(reg144)))) : reg146);
        end
      else
        begin
          reg154 <= $signed(reg148);
          reg155 <= (~$unsigned($unsigned(reg153[(3'h5):(2'h3)])));
          if ($unsigned(wire128[(3'h6):(2'h2)]))
            begin
              reg156 <= (~((&(((7'h40) ?
                      reg154 : wire131) <= $signed((8'haf)))) ?
                  (7'h44) : wire136[(5'h11):(1'h0)]));
              reg157 <= reg140[(3'h7):(3'h5)];
              reg158 <= (reg157 ?
                  {((reg155[(2'h2):(1'h1)] ?
                              (reg151 ?
                                  (8'had) : (8'ha7)) : (wire133 << wire135)) ?
                          wire135[(2'h3):(2'h3)] : reg137[(1'h0):(1'h0)]),
                      reg137[(2'h2):(1'h1)]} : (($unsigned((reg148 ?
                          reg156 : wire128)) << (!(reg139 & wire130))) ?
                      $signed((+{reg144, wire136})) : (7'h41)));
              reg159 <= wire130;
            end
          else
            begin
              reg156 <= wire132[(2'h2):(1'h1)];
              reg157 <= reg143;
              reg158 <= ((~&($signed((reg156 + reg148)) == reg146)) >>> $unsigned({((reg159 - wire128) ?
                      $unsigned(wire133) : $signed(reg159)),
                  (~^$signed((8'hab)))}));
              reg159 <= $signed(reg139[(2'h3):(1'h1)]);
              reg160 <= ((wire133[(1'h0):(1'h0)] ?
                      reg145[(3'h5):(1'h1)] : {{$signed(reg150), {reg145}},
                          reg145}) ?
                  ((~{$signed((8'hb2))}) ?
                      ($unsigned((&reg142)) ?
                          {(reg154 ? reg150 : reg137),
                              $signed(reg137)} : $unsigned((|reg156))) : (($unsigned(reg144) ?
                              $signed(wire134) : reg153[(3'h5):(1'h0)]) ?
                          (reg154 ~^ reg155[(4'ha):(4'ha)]) : ((reg153 + (8'haa)) ?
                              $unsigned(wire130) : $unsigned(wire130)))) : {$unsigned($signed((|wire135)))});
            end
        end
    end
  always
    @(posedge clk) begin
      reg161 <= $signed($signed({({reg151, reg138} ?
              $signed(wire128) : {reg145})}));
      reg162 <= reg147;
      if ({reg151[(4'h9):(3'h6)], $unsigned(reg152)})
        begin
          if ((($signed($unsigned((wire136 ?
                  reg148 : reg161))) & ((+{wire128}) > ({reg142,
                  reg141} * $signed(reg155)))) ?
              (^~($signed($unsigned(reg155)) <= ($signed((8'ha3)) ?
                  (wire128 ?
                      wire136 : reg160) : (reg157 & reg140)))) : ((+reg139) + reg138)))
            begin
              reg163 <= ($unsigned($signed((!(reg155 >> reg151)))) & reg160);
            end
          else
            begin
              reg163 <= ((($signed($unsigned((8'hb5))) ?
                          reg143[(5'h10):(2'h3)] : ((reg155 == reg156) ?
                              (reg140 << (8'hb5)) : $unsigned(reg142))) ?
                      $unsigned((reg156[(5'h10):(2'h2)] ?
                          (wire131 ^~ (8'h9d)) : (8'h9e))) : wire136) ?
                  (reg144 ?
                      $signed((~|wire129)) : ($unsigned((~reg153)) ?
                          wire133[(3'h6):(2'h2)] : (reg151 | (reg152 == reg147)))) : $signed(((reg156[(5'h14):(2'h2)] + (wire131 | reg156)) ?
                      (|((8'hab) ? wire130 : wire135)) : (^~$signed(reg142)))));
            end
          reg164 <= $signed($unsigned((-reg156)));
          reg165 <= (8'hb2);
          if ((^~reg142))
            begin
              reg166 <= ({({$unsigned(reg141), {reg162}} ?
                          (8'h9c) : ($unsigned(wire130) ?
                              (reg158 ?
                                  (8'hb3) : wire130) : $unsigned(wire131)))} ?
                  (|((|(wire132 ^~ reg154)) ^ (reg139 ?
                      (reg154 <= (8'ha9)) : (&reg149)))) : {(($unsigned(reg147) ?
                              (^reg141) : ((8'hb0) ? wire131 : wire131)) ?
                          ((reg143 ? reg153 : (8'hbd)) ?
                              wire135 : ((8'h9c) << wire135)) : ((reg162 >> wire132) ?
                              (reg153 << reg147) : {reg153, reg139}))});
              reg167 <= (-$signed(wire131[(3'h5):(3'h4)]));
              reg168 <= $unsigned(reg145);
              reg169 <= $unsigned($unsigned(((reg139 < (reg152 ?
                  reg149 : reg164)) << ((reg157 ? reg162 : reg141) ?
                  (wire129 <<< reg144) : ((8'haa) ? reg152 : reg149)))));
            end
          else
            begin
              reg166 <= $unsigned($signed((^~(|wire130))));
              reg167 <= wire133;
              reg168 <= $signed(reg145[(3'h6):(2'h2)]);
              reg169 <= reg159[(3'h4):(2'h3)];
              reg170 <= (($signed(reg137[(3'h4):(3'h4)]) ?
                      $signed(reg167) : {((reg139 >>> reg159) ?
                              (^~reg147) : (!reg154)),
                          ($unsigned((8'hae)) && $unsigned(wire130))}) ?
                  $signed(reg146) : $unsigned($signed((reg159 ?
                      reg163[(1'h0):(1'h0)] : reg137[(2'h2):(1'h1)]))));
            end
        end
      else
        begin
          reg163 <= reg153;
          reg164 <= (|((^~($signed(reg169) ?
                  $unsigned(wire136) : $unsigned(reg157))) ?
              (~&$unsigned($signed((8'hb2)))) : reg137));
        end
      reg171 <= reg170;
    end
  always
    @(posedge clk) begin
      if (reg141[(3'h5):(1'h0)])
        begin
          if (reg160)
            begin
              reg172 <= (wire129[(1'h1):(1'h1)] ?
                  reg149[(3'h6):(1'h1)] : (^~reg138[(2'h2):(1'h1)]));
              reg173 <= (^~wire131);
              reg174 <= ($unsigned(($unsigned((|reg164)) ~^ $unsigned((^wire132)))) || {($signed((reg160 ~^ reg150)) ?
                      $unsigned($unsigned(reg156)) : (~(^wire136)))});
              reg175 <= {(wire131 ?
                      (reg140 ?
                          (reg171 && $signed((7'h41))) : {(reg148 ^~ reg153)}) : $unsigned((((8'hbb) * reg160) ?
                          reg171 : {(8'hb8)}))),
                  $signed(((reg142[(1'h1):(1'h0)] ? (-(8'ha2)) : (~|reg167)) ?
                      ($signed(reg141) ?
                          $unsigned(reg163) : $signed(reg139)) : $signed((reg155 ?
                          reg160 : reg146))))};
            end
          else
            begin
              reg172 <= reg167[(3'h6):(3'h4)];
              reg173 <= $unsigned($signed({reg150, reg138}));
              reg174 <= reg170[(4'hd):(2'h2)];
              reg175 <= {(^($unsigned($signed((8'haa))) ?
                      (^(reg159 ? reg162 : reg151)) : $unsigned({reg143})))};
            end
        end
      else
        begin
          reg172 <= (reg161[(5'h14):(3'h4)] & {(($unsigned(reg175) && $signed(reg150)) < $unsigned(wire131[(3'h4):(1'h1)]))});
        end
      reg176 <= ($unsigned(({reg137[(3'h5):(3'h4)], reg146} ?
              reg158[(4'hd):(4'hb)] : (((8'ha4) && (8'ha9)) ?
                  (reg173 ? reg153 : (8'hb5)) : (reg145 & wire130)))) ?
          (wire130 >>> ($signed((reg140 ? reg139 : (8'h9e))) ?
              reg174 : $unsigned(reg146[(1'h1):(1'h0)]))) : ($signed(reg173[(4'h8):(3'h4)]) && $signed($unsigned((reg150 ?
              wire128 : reg168)))));
    end
  assign wire177 = (|$unsigned($unsigned(($unsigned(reg172) <= reg173))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module76  (y, clk, wire81, wire80, wire79, wire78, wire77);
  output wire [(32'h20f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire81;
  input wire [(4'hf):(1'h0)] wire80;
  input wire signed [(2'h3):(1'h0)] wire79;
  input wire [(5'h12):(1'h0)] wire78;
  input wire [(4'hb):(1'h0)] wire77;
  wire signed [(4'he):(1'h0)] wire124;
  wire [(5'h15):(1'h0)] wire123;
  wire signed [(4'hd):(1'h0)] wire122;
  wire signed [(3'h4):(1'h0)] wire121;
  wire signed [(5'h12):(1'h0)] wire120;
  wire [(4'h9):(1'h0)] wire119;
  wire [(4'hd):(1'h0)] wire118;
  reg signed [(3'h7):(1'h0)] reg117 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg116 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg115 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg114 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg113 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg112 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg110 = (1'h0);
  reg [(4'hd):(1'h0)] reg109 = (1'h0);
  reg [(2'h2):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg106 = (1'h0);
  reg [(5'h13):(1'h0)] reg105 = (1'h0);
  reg [(5'h12):(1'h0)] reg104 = (1'h0);
  reg [(5'h12):(1'h0)] reg103 = (1'h0);
  reg [(2'h3):(1'h0)] reg102 = (1'h0);
  reg [(4'h9):(1'h0)] reg101 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg100 = (1'h0);
  reg [(3'h5):(1'h0)] reg99 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg98 = (1'h0);
  reg [(5'h12):(1'h0)] reg97 = (1'h0);
  reg [(4'hc):(1'h0)] reg96 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire95;
  wire signed [(4'hc):(1'h0)] wire94;
  reg signed [(4'he):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg92 = (1'h0);
  reg [(4'hc):(1'h0)] reg91 = (1'h0);
  reg [(5'h15):(1'h0)] reg90 = (1'h0);
  reg [(4'he):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg88 = (1'h0);
  reg [(5'h14):(1'h0)] reg87 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg86 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg84 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg83 = (1'h0);
  reg [(5'h12):(1'h0)] reg82 = (1'h0);
  assign y = {wire124,
                 wire123,
                 wire122,
                 wire121,
                 wire120,
                 wire119,
                 wire118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 wire95,
                 wire94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire77[(4'h9):(3'h7)])
        begin
          reg82 <= wire81;
          reg83 <= (wire77[(1'h0):(1'h0)] >= $unsigned($unsigned(({wire80,
                  wire81} ?
              reg82 : wire79))));
          reg84 <= (|$signed(wire78[(4'he):(1'h0)]));
          reg85 <= (~(^~$unsigned((wire77 ?
              (wire81 ^ wire81) : (wire80 ~^ wire78)))));
          reg86 <= ($signed($signed(wire80[(1'h0):(1'h0)])) & (+(~(&(wire81 ?
              (8'hbf) : wire80)))));
        end
      else
        begin
          reg82 <= ($unsigned(reg84[(5'h10):(4'h8)]) >= wire77);
          reg83 <= ($unsigned(wire77) ? wire80 : (8'hb7));
          if ((~$signed(reg82[(4'he):(4'h8)])))
            begin
              reg84 <= ({$unsigned($unsigned((reg85 ? (8'hb3) : reg82))),
                  reg84} & (+(($unsigned(wire80) * $unsigned(reg83)) ?
                  (!(&(8'h9e))) : ({reg82} ?
                      $signed(wire78) : (wire79 | (8'hab))))));
            end
          else
            begin
              reg84 <= wire79;
              reg85 <= $signed({$unsigned(reg82), wire79});
              reg86 <= (|(~|$signed((~^reg86[(4'h9):(3'h5)]))));
              reg87 <= {wire78[(4'hd):(4'h9)],
                  ($unsigned($signed({wire81})) ?
                      reg84[(4'ha):(1'h1)] : wire79[(2'h3):(2'h3)])};
              reg88 <= $unsigned((~|(((~|wire78) ?
                      $unsigned(reg84) : reg86[(3'h6):(3'h4)]) ?
                  (|$signed(reg85)) : $unsigned((~&reg84)))));
            end
          if ((~^$unsigned($unsigned(wire80[(3'h7):(1'h0)]))))
            begin
              reg89 <= {$unsigned((wire80[(4'h8):(3'h4)] ?
                      {(-reg84), wire78} : $signed((|reg82))))};
              reg90 <= (~&(|($unsigned((wire80 >>> wire81)) ?
                  (reg84[(5'h11):(2'h2)] - $unsigned(wire78)) : $unsigned($unsigned(reg86)))));
              reg91 <= wire77;
              reg92 <= (($signed({{wire80},
                  ((8'hae) > wire81)}) <= reg82) < (($signed($signed(reg89)) ?
                  (~&reg83) : ($unsigned(reg91) == (~|wire78))) >> ((~^wire80[(3'h7):(2'h2)]) ?
                  $unsigned(wire79[(1'h1):(1'h0)]) : $signed((&reg86)))));
              reg93 <= ($signed(((+$unsigned(reg86)) * reg84)) ?
                  ($unsigned((~^(wire78 >> reg87))) != ((-reg91[(3'h4):(2'h2)]) ?
                      ({reg86, reg83} ?
                          $signed(reg88) : (|(7'h41))) : ((wire77 ?
                          reg86 : wire77) && $unsigned(reg92)))) : $unsigned({$signed(reg88)}));
            end
          else
            begin
              reg89 <= (({(!wire78), reg89} + ($signed((~^reg91)) ?
                  ((reg93 || wire77) || (reg91 ?
                      (8'h9f) : (8'ha6))) : $signed($signed(reg88)))) ^ $signed(($unsigned((~^reg89)) != (+$signed(reg88)))));
              reg90 <= $unsigned(((~^{(!reg90),
                  $unsigned(reg92)}) != (~reg92)));
              reg91 <= $signed($unsigned((|{wire79, (&reg83)})));
              reg92 <= {((|((reg93 >= reg83) ? (|(8'hba)) : (!wire77))) ?
                      (~^reg83) : {({(8'hb5)} ^ reg88), wire81}),
                  $unsigned($signed($unsigned(reg86)))};
              reg93 <= (8'ha3);
            end
        end
    end
  assign wire94 = (|(reg86 <= ((8'ha2) ?
                      ($unsigned(reg86) + reg93[(3'h5):(1'h0)]) : $unsigned(reg88))));
  assign wire95 = reg91[(4'h9):(2'h3)];
  always
    @(posedge clk) begin
      if (reg91[(2'h3):(2'h3)])
        begin
          reg96 <= ((({(wire80 ? wire81 : reg83),
                  {reg93, reg93}} <<< $signed({reg83})) <<< wire79) ?
              $unsigned($signed(({(8'ha4),
                  reg89} == $unsigned(reg91)))) : ({reg92[(2'h2):(1'h0)],
                      $signed(reg86)} ?
                  (wire77[(4'ha):(3'h6)] < ({wire95} ?
                      {reg83} : (~&(8'hbd)))) : ($unsigned(wire77[(4'h9):(1'h1)]) < $unsigned(wire95))));
          reg97 <= $signed((reg93 ^ $unsigned(wire77)));
        end
      else
        begin
          if ((~(($signed((reg88 <= wire79)) ?
              $signed($signed(reg86)) : ((wire95 ?
                  wire95 : reg85) & $signed((8'hac)))) <<< (~(+$unsigned(reg84))))))
            begin
              reg96 <= (((((reg82 <<< reg82) >> (7'h43)) ?
                      wire79 : reg90[(5'h12):(5'h10)]) ?
                  (~&(&(!wire77))) : ($signed({reg97}) << reg89)) + (((!((8'haf) ?
                          reg83 : reg87)) ?
                      ($unsigned(reg85) << $signed(reg92)) : reg91[(1'h0):(1'h0)]) ?
                  {$signed($unsigned(wire79)),
                      ((8'h9d) ?
                          reg91 : $unsigned(wire95))} : {$signed((reg87 > reg88)),
                      wire78}));
              reg97 <= (!$unsigned(({$unsigned(reg91)} ?
                  reg90 : (&(reg92 ? reg89 : reg97)))));
              reg98 <= $signed({(wire95[(3'h7):(3'h4)] ?
                      $signed(wire95[(4'h9):(3'h5)]) : reg97[(3'h4):(3'h4)])});
              reg99 <= (reg93 ^~ (8'hb6));
            end
          else
            begin
              reg96 <= (8'ha2);
              reg97 <= {(((+$unsigned(reg91)) ?
                          $signed($signed(reg96)) : (!(wire80 >>> wire94))) ?
                      ({(reg92 ? (8'ha4) : wire77),
                          reg92[(2'h2):(2'h2)]} & $signed($unsigned(reg91))) : (~&reg91[(3'h5):(2'h2)]))};
              reg98 <= (({$signed((reg90 ? wire77 : (8'h9c))),
                  $unsigned((reg87 ?
                      (8'ha1) : (8'hb2)))} ^ (~^reg86[(1'h1):(1'h1)])) - ((^{$signed(reg96),
                  $unsigned(reg82)}) <<< $unsigned($unsigned(((8'had) >= (8'hb5))))));
              reg99 <= (~(~|reg88[(3'h5):(2'h2)]));
              reg100 <= wire81;
            end
          if ($unsigned(((($signed(reg86) <<< reg85) < wire95) == (($unsigned(reg89) <<< (wire94 ?
              wire80 : reg88)) << (-$unsigned(wire95))))))
            begin
              reg101 <= reg85;
              reg102 <= ((8'hb5) - (|{(reg100 ?
                      (reg83 ? wire81 : wire95) : {(8'hb7), wire81})}));
              reg103 <= $signed($unsigned((^wire80[(1'h1):(1'h0)])));
              reg104 <= $unsigned((8'hb1));
              reg105 <= $unsigned(reg85);
            end
          else
            begin
              reg101 <= $unsigned((^$signed($signed(reg84))));
              reg102 <= ($unsigned({$unsigned({(8'hbc),
                      reg88})}) << (^{wire81}));
              reg103 <= ($signed((-$unsigned((+(8'hbf))))) ?
                  wire94 : ((reg86[(1'h0):(1'h0)] ?
                          $signed({reg105, reg96}) : (~$unsigned(wire81))) ?
                      {$signed((~^(8'hac))),
                          (reg98[(4'h9):(1'h0)] ?
                              reg97 : $signed(reg98))} : (-(|reg88[(4'hf):(4'h9)]))));
              reg104 <= wire95[(4'h8):(2'h3)];
            end
          if ({($unsigned(($unsigned(wire77) ?
                  ((8'hbd) >> reg104) : $unsigned(reg97))) <<< ($signed((+reg83)) & ((wire78 >> (8'ha0)) | $signed(reg92)))),
              ((~|((reg99 ? (7'h42) : reg104) & (wire94 ?
                  wire80 : reg89))) > (^~$signed(reg92[(1'h1):(1'h1)])))})
            begin
              reg106 <= (8'h9f);
              reg107 <= $unsigned(((~|(8'ha2)) ?
                  {reg90[(5'h12):(3'h4)],
                      $signed($unsigned(reg106))} : ($signed((^~reg86)) ^ {(reg101 * reg102)})));
              reg108 <= $unsigned(reg105[(4'he):(3'h4)]);
              reg109 <= $unsigned({$unsigned({(8'hbb), (wire77 ~^ wire79)})});
            end
          else
            begin
              reg106 <= reg83;
              reg107 <= reg103[(5'h10):(3'h7)];
              reg108 <= (!reg93[(2'h2):(1'h1)]);
              reg109 <= ((reg107 != $unsigned((~|reg90[(4'hc):(4'h9)]))) ?
                  (+reg86) : {$unsigned((wire81[(3'h4):(2'h3)] ?
                          {(8'hbd), reg92} : $unsigned(reg99))),
                      (reg85 <= ((-reg96) >> (wire79 ? wire80 : reg91)))});
              reg110 <= reg102[(2'h3):(1'h0)];
            end
          if (reg82)
            begin
              reg111 <= $unsigned($signed($unsigned(($signed(reg83) ?
                  {reg82} : {(8'ha2), (8'ha1)}))));
              reg112 <= $signed($signed(reg101[(4'h8):(3'h7)]));
              reg113 <= reg99[(2'h2):(2'h2)];
              reg114 <= (reg100 ?
                  reg102[(2'h3):(1'h1)] : $signed((~&$signed($unsigned(reg88)))));
              reg115 <= reg107;
            end
          else
            begin
              reg111 <= $signed((~|{($unsigned(reg98) | (!(8'hb0)))}));
              reg112 <= reg101;
            end
          reg116 <= (!$unsigned((($signed(reg106) < {wire80, reg83}) ?
              $unsigned((~|reg106)) : reg108)));
        end
      reg117 <= ({{$signed((!wire94)),
              $unsigned(reg109)}} <= $unsigned($signed($signed((~reg84)))));
    end
  assign wire118 = reg99;
  assign wire119 = reg96;
  assign wire120 = reg105[(5'h12):(1'h1)];
  assign wire121 = ($signed($unsigned(($signed((8'hbc)) ?
                       $unsigned(wire78) : $unsigned(reg98)))) << (&reg102));
  assign wire122 = reg105[(4'hb):(4'hb)];
  assign wire123 = wire94[(3'h7):(3'h6)];
  assign wire124 = (|reg111[(3'h6):(1'h0)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module35  (y, clk, wire39, wire38, wire37, wire36);
  output wire [(32'h166):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire39;
  input wire [(4'h8):(1'h0)] wire38;
  input wire [(4'hc):(1'h0)] wire37;
  input wire [(2'h2):(1'h0)] wire36;
  wire signed [(4'hc):(1'h0)] wire71;
  reg signed [(3'h6):(1'h0)] reg70 = (1'h0);
  reg [(4'he):(1'h0)] reg69 = (1'h0);
  reg [(4'h8):(1'h0)] reg68 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire67;
  wire [(4'hd):(1'h0)] wire66;
  reg signed [(3'h4):(1'h0)] reg65 = (1'h0);
  reg signed [(4'he):(1'h0)] reg64 = (1'h0);
  reg signed [(4'he):(1'h0)] reg63 = (1'h0);
  reg [(4'ha):(1'h0)] reg62 = (1'h0);
  reg [(3'h7):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg60 = (1'h0);
  reg [(2'h2):(1'h0)] reg59 = (1'h0);
  reg [(5'h12):(1'h0)] reg58 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg57 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg56 = (1'h0);
  reg [(3'h6):(1'h0)] reg55 = (1'h0);
  reg [(3'h7):(1'h0)] reg54 = (1'h0);
  reg [(5'h11):(1'h0)] reg53 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg52 = (1'h0);
  reg [(5'h11):(1'h0)] reg51 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg50 = (1'h0);
  reg [(4'h8):(1'h0)] reg49 = (1'h0);
  reg [(4'he):(1'h0)] reg48 = (1'h0);
  reg [(4'hb):(1'h0)] reg47 = (1'h0);
  reg [(5'h10):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg45 = (1'h0);
  reg [(4'hc):(1'h0)] reg44 = (1'h0);
  reg [(2'h3):(1'h0)] reg43 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg41 = (1'h0);
  reg [(4'hc):(1'h0)] reg40 = (1'h0);
  assign y = {wire71,
                 reg70,
                 reg69,
                 reg68,
                 wire67,
                 wire66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($signed(wire39))
        begin
          reg40 <= (|$signed({wire38[(3'h6):(1'h0)],
              ((wire36 ? wire37 : (8'h9e)) ?
                  wire39[(4'hf):(2'h2)] : wire38[(1'h0):(1'h0)])}));
          reg41 <= $unsigned(reg40[(2'h2):(1'h0)]);
        end
      else
        begin
          reg40 <= wire37[(3'h4):(2'h3)];
          reg41 <= wire37[(4'hb):(1'h1)];
          if ({$signed($signed((wire36[(1'h0):(1'h0)] ?
                  $unsigned(reg41) : $unsigned(reg41))))})
            begin
              reg42 <= ((wire39[(3'h7):(3'h6)] ? $signed(reg41) : {{reg40}}) ?
                  (({wire39, $signed(reg40)} ?
                          (!wire36[(1'h1):(1'h0)]) : wire39) ?
                      reg41 : ($signed(wire36[(1'h0):(1'h0)]) ?
                          ({wire38, (8'hbf)} ?
                              (~^wire39) : (wire37 ^ wire39)) : ($unsigned(reg40) ?
                              {(8'hab), reg40} : (wire39 ?
                                  (8'hb3) : wire36)))) : reg40);
              reg43 <= (!(+($signed($signed(wire36)) < wire36[(2'h2):(1'h1)])));
              reg44 <= (^wire38[(4'h8):(4'h8)]);
              reg45 <= $signed({(^~{$unsigned(reg43)})});
              reg46 <= (^~((reg41 ?
                      reg45 : ($unsigned(reg42) ?
                          $signed(wire39) : $unsigned(wire37))) ?
                  $unsigned(wire38) : (($unsigned(reg42) ?
                          (~&wire39) : wire39) ?
                      ((reg43 <= wire39) ?
                          reg44 : (^(8'ha9))) : $unsigned(reg41))));
            end
          else
            begin
              reg42 <= reg41[(4'hb):(4'ha)];
              reg43 <= wire39[(1'h0):(1'h0)];
              reg44 <= ({{wire39}, reg40[(3'h7):(3'h7)]} + reg42);
            end
        end
      reg47 <= ((-{($signed(reg45) <= reg40)}) >= $unsigned(reg42));
      reg48 <= reg41;
    end
  always
    @(posedge clk) begin
      reg49 <= $signed({reg46[(1'h0):(1'h0)]});
      if (reg43[(2'h2):(1'h0)])
        begin
          if (wire36[(1'h0):(1'h0)])
            begin
              reg50 <= $unsigned(((&$unsigned($signed(reg40))) > (reg48[(1'h0):(1'h0)] ?
                  (~&(~reg48)) : reg44[(4'hc):(4'hb)])));
            end
          else
            begin
              reg50 <= ((&$signed({(wire37 <= wire38), (^reg49)})) ?
                  reg50 : wire37[(3'h4):(1'h1)]);
              reg51 <= ($unsigned((^reg42)) ?
                  $signed((!{$unsigned(reg48)})) : $unsigned((reg50 == ($unsigned(reg50) >> (~|reg49)))));
            end
          reg52 <= reg45[(5'h14):(4'h8)];
        end
      else
        begin
          if ($signed((+reg50[(2'h2):(1'h0)])))
            begin
              reg50 <= (($signed({wire36}) + $unsigned({(+reg41),
                  reg49[(3'h7):(3'h5)]})) + wire37[(3'h6):(1'h0)]);
            end
          else
            begin
              reg50 <= ((+(^(^~reg42[(4'h8):(2'h2)]))) ? (~reg48) : reg40);
              reg51 <= $signed($unsigned(wire36));
            end
        end
      if (((~(reg49[(2'h3):(1'h1)] ?
              reg50[(1'h0):(1'h0)] : ({wire36} ^~ (reg51 ? reg47 : reg52)))) ?
          {(($signed((8'ha4)) != (reg48 == reg45)) ?
                  {reg48} : $unsigned(wire37)),
              (~|{reg42[(1'h1):(1'h0)]})} : ((^~(-(reg40 != reg49))) <= (!(!$unsigned(reg43))))))
        begin
          reg53 <= ((reg47[(1'h1):(1'h0)] ?
              $unsigned(((reg45 ?
                  reg44 : (8'ha8)) + wire39)) : {reg48[(4'he):(2'h3)]}) ^ (!$unsigned($unsigned(reg46))));
        end
      else
        begin
          reg53 <= $signed((reg52[(2'h2):(1'h0)] ?
              $unsigned(((reg46 && reg40) ? {reg40} : (&wire36))) : ((wire39 ?
                      $signed(reg52) : (wire37 * wire36)) ?
                  (+(wire38 ? reg41 : reg48)) : (~reg51[(4'he):(4'ha)]))));
          reg54 <= reg52[(4'hc):(4'h8)];
          reg55 <= $unsigned({wire37[(2'h3):(2'h3)],
              $signed(wire37[(4'h8):(3'h7)])});
          reg56 <= ((reg41 ~^ reg41) ^ reg52);
          reg57 <= ((((8'hac) + ((^~(8'hbe)) ^~ (reg44 >>> wire38))) >>> $unsigned(reg54[(3'h5):(2'h3)])) > $signed((wire36[(2'h2):(1'h0)] ?
              $signed((~reg43)) : reg56[(2'h2):(1'h1)])));
        end
      reg58 <= $unsigned(((8'h9e) ? {$signed((7'h40))} : reg51[(4'ha):(1'h1)]));
      if (((~^wire37[(3'h6):(3'h6)]) < {$signed($signed((reg56 ?
              reg57 : reg56)))}))
        begin
          reg59 <= ({$signed(reg45)} ?
              ((reg48[(3'h5):(3'h4)] && $signed($signed(reg44))) < (+wire36)) : reg53[(4'h9):(1'h0)]);
          reg60 <= ({{((~^(8'ha9)) ? reg44[(3'h5):(1'h1)] : {(8'hba)}),
                  wire36[(1'h0):(1'h0)]},
              reg41[(1'h0):(1'h0)]} >= (($unsigned($signed((8'ha3))) != {reg46}) ?
              reg45 : $unsigned(($signed(reg52) < (wire37 <= reg40)))));
        end
      else
        begin
          reg59 <= $unsigned(reg50[(1'h1):(1'h0)]);
          if (reg54[(1'h0):(1'h0)])
            begin
              reg60 <= reg54[(1'h1):(1'h1)];
              reg61 <= {$signed($unsigned(((|reg51) > ((8'ha3) ?
                      reg48 : reg48))))};
              reg62 <= $unsigned($signed(reg54[(1'h1):(1'h1)]));
              reg63 <= ((8'hb5) > ($unsigned($unsigned(reg61)) ?
                  $unsigned((reg62 >= {reg50,
                      reg45})) : {reg46[(5'h10):(1'h1)]}));
              reg64 <= reg59[(1'h0):(1'h0)];
            end
          else
            begin
              reg60 <= reg57[(1'h1):(1'h1)];
              reg61 <= reg50;
              reg62 <= reg52[(3'h5):(3'h5)];
              reg63 <= $signed(reg43);
              reg64 <= $unsigned({reg55, $signed((&reg54))});
            end
          reg65 <= reg51;
        end
    end
  assign wire66 = $signed(wire38[(1'h1):(1'h0)]);
  assign wire67 = (^$unsigned(reg55));
  always
    @(posedge clk) begin
      reg68 <= $signed(wire37[(2'h3):(1'h1)]);
      reg69 <= (wire36[(2'h2):(2'h2)] <<< reg48);
      reg70 <= (^(((~(|reg48)) + reg42) ?
          $signed($unsigned((~reg49))) : $unsigned({(reg61 ? reg52 : (8'ha2)),
              {(8'ha9), reg58}})));
    end
  assign wire71 = $signed(((reg50[(2'h2):(2'h2)] ?
                          reg64[(4'hc):(4'ha)] : ($unsigned(reg40) * (~reg69))) ?
                      ((8'hac) & (reg48 ?
                          reg49 : {reg46})) : $unsigned(reg70[(3'h5):(3'h5)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module239
#(parameter param316 = {(~&(&{(^~(7'h42))}))})
(y, clk, wire243, wire242, wire241, wire240);
  output wire [(32'h385):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire243;
  input wire [(4'hb):(1'h0)] wire242;
  input wire [(4'hb):(1'h0)] wire241;
  input wire signed [(5'h10):(1'h0)] wire240;
  wire signed [(5'h15):(1'h0)] wire315;
  reg signed [(5'h15):(1'h0)] reg314 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg313 = (1'h0);
  reg [(3'h4):(1'h0)] reg312 = (1'h0);
  wire [(4'hd):(1'h0)] wire311;
  wire signed [(5'h12):(1'h0)] wire310;
  wire signed [(4'h9):(1'h0)] wire309;
  wire signed [(4'h8):(1'h0)] wire308;
  reg [(4'h8):(1'h0)] reg307 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg306 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg305 = (1'h0);
  reg [(4'h9):(1'h0)] reg304 = (1'h0);
  reg [(5'h11):(1'h0)] reg303 = (1'h0);
  reg [(4'he):(1'h0)] reg302 = (1'h0);
  reg [(4'hc):(1'h0)] reg301 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg300 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg299 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg298 = (1'h0);
  reg [(5'h11):(1'h0)] reg297 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg296 = (1'h0);
  reg [(5'h12):(1'h0)] reg295 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg294 = (1'h0);
  reg [(5'h15):(1'h0)] reg293 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg291 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire290;
  wire [(3'h7):(1'h0)] wire289;
  wire signed [(2'h3):(1'h0)] wire288;
  reg signed [(4'hf):(1'h0)] reg287 = (1'h0);
  reg [(2'h3):(1'h0)] reg286 = (1'h0);
  reg [(5'h10):(1'h0)] reg285 = (1'h0);
  reg [(2'h3):(1'h0)] reg284 = (1'h0);
  reg [(4'hc):(1'h0)] reg283 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg282 = (1'h0);
  reg [(4'hb):(1'h0)] reg281 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire280;
  wire signed [(3'h4):(1'h0)] wire279;
  wire [(4'h9):(1'h0)] wire278;
  wire [(3'h4):(1'h0)] wire277;
  reg signed [(5'h15):(1'h0)] reg276 = (1'h0);
  reg signed [(4'he):(1'h0)] reg275 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg274 = (1'h0);
  reg [(5'h11):(1'h0)] reg273 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg272 = (1'h0);
  reg [(3'h7):(1'h0)] reg271 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg269 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg268 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg267 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg266 = (1'h0);
  reg [(5'h14):(1'h0)] reg265 = (1'h0);
  reg [(5'h14):(1'h0)] reg264 = (1'h0);
  reg [(4'ha):(1'h0)] reg263 = (1'h0);
  reg signed [(4'he):(1'h0)] reg262 = (1'h0);
  reg [(4'hd):(1'h0)] reg261 = (1'h0);
  reg [(4'hf):(1'h0)] reg260 = (1'h0);
  reg [(5'h15):(1'h0)] reg259 = (1'h0);
  reg [(5'h10):(1'h0)] reg258 = (1'h0);
  reg [(5'h15):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg256 = (1'h0);
  wire [(4'hc):(1'h0)] wire255;
  wire [(5'h12):(1'h0)] wire254;
  reg [(4'hb):(1'h0)] reg253 = (1'h0);
  reg [(2'h2):(1'h0)] reg252 = (1'h0);
  reg [(5'h11):(1'h0)] reg251 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg250 = (1'h0);
  reg [(5'h11):(1'h0)] reg249 = (1'h0);
  reg [(3'h5):(1'h0)] reg248 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg246 = (1'h0);
  wire [(3'h5):(1'h0)] wire245;
  wire signed [(4'h8):(1'h0)] wire244;
  assign y = {wire315,
                 reg314,
                 reg313,
                 reg312,
                 wire311,
                 wire310,
                 wire309,
                 wire308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 wire290,
                 wire289,
                 wire288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 wire280,
                 wire279,
                 wire278,
                 wire277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 wire255,
                 wire254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 wire245,
                 wire244,
                 (1'h0)};
  assign wire244 = (wire242[(1'h1):(1'h1)] ?
                       ($signed(wire240) ^~ {$signed((&(8'hb9)))}) : $unsigned((^$signed((^wire241)))));
  assign wire245 = (~|$unsigned($signed(((wire243 ^~ wire244) << (~|wire244)))));
  always
    @(posedge clk) begin
      if (((-$unsigned(wire245)) ? $signed((8'hbf)) : wire245))
        begin
          reg246 <= ((wire243 ?
              (~|((-wire243) + (wire244 ?
                  wire243 : wire243))) : ($unsigned({(8'ha9), wire243}) ?
                  $unsigned($signed(wire241)) : ((-(7'h40)) | (wire244 | wire242)))) ~^ wire242);
          reg247 <= (($unsigned(wire242[(3'h4):(1'h0)]) == $unsigned({$unsigned((8'hbc)),
                  (^wire241)})) ?
              wire240 : $unsigned(wire241[(3'h6):(2'h3)]));
          reg248 <= (!(($unsigned($unsigned(wire243)) >>> ($signed((8'hac)) > $unsigned(reg247))) <= $unsigned(wire244[(2'h3):(1'h0)])));
        end
      else
        begin
          if (wire244[(2'h3):(1'h0)])
            begin
              reg246 <= (reg246[(4'hc):(4'h8)] || (8'hb1));
              reg247 <= wire241;
            end
          else
            begin
              reg246 <= ({$unsigned({$unsigned(wire243)}),
                      wire242[(3'h5):(3'h4)]} ?
                  (($signed((!wire245)) << (~|$unsigned((8'hb4)))) ?
                      wire240 : wire241[(1'h1):(1'h0)]) : (-reg247[(1'h1):(1'h0)]));
              reg247 <= wire241;
              reg248 <= ($signed($signed(((-(7'h42)) ?
                      (reg246 != (8'hb9)) : $unsigned(reg246)))) ?
                  ((8'hb8) ?
                      $signed($unsigned((wire241 ?
                          (7'h41) : reg247))) : reg247[(3'h5):(2'h3)]) : wire243);
              reg249 <= $unsigned(wire240[(1'h0):(1'h0)]);
            end
        end
      reg250 <= $signed(wire244);
      if (((^wire245[(2'h3):(2'h2)]) ? wire240[(4'hc):(1'h1)] : (7'h42)))
        begin
          reg251 <= (&(-($unsigned($signed(wire245)) ?
              {$unsigned((8'hab))} : $signed($signed(wire243)))));
        end
      else
        begin
          reg251 <= $signed((({$signed(reg248),
              $unsigned(wire244)} && ($signed(wire241) ?
              (reg249 ?
                  wire242 : reg246) : (!reg249))) != wire245[(1'h0):(1'h0)]));
        end
      reg252 <= reg250;
      reg253 <= (wire243[(4'he):(4'hb)] >= (reg250 >= (~^(((8'h9e) & reg250) ?
          ((8'hb8) ? reg246 : reg251) : (^~(8'hb5))))));
    end
  assign wire254 = $signed(({(!wire244[(1'h0):(1'h0)]),
                           (reg249 + (wire244 <= reg247))} ?
                       reg248[(2'h3):(2'h3)] : (-{$signed(reg248)})));
  assign wire255 = {($unsigned((&(8'ha3))) ?
                           $unsigned(((reg253 == reg246) | (wire241 ?
                               wire244 : reg251))) : reg249[(5'h11):(2'h3)])};
  always
    @(posedge clk) begin
      reg256 <= $unsigned((reg247[(4'h8):(3'h6)] ?
          $signed((((8'hb2) > wire240) == $unsigned(wire242))) : reg253[(3'h7):(1'h0)]));
      if (($unsigned(wire244) ?
          ((($signed(reg251) | (reg246 | reg247)) ?
              (((7'h43) | wire254) ^ $signed((7'h40))) : reg253) * (&(~&wire242))) : $unsigned((reg250 != ((reg251 ?
              (8'h9f) : reg253) * {wire255})))))
        begin
          reg257 <= wire245;
          reg258 <= (^~wire244[(2'h2):(1'h0)]);
          if (((~^$unsigned(wire255[(1'h0):(1'h0)])) ^~ $unsigned(wire243[(2'h3):(2'h2)])))
            begin
              reg259 <= (~|(!reg252));
            end
          else
            begin
              reg259 <= (($unsigned(wire241) ^~ ({(reg257 ? reg251 : (7'h44)),
                      $signed(wire255)} >= (+((8'hb5) ? reg256 : (8'hb1))))) ?
                  ((8'haa) ?
                      wire241 : $signed($signed((reg253 >> reg250)))) : (~&wire244));
              reg260 <= ({$unsigned(($unsigned(reg257) | wire255)),
                      ({$unsigned(wire244), reg248[(2'h3):(2'h2)]} ?
                          $unsigned($signed(wire255)) : reg246)} ?
                  reg256 : $signed(((-$signed((7'h43))) ?
                      $unsigned((8'hb4)) : (reg257[(3'h6):(1'h0)] ~^ $unsigned(reg256)))));
              reg261 <= $unsigned((!((((8'hb1) | wire254) - $unsigned(wire255)) ?
                  $signed((8'h9c)) : $unsigned((^reg257)))));
            end
          if ({((-$unsigned($unsigned(reg248))) <<< (reg258[(3'h7):(2'h2)] & wire245)),
              ((reg261 ? {(-reg248)} : reg260) ?
                  $unsigned(reg253[(4'hb):(4'ha)]) : reg248)})
            begin
              reg262 <= $unsigned(reg250);
              reg263 <= reg247[(2'h2):(1'h0)];
              reg264 <= (wire244 >= reg262);
            end
          else
            begin
              reg262 <= $unsigned(reg264);
              reg263 <= ($unsigned(wire242[(2'h2):(2'h2)]) ?
                  reg258 : (~(((wire240 ? reg249 : reg246) ?
                          reg249[(4'hb):(4'h9)] : ((8'ha4) ?
                              wire255 : reg259)) ?
                      {(wire243 ~^ reg262)} : $signed($signed((8'hb1))))));
              reg264 <= ($signed(wire245) < {(reg251 == {$signed((8'ha5))})});
              reg265 <= ({$signed(wire254),
                  (wire245[(3'h4):(2'h2)] | $signed(((8'hb5) <<< reg246)))} == reg257[(4'ha):(2'h3)]);
            end
          reg266 <= $unsigned($unsigned((($unsigned((7'h44)) <<< (8'hb0)) ~^ reg248)));
        end
      else
        begin
          reg257 <= $signed({$signed($unsigned($unsigned(reg266))),
              wire245[(3'h5):(1'h0)]});
          reg258 <= {(($signed({(8'had), reg250}) ?
                  reg259 : $unsigned(wire240)) > (~|$unsigned((&reg266)))),
              ({(reg246[(2'h3):(2'h2)] < reg256[(2'h2):(1'h0)]),
                      $unsigned((reg248 ? wire245 : wire255))} ?
                  $signed((8'ha7)) : ((~^$unsigned(wire240)) ?
                      reg266[(1'h0):(1'h0)] : reg257[(4'hf):(1'h0)]))};
          if (((!(&$signed((reg259 < reg258)))) ?
              reg256[(5'h10):(3'h6)] : ($signed((&(reg256 | reg264))) - ((|(reg258 & reg252)) ?
                  reg249[(4'h9):(4'h8)] : (((7'h44) <<< reg252) ?
                      {reg253} : reg261[(1'h0):(1'h0)])))))
            begin
              reg259 <= {((!(wire242 ?
                      (|reg257) : (reg248 ?
                          reg248 : (8'hab)))) || reg248[(1'h1):(1'h0)]),
                  $signed((reg259[(5'h12):(2'h3)] ?
                      reg261[(4'ha):(1'h0)] : ({(8'hb7)} ?
                          $unsigned((7'h43)) : wire242)))};
              reg260 <= $signed(reg252);
            end
          else
            begin
              reg259 <= reg250[(4'hd):(3'h6)];
              reg260 <= $signed((wire242 ?
                  (-(reg263[(4'ha):(2'h3)] ?
                      $unsigned(reg260) : (~|wire240))) : reg262[(4'hc):(1'h1)]));
            end
          reg261 <= $signed(wire241);
          if (reg251[(2'h3):(1'h0)])
            begin
              reg262 <= $signed(wire240[(3'h6):(3'h4)]);
              reg263 <= $unsigned($signed(wire243[(4'hb):(3'h5)]));
            end
          else
            begin
              reg262 <= $signed(reg266[(4'h9):(3'h4)]);
              reg263 <= (wire254 || {reg257, reg256});
            end
        end
      reg267 <= (~^($unsigned(wire245) < $unsigned($unsigned((&reg257)))));
      if (reg260)
        begin
          reg268 <= ((reg246 >= ($unsigned((wire244 * (8'hbd))) ?
              reg261 : ($unsigned(wire255) >> (wire241 != (7'h43))))) > (+reg260[(3'h5):(3'h5)]));
          reg269 <= $unsigned(wire244);
          reg270 <= {(-reg266[(1'h1):(1'h1)]),
              (^~$signed((reg264 & ((8'ha0) ? reg250 : reg268))))};
        end
      else
        begin
          if ((($unsigned(reg259[(5'h12):(4'hb)]) ?
              {{(~(8'hb6))}} : (8'hb2)) || $signed(reg268[(1'h1):(1'h1)])))
            begin
              reg268 <= wire254;
            end
          else
            begin
              reg268 <= {$signed(reg269[(4'hb):(3'h7)])};
              reg269 <= (^(reg259 ?
                  $unsigned($unsigned($signed((8'had)))) : $signed(((reg259 ?
                      (8'hb1) : (8'hbc)) < wire245[(1'h1):(1'h0)]))));
              reg270 <= wire254[(2'h2):(2'h2)];
            end
          if ($signed((wire254[(3'h7):(1'h0)] ?
              $signed($unsigned((reg261 ?
                  reg258 : reg265))) : $signed(((wire245 ? wire241 : reg261) ?
                  (reg269 - reg250) : (reg252 ? reg256 : reg269))))))
            begin
              reg271 <= wire243[(4'h8):(2'h2)];
              reg272 <= {(^($unsigned((reg251 ? reg260 : reg262)) ?
                      {$signed(wire245),
                          $unsigned((7'h43))} : {$signed(reg261)}))};
              reg273 <= (^~reg248);
              reg274 <= $signed((!($unsigned(reg263) ?
                  {(wire244 ? wire241 : (7'h43)),
                      (reg247 ? reg252 : wire242)} : (8'ha4))));
            end
          else
            begin
              reg271 <= reg248;
            end
          reg275 <= $unsigned(reg246[(4'ha):(2'h2)]);
        end
      reg276 <= $signed((~|{$signed(reg265[(3'h5):(2'h2)])}));
    end
  assign wire277 = $unsigned($signed((&(!reg264[(5'h13):(4'hf)]))));
  assign wire278 = ($unsigned((reg264[(4'hd):(4'h9)] ^ reg275)) << ($signed((reg265[(5'h12):(3'h5)] && $signed(wire240))) >>> $unsigned((!(~&reg258)))));
  assign wire279 = ((($signed($signed(reg272)) == reg261[(3'h4):(1'h0)]) >= $signed((-(reg256 ?
                           reg264 : reg275)))) ?
                       (8'h9d) : (!wire277[(2'h3):(1'h1)]));
  assign wire280 = reg265;
  always
    @(posedge clk) begin
      reg281 <= $unsigned((wire243[(2'h3):(2'h2)] ?
          {reg252} : (-({reg256} ? wire255 : (~reg258)))));
      if ({(|(reg257 ? (wire241 <= (|reg269)) : (&(wire280 && reg262)))),
          ($unsigned({(reg253 && reg263), $signed(reg259)}) ?
              (!reg250) : $unsigned(reg249))})
        begin
          reg282 <= reg260[(2'h2):(1'h1)];
          reg283 <= $signed(wire254);
          reg284 <= (^(|(!reg276)));
        end
      else
        begin
          reg282 <= {$unsigned((~^$unsigned(reg262)))};
        end
      if ((&reg275[(4'ha):(2'h3)]))
        begin
          if ((reg276[(3'h5):(2'h2)] ?
              reg273[(4'hf):(3'h6)] : reg275[(4'he):(1'h1)]))
            begin
              reg285 <= ((&(reg283[(2'h2):(1'h1)] ?
                      ($unsigned(wire279) != ((7'h43) ?
                          reg262 : reg274)) : reg247)) ?
                  reg249 : (reg261[(3'h4):(2'h2)] != ((((8'hac) ?
                      reg253 : reg267) | (reg269 ?
                      reg257 : wire243)) != (reg274 ?
                      wire244 : $unsigned(reg251)))));
            end
          else
            begin
              reg285 <= $unsigned(reg256);
            end
          reg286 <= $unsigned(($signed(reg262[(4'h8):(2'h2)]) ?
              (~reg246[(4'h8):(3'h7)]) : (-$unsigned((reg246 <<< reg251)))));
          reg287 <= reg286[(2'h3):(1'h0)];
        end
      else
        begin
          reg285 <= ((-$unsigned({(~wire242)})) ? wire278 : reg269);
          reg286 <= {$unsigned((($signed(reg250) ^ (~&reg251)) >= ((wire241 ~^ reg273) < {reg282})))};
          reg287 <= ({wire243[(5'h10):(2'h3)]} || wire243);
        end
    end
  assign wire288 = ($signed(wire243) >= ($unsigned(($signed(reg268) ^~ (wire241 >= reg286))) ?
                       reg266 : (!(wire255 ?
                           $signed(wire278) : reg276[(5'h15):(1'h1)]))));
  assign wire289 = (^(reg266 != {(~(reg287 ? reg282 : reg260))}));
  assign wire290 = $unsigned(((^~reg262[(1'h1):(1'h0)]) >>> (reg252[(1'h0):(1'h0)] ?
                       $signed(reg270[(1'h0):(1'h0)]) : (8'h9f))));
  always
    @(posedge clk) begin
      reg291 <= (+reg283[(3'h5):(2'h2)]);
      if ({reg252})
        begin
          reg292 <= (reg259[(1'h0):(1'h0)] == reg264);
          reg293 <= {(-(reg271[(1'h1):(1'h1)] ?
                  $signed(wire288) : $unsigned($signed((8'hbc))))),
              ((-(wire279 - reg262[(3'h6):(3'h6)])) ?
                  (wire277 == ((wire279 <= reg258) ?
                      $signed((8'hb3)) : {reg291, reg251})) : (((~wire240) ?
                      $unsigned(reg264) : (~wire254)) + (8'hb1)))};
        end
      else
        begin
          reg292 <= {{$signed(reg281[(2'h3):(1'h1)])},
              (reg286[(1'h1):(1'h1)] ?
                  ($signed($unsigned(reg257)) ~^ {(8'ha4)}) : {(^~wire254),
                      ({reg261, reg273} ? (~^reg283) : reg248)})};
        end
      reg294 <= {((~|$signed((wire244 < reg253))) ?
              ($signed($unsigned(reg292)) ?
                  reg246 : {$signed(reg251), reg286}) : (+{reg252})),
          reg285};
    end
  always
    @(posedge clk) begin
      if (reg256)
        begin
          reg295 <= ((~{reg260[(4'hf):(4'ha)]}) ^~ (7'h43));
          if ((~$signed((-(^{reg287, reg276})))))
            begin
              reg296 <= reg251;
              reg297 <= $signed(reg260[(3'h5):(2'h2)]);
              reg298 <= $signed(reg249[(3'h5):(3'h5)]);
            end
          else
            begin
              reg296 <= $unsigned((reg260[(3'h5):(3'h5)] & reg266));
              reg297 <= {{(reg251[(1'h1):(1'h1)] ?
                          ($signed(reg296) ?
                              (&reg296) : (reg260 ^~ wire255)) : ($signed(wire278) ?
                              $unsigned(reg287) : (reg276 ? wire289 : reg275))),
                      reg250}};
              reg298 <= $signed((8'ha7));
              reg299 <= wire245[(1'h1):(1'h0)];
              reg300 <= ($signed((wire288[(2'h3):(2'h3)] != reg298[(4'hd):(3'h6)])) ~^ $unsigned((&{reg297[(4'hc):(3'h6)],
                  wire255[(2'h2):(2'h2)]})));
            end
          reg301 <= $signed(reg292);
        end
      else
        begin
          if ($unsigned($unsigned((^~reg295))))
            begin
              reg295 <= (~&({$unsigned(((8'hb3) ? wire242 : reg271)),
                  $signed((reg257 ?
                      (8'ha4) : (8'ha3)))} & $unsigned((reg276[(4'h9):(3'h5)] && wire280))));
              reg296 <= $unsigned((~&$signed((~^reg298[(4'hb):(4'hb)]))));
              reg297 <= $unsigned($signed((-(!(reg248 >= reg285)))));
              reg298 <= ((&(~|$unsigned((wire245 > wire289)))) + $signed(reg263[(1'h0):(1'h0)]));
              reg299 <= {$unsigned($unsigned($unsigned((~^reg295))))};
            end
          else
            begin
              reg295 <= reg256;
              reg296 <= reg294[(4'h8):(3'h5)];
              reg297 <= wire289[(3'h6):(1'h1)];
              reg298 <= (~|reg281[(3'h6):(1'h1)]);
            end
        end
      if ($unsigned((~$unsigned($signed($signed(wire290))))))
        begin
          reg302 <= $unsigned(reg262);
          reg303 <= wire244[(1'h0):(1'h0)];
          reg304 <= (~reg261);
          reg305 <= (reg292[(2'h3):(2'h3)] ?
              wire242[(3'h4):(1'h1)] : (~|($unsigned({reg266}) && reg248)));
          if ($signed({reg305}))
            begin
              reg306 <= {((((^reg295) >= $unsigned(wire280)) | (~|reg268)) ?
                      $signed(wire245[(2'h2):(1'h1)]) : $unsigned(reg302))};
            end
          else
            begin
              reg306 <= (~&($unsigned(wire279) ?
                  reg275[(4'hd):(1'h1)] : ($unsigned(reg302) ?
                      (reg269 - $signed(wire242)) : ($signed(reg300) ?
                          $unsigned(wire289) : reg299))));
              reg307 <= (-((8'hbb) << {reg284[(2'h2):(1'h1)],
                  wire279[(1'h0):(1'h0)]}));
            end
        end
      else
        begin
          if (reg257)
            begin
              reg302 <= {$signed((!(wire289 ?
                      (wire240 ? reg300 : (8'ha4)) : (wire288 ?
                          wire245 : reg275)))),
                  (^~reg259)};
              reg303 <= (!{(reg291 > reg307[(2'h3):(1'h0)])});
            end
          else
            begin
              reg302 <= {$signed({(reg299[(2'h2):(1'h1)] ?
                          {reg248, (8'haf)} : (8'ha3)),
                      (((8'h9f) ? reg263 : reg291) ? (^wire241) : wire280)}),
                  (wire290[(1'h0):(1'h0)] ?
                      $signed(({reg286, reg276} ?
                          (wire289 ~^ reg286) : (~^wire277))) : $signed($unsigned((wire242 <<< reg303))))};
              reg303 <= {(-reg267[(2'h3):(2'h3)]), (8'hb7)};
            end
        end
    end
  assign wire308 = (((~|reg248[(2'h2):(1'h1)]) ?
                       reg275 : reg246) <<< {$signed(reg307[(4'h8):(1'h0)])});
  assign wire309 = (~|(~|(reg286 || $unsigned($signed((8'hae))))));
  assign wire310 = {$unsigned(reg248[(2'h2):(2'h2)])};
  assign wire311 = (&reg272[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg312 <= (!(^~$unsigned((~&$unsigned(reg273)))));
      reg313 <= reg302[(2'h2):(1'h1)];
      reg314 <= (!(reg313 >>> $unsigned(wire308[(2'h3):(1'h1)])));
    end
  assign wire315 = $signed((wire290[(4'h9):(4'h8)] >= reg272[(1'h0):(1'h0)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module346
#( parameter param386 = ((+(~|({(8'hab), (8'ha8)} != {(8'hbb), (8'had)}))) * (^~(8'hbe)))
, parameter param387 = param386 )
(y, clk, wire350, wire349, wire348, wire347);
  output wire [(32'h184):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire350;
  input wire [(4'ha):(1'h0)] wire349;
  input wire [(5'h12):(1'h0)] wire348;
  input wire signed [(2'h2):(1'h0)] wire347;
  reg signed [(4'h9):(1'h0)] reg385 = (1'h0);
  reg signed [(4'he):(1'h0)] reg384 = (1'h0);
  reg [(5'h11):(1'h0)] reg383 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg382 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg381 = (1'h0);
  reg [(5'h13):(1'h0)] reg380 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg379 = (1'h0);
  reg [(2'h2):(1'h0)] reg378 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg377 = (1'h0);
  reg [(3'h5):(1'h0)] reg376 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg375 = (1'h0);
  reg [(4'hd):(1'h0)] reg374 = (1'h0);
  reg [(3'h7):(1'h0)] reg373 = (1'h0);
  reg [(4'hf):(1'h0)] reg372 = (1'h0);
  wire [(4'ha):(1'h0)] wire371;
  wire signed [(4'ha):(1'h0)] wire370;
  wire [(5'h12):(1'h0)] wire369;
  wire signed [(5'h13):(1'h0)] wire368;
  wire [(4'he):(1'h0)] wire367;
  wire signed [(3'h6):(1'h0)] wire366;
  reg [(4'hd):(1'h0)] reg365 = (1'h0);
  wire [(5'h11):(1'h0)] wire364;
  reg signed [(4'h9):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg362 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg361 = (1'h0);
  reg [(5'h11):(1'h0)] reg360 = (1'h0);
  reg [(3'h4):(1'h0)] reg359 = (1'h0);
  reg [(4'h9):(1'h0)] reg358 = (1'h0);
  reg [(5'h12):(1'h0)] reg357 = (1'h0);
  reg [(3'h7):(1'h0)] reg356 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg355 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg354 = (1'h0);
  reg [(2'h3):(1'h0)] reg353 = (1'h0);
  reg [(3'h5):(1'h0)] reg352 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg351 = (1'h0);
  assign y = {reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 wire371,
                 wire370,
                 wire369,
                 wire368,
                 wire367,
                 wire366,
                 reg365,
                 wire364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg351 <= $signed($unsigned($signed(({wire349, (8'hae)} ^ (8'hb5)))));
      if (wire349)
        begin
          if ($signed(wire349[(3'h6):(1'h0)]))
            begin
              reg352 <= wire350;
              reg353 <= (wire349[(3'h7):(1'h1)] ?
                  (^(^({wire347, wire349} ?
                      wire348[(3'h5):(2'h3)] : $unsigned(reg352)))) : (($unsigned($signed(wire350)) < wire348) - wire347[(1'h1):(1'h1)]));
            end
          else
            begin
              reg352 <= (reg351 ?
                  $unsigned((~&reg351[(3'h6):(1'h1)])) : wire348);
              reg353 <= reg353;
              reg354 <= $signed((8'ha2));
              reg355 <= (reg351 ?
                  ($signed((((8'ha1) >> wire347) & (|(8'ha5)))) ?
                      {((wire347 - wire350) <<< (8'ha1))} : $signed((8'ha2))) : (wire349[(4'h8):(3'h4)] - reg351));
              reg356 <= ((8'hb0) ?
                  $unsigned(wire349) : ($unsigned(reg354[(1'h1):(1'h1)]) ^ (reg354 || (~^(wire347 ?
                      reg351 : wire350)))));
            end
          reg357 <= wire347;
          reg358 <= $signed(wire348);
          if ($signed(reg355))
            begin
              reg359 <= reg358[(4'h8):(4'h8)];
              reg360 <= wire350;
            end
          else
            begin
              reg359 <= {(~&(^~reg352))};
              reg360 <= reg354;
              reg361 <= (wire347 || reg352);
              reg362 <= (8'hbf);
              reg363 <= reg352[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg352 <= reg354;
          reg353 <= {(reg352[(2'h3):(2'h2)] & reg359[(2'h2):(1'h1)]),
              wire349[(4'h8):(4'h8)]};
          reg354 <= reg355[(2'h3):(1'h1)];
        end
    end
  assign wire364 = $unsigned(reg352[(2'h2):(1'h0)]);
  always
    @(posedge clk) begin
      reg365 <= $unsigned((~^(reg363[(4'h9):(2'h2)] >= reg361[(4'h9):(1'h1)])));
    end
  assign wire366 = reg363[(4'h8):(2'h2)];
  assign wire367 = (~|$signed(reg352[(3'h4):(2'h3)]));
  assign wire368 = ($signed((~^$signed({wire366, reg358}))) ?
                       ((((reg357 ? wire348 : reg357) ^ $unsigned(reg353)) ?
                               $signed(wire349) : ({reg363} ?
                                   $signed(reg353) : reg354)) ?
                           ({(~reg362)} ?
                               {$signed(reg361),
                                   $signed(reg351)} : ((~reg363) ^~ $unsigned(wire367))) : reg362[(2'h3):(1'h1)]) : {$signed($unsigned(wire366)),
                           $signed(reg365)});
  assign wire369 = wire347;
  assign wire370 = ((($signed((8'hbf)) ?
                       (&wire366) : reg363) == wire350) >= reg359);
  assign wire371 = $unsigned(reg354);
  always
    @(posedge clk) begin
      reg372 <= (({{(8'hbf),
              $signed(wire364)}} == wire367) ~^ (reg356[(3'h4):(2'h3)] ?
          ($unsigned(wire366[(3'h6):(3'h4)]) >>> wire370[(2'h2):(1'h0)]) : (-(reg363 ~^ (~&(7'h43))))));
      reg373 <= $signed({$unsigned($unsigned($unsigned((8'hb0))))});
      if ({$unsigned(wire367[(4'h9):(2'h3)])})
        begin
          reg374 <= (|reg360[(4'hc):(4'h8)]);
          reg375 <= {(reg356[(3'h6):(2'h2)] - reg362)};
          if (wire371[(4'h8):(1'h0)])
            begin
              reg376 <= {$unsigned({((reg359 << reg372) ?
                          (^~(8'ha2)) : reg375[(3'h6):(2'h3)])}),
                  reg361[(1'h1):(1'h1)]};
              reg377 <= reg354;
              reg378 <= (-$signed(($unsigned(reg362) ?
                  (~^reg355) : wire366[(1'h0):(1'h0)])));
              reg379 <= reg352;
              reg380 <= wire371;
            end
          else
            begin
              reg376 <= (wire366[(2'h2):(2'h2)] ?
                  wire369[(5'h10):(4'h8)] : {$unsigned(reg352[(1'h1):(1'h0)]),
                      $signed(({reg373} ? (~^reg378) : (^~(7'h42))))});
              reg377 <= reg380[(3'h5):(2'h2)];
              reg378 <= $signed((wire347[(1'h1):(1'h0)] >> $signed(reg365)));
              reg379 <= {$unsigned($unsigned((8'ha8)))};
            end
          if ((reg351 ?
              $unsigned((-$signed(((8'hb6) ?
                  wire350 : reg376)))) : reg358[(2'h2):(2'h2)]))
            begin
              reg381 <= (-($signed(((reg357 ?
                      (8'hbe) : reg362) & $unsigned((8'hb3)))) ?
                  $signed({((7'h40) ^ wire364)}) : wire367[(4'h8):(3'h7)]));
              reg382 <= $signed({{($signed(reg356) ?
                          $unsigned(reg355) : wire369),
                      (!reg356)},
                  $signed(wire350[(3'h7):(1'h1)])});
              reg383 <= $unsigned($unsigned($unsigned(((reg374 ~^ (8'hab)) ^ (!wire347)))));
            end
          else
            begin
              reg381 <= $signed(reg363);
              reg382 <= reg365;
              reg383 <= $signed(reg372);
              reg384 <= reg375;
              reg385 <= ((reg376[(3'h4):(2'h2)] ?
                  (-$unsigned(wire348[(5'h11):(1'h0)])) : {$unsigned($signed(reg377))}) * reg376);
            end
        end
      else
        begin
          if ($unsigned({$signed({(~|(8'hbe)), reg353})}))
            begin
              reg374 <= (reg376[(1'h0):(1'h0)] ~^ (($signed((reg356 ?
                          reg374 : reg378)) ?
                      wire369 : $signed((reg359 ^ reg360))) ?
                  wire348[(4'hc):(1'h0)] : (-reg354)));
              reg375 <= $signed($unsigned($unsigned($signed(reg359))));
              reg376 <= ($signed((8'h9c)) ?
                  wire370[(3'h6):(2'h2)] : ({reg384} ^ ($unsigned(reg383[(2'h2):(1'h1)]) ?
                      {wire349[(2'h2):(1'h0)],
                          (reg353 >>> reg374)} : wire371[(3'h7):(3'h4)])));
              reg377 <= reg382[(3'h7):(1'h1)];
            end
          else
            begin
              reg374 <= $signed((((reg354[(1'h1):(1'h1)] && {reg374}) ?
                      ((wire347 >> reg379) ?
                          (^~reg385) : $unsigned(reg365)) : reg365[(2'h2):(1'h1)]) ?
                  reg373 : $unsigned((reg373 != (!reg378)))));
              reg375 <= reg378;
              reg376 <= $unsigned((^(~^(!(reg356 << wire369)))));
              reg377 <= $signed({reg376[(2'h2):(1'h0)], reg354});
              reg378 <= $signed((^~$unsigned((+reg362[(1'h0):(1'h0)]))));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module420
#( parameter param613 = (!(((&(^~(8'hb4))) ? (((8'hb8) ? (8'hbf) : (8'ha4)) ? (8'ha0) : ((8'ha0) ? (8'hb1) : (8'h9d))) : ({(8'h9c), (8'haa)} - ((8'hb1) > (8'hb1)))) & {(^~{(8'hb6)})})) )
(y, clk, wire425, wire424, wire423, wire422, wire421);
  output wire [(32'h2fb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire425;
  input wire [(4'hd):(1'h0)] wire424;
  input wire [(5'h11):(1'h0)] wire423;
  input wire [(4'h8):(1'h0)] wire422;
  input wire signed [(5'h14):(1'h0)] wire421;
  wire [(4'he):(1'h0)] wire612;
  reg [(5'h11):(1'h0)] reg611 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire610;
  reg [(4'h8):(1'h0)] reg609 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg608 = (1'h0);
  reg [(3'h5):(1'h0)] reg607 = (1'h0);
  reg [(4'hf):(1'h0)] reg606 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg605 = (1'h0);
  reg [(5'h14):(1'h0)] reg604 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire602;
  wire signed [(4'he):(1'h0)] wire558;
  wire [(3'h4):(1'h0)] wire557;
  wire [(4'h9):(1'h0)] wire556;
  wire signed [(4'hf):(1'h0)] wire555;
  wire signed [(5'h15):(1'h0)] wire554;
  wire [(2'h3):(1'h0)] wire552;
  wire [(4'h9):(1'h0)] wire478;
  reg [(2'h3):(1'h0)] reg477 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg476 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg475 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg474 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg473 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg472 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg471 = (1'h0);
  reg [(4'hc):(1'h0)] reg470 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg469 = (1'h0);
  wire [(3'h4):(1'h0)] wire468;
  reg signed [(2'h3):(1'h0)] reg467 = (1'h0);
  reg [(5'h11):(1'h0)] reg466 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg465 = (1'h0);
  reg [(3'h4):(1'h0)] reg464 = (1'h0);
  reg [(4'he):(1'h0)] reg463 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg462 = (1'h0);
  reg [(5'h12):(1'h0)] reg461 = (1'h0);
  reg [(4'ha):(1'h0)] reg460 = (1'h0);
  reg [(4'hc):(1'h0)] reg459 = (1'h0);
  reg [(2'h2):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg457 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg456 = (1'h0);
  reg [(4'hb):(1'h0)] reg455 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg453 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg452 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg451 = (1'h0);
  reg [(5'h15):(1'h0)] reg450 = (1'h0);
  reg [(5'h14):(1'h0)] reg449 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire448;
  reg [(4'hd):(1'h0)] reg447 = (1'h0);
  reg [(4'ha):(1'h0)] reg446 = (1'h0);
  reg [(2'h3):(1'h0)] reg445 = (1'h0);
  reg [(5'h10):(1'h0)] reg444 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg443 = (1'h0);
  reg [(3'h4):(1'h0)] reg442 = (1'h0);
  reg [(4'h9):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg440 = (1'h0);
  reg [(4'hf):(1'h0)] reg439 = (1'h0);
  reg [(5'h11):(1'h0)] reg438 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg437 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg436 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg435 = (1'h0);
  reg [(4'ha):(1'h0)] reg434 = (1'h0);
  reg [(5'h12):(1'h0)] reg433 = (1'h0);
  reg [(4'h9):(1'h0)] reg432 = (1'h0);
  reg [(5'h10):(1'h0)] reg431 = (1'h0);
  reg [(2'h3):(1'h0)] reg430 = (1'h0);
  reg [(4'hb):(1'h0)] reg429 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg428 = (1'h0);
  reg [(3'h6):(1'h0)] reg427 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire426;
  assign y = {wire612,
                 reg611,
                 wire610,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 wire602,
                 wire558,
                 wire557,
                 wire556,
                 wire555,
                 wire554,
                 wire552,
                 wire478,
                 reg477,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 reg469,
                 wire468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 wire448,
                 reg447,
                 reg446,
                 reg445,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 wire426,
                 (1'h0)};
  assign wire426 = {(|wire421)};
  always
    @(posedge clk) begin
      reg427 <= ($unsigned($signed(wire426)) ?
          wire425[(4'hd):(4'h8)] : $signed(((!wire423[(4'hb):(4'h9)]) || $signed((wire421 & wire426)))));
      if ({{wire421}})
        begin
          reg428 <= reg427;
          if ($unsigned($signed(wire425)))
            begin
              reg429 <= $unsigned($unsigned((!wire421[(4'h9):(4'h8)])));
              reg430 <= $unsigned(($signed($signed($signed(reg429))) >> ({(^~wire425),
                  ((8'hb9) ? wire421 : (8'h9c))} >> reg429[(4'h9):(1'h1)])));
            end
          else
            begin
              reg429 <= ($unsigned($signed((~&(!wire424)))) >>> ((((wire425 ^ reg429) ?
                      $signed(wire426) : wire421) ?
                  (~^$signed(wire424)) : $unsigned(wire422)) >> $signed(((reg427 >>> reg428) ?
                  $unsigned(wire424) : reg428[(2'h2):(2'h2)]))));
            end
          reg431 <= reg428[(3'h4):(2'h2)];
        end
      else
        begin
          reg428 <= $unsigned(((8'ha6) ?
              ($signed($unsigned(wire422)) ?
                  (~&reg430) : $signed((8'hb0))) : $signed((8'hba))));
          reg429 <= reg431;
        end
      if ((wire424 ^ wire425[(4'h9):(2'h2)]))
        begin
          reg432 <= $unsigned((({$signed((8'hac))} ?
              reg431[(4'ha):(4'ha)] : $signed((reg430 == reg428))) <= $unsigned((reg430 | (reg428 * reg430)))));
          reg433 <= ($signed(wire425[(4'hf):(4'he)]) <= ((|(~^{wire422,
                  reg432})) ?
              $signed(($signed(wire421) == (-reg430))) : $unsigned($unsigned({(8'hbf),
                  reg432}))));
        end
      else
        begin
          reg432 <= $unsigned($signed(reg430));
          reg433 <= $unsigned($unsigned(wire425));
          reg434 <= $unsigned($signed((-reg430)));
          reg435 <= $unsigned({reg431, {(7'h42)}});
        end
      if ($unsigned(wire424))
        begin
          reg436 <= (reg431 < (~|({$signed(wire421)} ?
              ((wire425 ?
                  wire425 : wire422) >>> $unsigned(reg429)) : reg428[(1'h1):(1'h0)])));
          reg437 <= reg436;
          reg438 <= ((!(^~wire425)) ? wire426 : wire426[(1'h0):(1'h0)]);
        end
      else
        begin
          reg436 <= {(wire422 ?
                  $unsigned($signed((wire423 ? wire426 : wire425))) : ((8'ha2) ?
                      {{reg438},
                          $signed(reg437)} : ((7'h40) << (reg429 > reg434))))};
          if ((($unsigned($signed(((8'hae) <<< reg433))) ?
              reg430 : (($unsigned(reg430) ?
                  $unsigned(reg437) : (reg434 ?
                      (8'ha7) : wire421)) >> $signed($signed(reg431)))) | wire422[(1'h1):(1'h0)]))
            begin
              reg437 <= ($signed(($signed({wire421}) ?
                  (~^$signed(wire423)) : $unsigned(reg429[(2'h2):(2'h2)]))) + $signed($unsigned((reg427[(1'h1):(1'h1)] < reg435))));
              reg438 <= (-($signed($signed($signed(reg430))) << (reg430[(2'h2):(2'h2)] | wire425)));
            end
          else
            begin
              reg437 <= reg435[(3'h6):(2'h3)];
              reg438 <= wire424;
              reg439 <= $signed((-($signed((reg436 >> (8'hb8))) ?
                  (^~(|reg435)) : reg431[(4'hb):(1'h0)])));
              reg440 <= $signed($unsigned($unsigned((reg435 != wire426))));
              reg441 <= $unsigned((reg433[(5'h10):(4'hd)] ?
                  $signed($unsigned($unsigned((8'hba)))) : $signed($signed((!(8'h9d))))));
            end
          if ((-wire421))
            begin
              reg442 <= (reg440 ?
                  (((8'hb6) * reg427) ?
                      reg430[(2'h3):(1'h1)] : ($unsigned(((7'h41) ?
                          reg441 : wire425)) <= {(reg429 ? (7'h44) : wire425),
                          (^reg431)})) : (!$unsigned(reg438[(5'h11):(3'h6)])));
              reg443 <= reg441;
              reg444 <= (($signed(reg432[(2'h2):(2'h2)]) ^~ $unsigned($signed((wire421 ?
                  reg431 : reg434)))) || (-$signed((^~$unsigned(reg435)))));
              reg445 <= (wire424 ? reg440 : $unsigned((-reg427)));
              reg446 <= reg441[(3'h7):(3'h4)];
            end
          else
            begin
              reg442 <= wire426[(2'h2):(2'h2)];
              reg443 <= reg439[(4'hb):(4'h9)];
              reg444 <= $signed(reg432[(4'h9):(1'h0)]);
              reg445 <= reg436[(2'h2):(2'h2)];
            end
          reg447 <= $signed(((($signed((8'hbf)) + reg435) >> (reg444[(4'he):(4'hc)] & reg442)) ?
              ($signed($signed(reg439)) | ((wire421 > reg427) ?
                  (!wire425) : $unsigned(reg440))) : $signed((reg442 ?
                  (reg440 ? wire425 : (8'hb4)) : reg442))));
        end
    end
  assign wire448 = reg441[(4'h9):(1'h1)];
  always
    @(posedge clk) begin
      if ((-(($unsigned(reg439) ^~ $unsigned($signed(wire421))) >= reg431[(2'h2):(1'h0)])))
        begin
          if ((wire448[(2'h3):(2'h2)] ?
              (+reg437[(3'h4):(3'h4)]) : reg431[(3'h4):(3'h4)]))
            begin
              reg449 <= (wire448 > reg447[(4'ha):(3'h7)]);
              reg450 <= (reg444[(4'hd):(4'h8)] ?
                  $signed(((reg428 * $unsigned(reg432)) >>> ((wire424 ?
                          wire426 : reg440) ?
                      reg437 : reg431))) : reg434[(3'h5):(2'h2)]);
              reg451 <= reg445[(1'h1):(1'h0)];
              reg452 <= $signed($unsigned(reg451));
              reg453 <= $signed($unsigned($signed((7'h44))));
            end
          else
            begin
              reg449 <= reg450[(4'he):(3'h5)];
              reg450 <= reg445[(2'h2):(2'h2)];
            end
          reg454 <= $unsigned($signed(wire448[(2'h3):(2'h3)]));
          if ({(|(+$unsigned((^reg449))))})
            begin
              reg455 <= reg450;
            end
          else
            begin
              reg455 <= reg444;
              reg456 <= (wire422 ?
                  reg450 : ((8'hac) ?
                      {$unsigned($unsigned((7'h42))),
                          reg450[(4'h8):(3'h7)]} : reg434));
            end
          reg457 <= (-$signed((8'hb3)));
        end
      else
        begin
          if ((reg452[(1'h1):(1'h1)] ?
              $unsigned((~^(^~(^reg451)))) : $unsigned($signed(((reg445 >>> reg427) != (reg433 ?
                  reg439 : reg433))))))
            begin
              reg449 <= (8'ha9);
              reg450 <= reg446[(3'h6):(3'h6)];
              reg451 <= reg451;
              reg452 <= ((((~(reg455 ? reg450 : reg440)) ?
                  (~&(reg429 ? reg456 : reg434)) : ($signed(reg428) + ((8'had) ?
                      reg452 : reg429))) ^ (~|((reg436 >= wire425) ?
                  $unsigned(reg436) : {(7'h41), reg435}))) & reg428);
              reg453 <= (^reg437[(3'h5):(3'h5)]);
            end
          else
            begin
              reg449 <= (~|(~($signed((reg445 >= reg456)) ?
                  ({reg453} ?
                      {wire424,
                          (8'ha9)} : reg445) : ($unsigned(reg452) >>> $unsigned(reg457)))));
              reg450 <= (($unsigned(($signed(reg439) | {(7'h42),
                      (8'ha0)})) && (($signed((8'ha1)) ?
                      (reg441 ^~ reg443) : (reg445 ?
                          (7'h44) : reg434)) ~^ (reg452[(2'h2):(2'h2)] ?
                      (~^reg427) : reg444))) ?
                  (!{($unsigned(reg453) ?
                          reg447[(4'h8):(4'h8)] : $signed((8'had)))}) : $signed($signed(reg453[(4'h8):(2'h2)])));
              reg451 <= $unsigned((|reg438[(2'h2):(1'h1)]));
              reg452 <= $unsigned(reg454);
            end
          if (reg453)
            begin
              reg454 <= ({$signed((reg430[(1'h1):(1'h1)] ?
                          reg428 : {reg440, wire423}))} ?
                  reg441 : reg428[(4'hb):(1'h0)]);
              reg455 <= (reg428[(1'h0):(1'h0)] == reg437);
            end
          else
            begin
              reg454 <= $unsigned(wire421);
              reg455 <= $unsigned({$unsigned($unsigned($unsigned(wire422)))});
              reg456 <= {{reg452[(1'h0):(1'h0)]}};
              reg457 <= $unsigned((~{(reg446 == {reg444, reg457}),
                  ((reg432 + (8'ha8)) ?
                      wire425[(5'h14):(4'h9)] : ((8'hac) ?
                          reg428 : (8'hb5)))}));
            end
          reg458 <= $signed(reg440[(4'hb):(2'h2)]);
        end
      if (wire421)
        begin
          if (wire422[(2'h3):(2'h3)])
            begin
              reg459 <= (reg432[(3'h5):(2'h3)] ?
                  reg455[(1'h1):(1'h0)] : (~(8'hb5)));
              reg460 <= reg447[(3'h4):(2'h2)];
            end
          else
            begin
              reg459 <= (reg453[(5'h12):(4'hb)] <<< $signed((reg445[(2'h3):(1'h0)] < $signed({(7'h42),
                  (8'hb7)}))));
              reg460 <= reg453;
              reg461 <= $unsigned(((^~(reg433 ?
                  $unsigned((8'hb5)) : $unsigned(reg431))) && $unsigned(reg444)));
              reg462 <= $unsigned((((~^(reg438 ?
                      wire421 : wire424)) <= reg428[(4'ha):(1'h0)]) ?
                  $unsigned(reg431[(1'h1):(1'h0)]) : (8'h9c)));
            end
          if ((((~&$unsigned((wire422 ? reg433 : reg433))) ?
                  reg439[(4'hb):(2'h3)] : {reg442,
                      $unsigned(((8'hab) >= reg443))}) ?
              (+$unsigned($signed((reg433 ?
                  wire424 : reg433)))) : reg440[(1'h0):(1'h0)]))
            begin
              reg463 <= {$unsigned(reg428), $unsigned($unsigned(reg453))};
              reg464 <= ($signed({((reg440 ?
                      reg428 : wire426) & (reg429 < (7'h40))),
                  $signed(reg440)}) <= (~^($unsigned($signed(reg443)) ?
                  $unsigned((|reg450)) : (!$unsigned((8'hb0))))));
              reg465 <= $signed(reg457[(3'h4):(2'h2)]);
              reg466 <= reg443[(5'h10):(4'h8)];
            end
          else
            begin
              reg463 <= (reg463 < (^~(reg453 ?
                  ((|reg457) ?
                      (reg440 ?
                          wire424 : reg453) : (reg459 & (8'hb7))) : ($signed(reg452) ?
                      reg464 : (reg462 ? reg428 : reg429)))));
              reg464 <= $unsigned((8'hae));
              reg465 <= reg464;
              reg466 <= $unsigned($unsigned($unsigned(wire423[(5'h11):(1'h1)])));
              reg467 <= (+({(^(wire426 ?
                      reg436 : (8'ha5)))} < $signed($unsigned({reg439,
                  reg444}))));
            end
        end
      else
        begin
          reg459 <= $signed(reg467);
          reg460 <= ($signed(($signed($unsigned(reg456)) <= (+wire423[(4'ha):(1'h1)]))) <= (({$signed(reg441)} >= ((reg455 ?
                      reg445 : reg432) ?
                  (8'ha1) : reg464[(1'h1):(1'h1)])) ?
              wire425[(4'ha):(1'h1)] : reg447));
          reg461 <= (reg447 - reg462);
          reg462 <= $signed($unsigned($signed(reg463[(1'h1):(1'h0)])));
        end
    end
  assign wire468 = ($signed($unsigned(reg456)) ?
                       reg445[(2'h3):(2'h2)] : (reg460 ?
                           $signed((reg459 + (wire448 ?
                               (8'haa) : (8'haf)))) : reg463[(1'h1):(1'h0)]));
  always
    @(posedge clk) begin
      if ((+wire448[(1'h1):(1'h0)]))
        begin
          reg469 <= (~|$unsigned((reg447 ?
              $signed((reg428 ? reg443 : reg464)) : ($unsigned(reg465) ?
                  (reg457 >= reg455) : $signed(reg446)))));
          if ($signed((!(reg431 ?
              ({(8'ha6)} * {reg434, reg437}) : ($signed(wire426) ?
                  (reg437 * reg429) : (reg466 ? (8'hb9) : wire448))))))
            begin
              reg470 <= (^~$unsigned(($signed({reg429}) ?
                  reg441[(3'h5):(1'h0)] : $unsigned(((8'hae) && wire422)))));
              reg471 <= ($unsigned($signed((~|reg455))) ?
                  $unsigned(wire425[(3'h6):(2'h3)]) : $unsigned(reg449[(3'h6):(3'h4)]));
              reg472 <= $signed($signed({((+reg462) ?
                      reg451[(1'h1):(1'h0)] : (^reg465)),
                  wire424[(1'h0):(1'h0)]}));
            end
          else
            begin
              reg470 <= $signed(reg443[(1'h1):(1'h1)]);
              reg471 <= $signed(reg437);
              reg472 <= wire424;
              reg473 <= ($signed($unsigned(((reg437 <= reg438) | $unsigned(reg435)))) != $signed($signed((~(-(8'hb3))))));
            end
        end
      else
        begin
          reg469 <= $signed({reg427, reg462});
        end
      reg474 <= (wire468[(1'h0):(1'h0)] <= (reg436[(2'h2):(1'h1)] - ($signed({reg427}) ?
          ((~|wire448) ? (reg455 > reg466) : (~reg456)) : (8'hba))));
      reg475 <= (~^$signed(reg453[(4'h8):(2'h3)]));
      reg476 <= reg463;
      reg477 <= ($unsigned(reg430[(1'h1):(1'h1)]) && $unsigned($unsigned(reg428)));
    end
  assign wire478 = wire422;
  module479 modinst553 (wire552, clk, reg427, reg450, reg431, reg459);
  assign wire554 = $unsigned((((+(reg441 != (8'h9e))) >= reg447) ?
                       (~$unsigned($signed(reg429))) : wire552));
  assign wire555 = $signed((~$signed($signed($unsigned((8'hb1))))));
  assign wire556 = $signed((~|$unsigned({$signed(reg442), wire423})));
  assign wire557 = $signed((^(reg447[(4'h8):(1'h1)] ?
                       ({wire426, reg437} >>> $unsigned(wire555)) : reg467)));
  assign wire558 = (wire468[(3'h4):(1'h0)] ?
                       {(reg441 ?
                               reg429 : $signed((reg435 ? wire422 : (8'ha5)))),
                           (((&reg441) << reg456[(1'h1):(1'h0)]) ?
                               (!wire555) : (((8'ha6) ?
                                   reg456 : reg458) != (wire554 ?
                                   reg444 : reg474)))} : {((8'ha6) <= (|((8'ha8) == reg463)))});
  module559 modinst603 (wire602, clk, wire425, wire558, wire554, reg428);
  always
    @(posedge clk) begin
      if ($unsigned(reg430[(1'h1):(1'h0)]))
        begin
          if ($unsigned((wire558 != ({(wire422 ? reg438 : reg439)} ?
              {(^(8'hb9)), (reg466 ? reg452 : reg446)} : reg439))))
            begin
              reg604 <= (reg441[(2'h2):(1'h1)] <<< $signed((($signed(reg441) ?
                      reg430 : {reg475, wire422}) ?
                  ($signed(reg452) == reg464[(3'h4):(2'h3)]) : wire552[(1'h0):(1'h0)])));
              reg605 <= ($signed($signed(reg473)) ?
                  $signed($unsigned($signed(reg438[(4'he):(3'h6)]))) : $unsigned($signed(reg473)));
              reg606 <= {($unsigned(wire421) & $signed(($signed((7'h42)) || reg470))),
                  $unsigned(($unsigned((~(8'hb5))) ?
                      ((reg429 ?
                          wire552 : reg433) > reg460[(3'h4):(2'h3)]) : ((reg435 | reg469) <<< $signed(wire552))))};
              reg607 <= reg455;
            end
          else
            begin
              reg604 <= reg455;
              reg605 <= reg460;
            end
          reg608 <= ({(7'h42),
              ($unsigned((reg476 * reg430)) == (wire424 ?
                  reg432 : reg465))} != reg427[(1'h1):(1'h1)]);
          reg609 <= $unsigned((^~(reg464[(2'h3):(1'h1)] ?
              (^$unsigned(reg476)) : (((8'ha8) ? reg604 : reg608) > reg465))));
        end
      else
        begin
          reg604 <= $signed($unsigned(reg464[(1'h1):(1'h0)]));
        end
    end
  assign wire610 = $unsigned({$signed($signed({reg604})), (^(~|(!wire425)))});
  always
    @(posedge clk) begin
      reg611 <= (($signed(((wire423 ? wire448 : reg442) < (reg452 ?
                  reg458 : reg428))) ?
              (~|reg460) : reg459[(4'hc):(1'h0)]) ?
          $signed((+reg437[(2'h3):(2'h2)])) : reg435);
    end
  assign wire612 = (^reg606[(4'hd):(2'h2)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module559  (y, clk, wire563, wire562, wire561, wire560);
  output wire [(32'h1af):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire563;
  input wire [(4'he):(1'h0)] wire562;
  input wire signed [(4'hb):(1'h0)] wire561;
  input wire signed [(5'h12):(1'h0)] wire560;
  wire [(4'h9):(1'h0)] wire601;
  wire [(2'h2):(1'h0)] wire600;
  wire [(2'h2):(1'h0)] wire599;
  wire signed [(4'ha):(1'h0)] wire598;
  wire [(4'he):(1'h0)] wire597;
  wire [(4'h9):(1'h0)] wire596;
  wire [(4'ha):(1'h0)] wire595;
  wire [(4'he):(1'h0)] wire594;
  wire [(4'h9):(1'h0)] wire593;
  wire [(4'ha):(1'h0)] wire592;
  reg signed [(2'h3):(1'h0)] reg591 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg590 = (1'h0);
  reg [(5'h13):(1'h0)] reg589 = (1'h0);
  reg [(4'hb):(1'h0)] reg588 = (1'h0);
  reg [(5'h10):(1'h0)] reg587 = (1'h0);
  reg [(3'h6):(1'h0)] reg586 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg585 = (1'h0);
  reg [(2'h3):(1'h0)] reg584 = (1'h0);
  reg [(4'he):(1'h0)] reg583 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg581 = (1'h0);
  reg [(3'h5):(1'h0)] reg580 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg579 = (1'h0);
  reg [(4'hd):(1'h0)] reg578 = (1'h0);
  reg [(5'h15):(1'h0)] reg577 = (1'h0);
  reg [(4'he):(1'h0)] reg576 = (1'h0);
  reg [(4'h8):(1'h0)] reg575 = (1'h0);
  reg [(5'h15):(1'h0)] reg574 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg573 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg572 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire571;
  wire signed [(4'hc):(1'h0)] wire570;
  reg [(2'h3):(1'h0)] reg569 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire568;
  wire [(5'h12):(1'h0)] wire567;
  wire signed [(5'h14):(1'h0)] wire566;
  wire [(5'h15):(1'h0)] wire565;
  wire signed [(5'h10):(1'h0)] wire564;
  assign y = {wire601,
                 wire600,
                 wire599,
                 wire598,
                 wire597,
                 wire596,
                 wire595,
                 wire594,
                 wire593,
                 wire592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 reg579,
                 reg578,
                 reg577,
                 reg576,
                 reg575,
                 reg574,
                 reg573,
                 reg572,
                 wire571,
                 wire570,
                 reg569,
                 wire568,
                 wire567,
                 wire566,
                 wire565,
                 wire564,
                 (1'h0)};
  assign wire564 = ((wire560[(5'h12):(4'hb)] * (($unsigned(wire562) ?
                               wire562 : (wire562 ? wire563 : wire563)) ?
                           wire562 : wire563[(4'h8):(3'h7)])) ?
                       $unsigned((($unsigned(wire563) & wire563[(2'h3):(1'h0)]) ^~ $signed((~&wire560)))) : (wire561 ?
                           (({wire563} ? wire561[(1'h0):(1'h0)] : wire562) ?
                               (((8'hae) ^ wire563) ?
                                   {wire562} : $unsigned(wire563)) : $unsigned((wire560 ?
                                   wire560 : wire561))) : ((~&(wire563 - wire563)) <<< $signed({wire563,
                               (8'ha1)}))));
  assign wire565 = wire564;
  assign wire566 = (-$signed($unsigned({((8'hb5) ? wire565 : wire565),
                       wire563[(1'h0):(1'h0)]})));
  assign wire567 = wire561[(2'h3):(2'h2)];
  assign wire568 = wire563[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg569 <= (wire562[(3'h6):(2'h2)] ?
          wire566 : (wire565 || ($signed(wire566[(1'h1):(1'h0)]) < ((wire565 ?
                  wire563 : wire563) ?
              wire560[(4'he):(4'he)] : $unsigned(wire562)))));
    end
  assign wire570 = {wire560[(5'h11):(4'he)]};
  assign wire571 = $unsigned($signed((((+wire560) <<< $signed((8'hac))) ?
                       wire564[(3'h5):(2'h3)] : wire564[(2'h2):(1'h0)])));
  always
    @(posedge clk) begin
      if ($signed(((8'hbd) ?
          $unsigned($unsigned($signed(wire570))) : {((~wire570) < wire571[(2'h3):(1'h1)]),
              wire567[(4'hb):(3'h6)]})))
        begin
          reg572 <= ((^wire567) | (wire571 ?
              ($unsigned($signed((8'ha5))) ?
                  ($unsigned(wire563) ?
                      wire565 : (wire567 >> wire560)) : ($unsigned(wire564) ~^ wire570[(3'h6):(2'h2)])) : wire568));
          reg573 <= ($signed(wire570[(4'ha):(3'h7)]) < wire567[(4'hc):(4'ha)]);
        end
      else
        begin
          if ((wire571 ? $unsigned({(8'hb7)}) : wire562))
            begin
              reg572 <= wire571[(2'h2):(2'h2)];
              reg573 <= ((wire568[(5'h10):(4'hb)] && (({wire565} ?
                      (wire560 ? wire565 : wire566) : (+wire567)) & wire567)) ?
                  wire561[(3'h6):(3'h6)] : (&((~(wire571 ? wire563 : wire568)) ?
                      (reg572[(3'h5):(1'h0)] ?
                          (~|(8'hb3)) : $unsigned(reg572)) : reg572)));
              reg574 <= ((|{wire570,
                  {(wire570 ? wire570 : reg569),
                      (wire564 - (7'h40))}}) * $unsigned($signed(reg572[(1'h1):(1'h1)])));
              reg575 <= reg573[(3'h5):(3'h4)];
            end
          else
            begin
              reg572 <= (($signed(({reg572,
                      (8'hb5)} >> $signed(reg574))) >> (^{reg569, (8'ha3)})) ?
                  $signed((^wire567)) : $signed($unsigned($signed((reg575 ?
                      wire564 : reg573)))));
              reg573 <= ((wire571 < $signed($unsigned((^wire570)))) ^~ $signed(reg569[(1'h0):(1'h0)]));
              reg574 <= ((+{reg575, (&(8'ha6))}) ?
                  (($unsigned({reg575, wire561}) >= wire563) ?
                      wire560[(2'h3):(2'h3)] : wire567) : wire564[(4'hb):(3'h6)]);
              reg575 <= reg572[(2'h2):(1'h1)];
            end
          reg576 <= (+{(7'h41)});
          reg577 <= wire568[(5'h10):(3'h4)];
          reg578 <= $unsigned(wire564[(1'h0):(1'h0)]);
        end
      if (reg574)
        begin
          reg579 <= $unsigned((+(+(~(wire568 ? (8'hb2) : wire562)))));
          reg580 <= $unsigned(({$unsigned((reg579 ?
                  wire565 : wire564))} && $unsigned({wire568})));
          reg581 <= (8'hb8);
          if (wire564)
            begin
              reg582 <= $unsigned({reg576});
            end
          else
            begin
              reg582 <= (({($signed(reg580) ?
                              wire564[(2'h2):(1'h1)] : $unsigned((8'ha7)))} ?
                      (-$signed($signed(wire561))) : ($signed((!wire567)) | $unsigned((wire570 ?
                          reg580 : reg580)))) ?
                  (|(((-wire571) >>> (!(8'hbb))) ?
                      reg569 : ((reg578 == reg579) << (&wire571)))) : $signed((wire568 ?
                      (reg569 <<< (~&reg578)) : ($unsigned(wire563) ?
                          reg578 : $signed(wire560)))));
              reg583 <= (reg576[(2'h2):(1'h1)] ?
                  reg572 : (wire565 ? (~(-reg582)) : wire562));
            end
        end
      else
        begin
          reg579 <= reg574;
          reg580 <= (($unsigned((&reg569)) ?
                  (wire564[(1'h0):(1'h0)] ?
                      ((wire563 ?
                          wire564 : (8'haa)) ~^ $signed(wire561)) : $signed(reg578)) : reg582) ?
              (7'h44) : ((wire562[(3'h7):(3'h5)] ?
                  (~^$unsigned((8'hb1))) : reg582) & {reg569[(1'h1):(1'h1)]}));
        end
      if (wire561[(3'h6):(2'h2)])
        begin
          reg584 <= $unsigned((reg581 ^~ $signed($signed((-(8'ha7))))));
          reg585 <= (8'haa);
          reg586 <= (((~^($unsigned(wire570) ?
              $signed(wire562) : (8'hbc))) < wire568[(3'h5):(1'h1)]) + (~(($signed(wire568) >= (wire567 <= wire564)) ?
              (|((8'hb3) ? reg576 : wire564)) : $signed($signed(wire571)))));
          reg587 <= wire562;
        end
      else
        begin
          reg584 <= (wire566[(4'hb):(1'h0)] ?
              $unsigned((^$signed((-wire565)))) : reg579[(3'h5):(1'h0)]);
          reg585 <= (!{reg579[(1'h0):(1'h0)],
              ((8'ha9) <<< (wire567[(3'h4):(3'h4)] >> (-reg586)))});
          if ($unsigned($signed((^$signed((reg577 ? (8'hb9) : wire562))))))
            begin
              reg586 <= $signed(reg585[(3'h4):(2'h2)]);
              reg587 <= $signed((reg576[(2'h3):(1'h1)] ?
                  $signed(reg574[(5'h11):(4'hc)]) : (&reg575[(3'h6):(1'h1)])));
            end
          else
            begin
              reg586 <= reg579;
              reg587 <= reg575;
              reg588 <= reg576;
            end
          reg589 <= (~^(reg576 ?
              {(^(reg580 ?
                      wire566 : (8'ha9)))} : ((-{reg583}) > reg584[(2'h2):(2'h2)])));
        end
      reg590 <= $signed(((!reg577[(2'h2):(1'h1)]) ^ $unsigned(reg572[(1'h1):(1'h1)])));
      reg591 <= $signed(((reg588 >> ((-reg573) | wire570[(4'h8):(3'h6)])) ?
          ((^~reg583[(3'h6):(1'h1)]) ^ {wire570[(1'h1):(1'h0)],
              $signed((8'ha2))}) : ($unsigned($signed(reg587)) >= $signed((reg572 ?
              reg579 : reg573)))));
    end
  assign wire592 = wire570;
  assign wire593 = reg573[(3'h4):(1'h1)];
  assign wire594 = (reg588 >= (8'had));
  assign wire595 = ($signed($unsigned($signed($unsigned(reg583)))) ^~ wire566[(1'h1):(1'h0)]);
  assign wire596 = $signed({wire561[(4'ha):(3'h7)],
                       (+(!reg577[(4'h9):(3'h5)]))});
  assign wire597 = {wire567};
  assign wire598 = (~&(reg583[(1'h0):(1'h0)] - (8'ha0)));
  assign wire599 = reg583[(1'h0):(1'h0)];
  assign wire600 = $unsigned(wire597[(2'h3):(2'h3)]);
  assign wire601 = (^$signed((~^(-wire566[(2'h3):(2'h3)]))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module479
#( parameter param550 = ((^~{((!(8'ha9)) ? (!(8'h9f)) : (^(8'ha4)))}) | (((|((8'ha3) == (7'h40))) ^ ((~&(8'hb8)) != (~(8'hb6)))) ? (({(8'had)} ? ((8'ha5) <<< (8'hab)) : ((8'hb6) ? (8'ha4) : (8'ha0))) && ((^~(8'ha3)) > ((8'hba) ? (8'ha8) : (7'h40)))) : (~|((|(8'h9e)) < ((8'h9d) >>> (8'hb0))))))
, parameter param551 = (8'hb0) )
(y, clk, wire483, wire482, wire481, wire480);
  output wire [(32'h2c0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire483;
  input wire [(5'h15):(1'h0)] wire482;
  input wire signed [(5'h10):(1'h0)] wire481;
  input wire [(3'h5):(1'h0)] wire480;
  wire signed [(4'ha):(1'h0)] wire549;
  wire signed [(5'h15):(1'h0)] wire548;
  wire [(5'h13):(1'h0)] wire547;
  wire signed [(3'h5):(1'h0)] wire546;
  wire [(4'hd):(1'h0)] wire545;
  wire [(4'h9):(1'h0)] wire544;
  reg signed [(3'h7):(1'h0)] reg543 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg542 = (1'h0);
  reg [(4'h8):(1'h0)] reg541 = (1'h0);
  wire [(3'h6):(1'h0)] wire540;
  wire signed [(3'h6):(1'h0)] wire539;
  reg [(5'h12):(1'h0)] reg538 = (1'h0);
  reg [(4'ha):(1'h0)] reg537 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg536 = (1'h0);
  reg [(2'h2):(1'h0)] reg535 = (1'h0);
  reg [(3'h5):(1'h0)] reg534 = (1'h0);
  reg [(4'hd):(1'h0)] reg533 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg532 = (1'h0);
  reg [(4'h8):(1'h0)] reg531 = (1'h0);
  reg [(4'hb):(1'h0)] reg530 = (1'h0);
  reg [(2'h3):(1'h0)] reg529 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg528 = (1'h0);
  reg [(3'h6):(1'h0)] reg527 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg526 = (1'h0);
  reg [(4'hf):(1'h0)] reg525 = (1'h0);
  reg [(5'h13):(1'h0)] reg524 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg523 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg522 = (1'h0);
  wire [(3'h4):(1'h0)] wire521;
  wire signed [(3'h5):(1'h0)] wire520;
  reg signed [(4'ha):(1'h0)] reg519 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg518 = (1'h0);
  reg [(4'h8):(1'h0)] reg517 = (1'h0);
  reg [(4'hc):(1'h0)] reg516 = (1'h0);
  reg [(5'h12):(1'h0)] reg515 = (1'h0);
  reg [(5'h10):(1'h0)] reg514 = (1'h0);
  reg [(5'h15):(1'h0)] reg513 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg512 = (1'h0);
  reg signed [(4'he):(1'h0)] reg511 = (1'h0);
  reg [(2'h2):(1'h0)] reg510 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg509 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg508 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg507 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg506 = (1'h0);
  reg [(5'h13):(1'h0)] reg505 = (1'h0);
  reg [(5'h14):(1'h0)] reg504 = (1'h0);
  reg [(4'hc):(1'h0)] reg503 = (1'h0);
  reg [(3'h5):(1'h0)] reg502 = (1'h0);
  reg [(3'h7):(1'h0)] reg501 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg500 = (1'h0);
  reg [(5'h15):(1'h0)] reg499 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg498 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg497 = (1'h0);
  reg [(3'h4):(1'h0)] reg496 = (1'h0);
  reg [(5'h11):(1'h0)] reg495 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg494 = (1'h0);
  reg [(3'h4):(1'h0)] reg493 = (1'h0);
  reg [(4'hd):(1'h0)] reg492 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg491 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg490 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg489 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire488;
  wire signed [(5'h15):(1'h0)] wire487;
  wire [(3'h5):(1'h0)] wire486;
  wire signed [(4'h9):(1'h0)] wire485;
  wire signed [(5'h13):(1'h0)] wire484;
  assign y = {wire549,
                 wire548,
                 wire547,
                 wire546,
                 wire545,
                 wire544,
                 reg543,
                 reg542,
                 reg541,
                 wire540,
                 wire539,
                 reg538,
                 reg537,
                 reg536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 reg522,
                 wire521,
                 wire520,
                 reg519,
                 reg518,
                 reg517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 reg501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 reg491,
                 reg490,
                 reg489,
                 wire488,
                 wire487,
                 wire486,
                 wire485,
                 wire484,
                 (1'h0)};
  assign wire484 = {wire480[(2'h3):(1'h0)]};
  assign wire485 = {wire484};
  assign wire486 = $signed(wire484);
  assign wire487 = (~^$unsigned((wire481[(3'h7):(3'h7)] ?
                       wire483[(1'h0):(1'h0)] : (wire485[(3'h6):(3'h4)] ?
                           {(8'ha3), wire481} : {wire480}))));
  assign wire488 = ((($signed($unsigned(wire481)) ?
                           (^~(wire486 - wire485)) : $signed($unsigned(wire484))) ?
                       $unsigned(wire485[(3'h4):(1'h0)]) : (wire486 << (~^$signed(wire480)))) && wire484[(5'h10):(4'hb)]);
  always
    @(posedge clk) begin
      if ($unsigned(wire484))
        begin
          reg489 <= ({$unsigned($unsigned((+wire485)))} ?
              wire480 : wire488[(2'h2):(2'h2)]);
          if (wire481[(4'hd):(4'ha)])
            begin
              reg490 <= wire480;
              reg491 <= $unsigned((+({$unsigned(wire482),
                      reg489[(2'h2):(2'h2)]} ?
                  ((reg489 ^~ reg490) ?
                      $unsigned(wire482) : (&wire487)) : $signed((wire486 <<< wire481)))));
              reg492 <= ($unsigned($unsigned(((&wire488) >>> (8'hab)))) && wire486);
            end
          else
            begin
              reg490 <= ($unsigned((wire481[(2'h3):(2'h3)] - (8'hba))) && (!wire488));
              reg491 <= {(wire487 ?
                      $unsigned((wire482[(3'h7):(1'h1)] & {wire485,
                          wire480})) : $signed(((wire482 ?
                          reg492 : (8'hb4)) <= (wire486 & (8'hbd)))))};
              reg492 <= $unsigned((~&{wire487[(4'h9):(2'h3)]}));
              reg493 <= $signed(($unsigned((wire488[(3'h4):(3'h4)] | wire484)) ?
                  reg489[(2'h2):(2'h2)] : $unsigned($signed((wire481 == wire483)))));
            end
          reg494 <= ($unsigned((wire488[(1'h0):(1'h0)] ^~ (!wire487[(3'h6):(3'h5)]))) ?
              wire481 : (8'ha0));
          if (((({$signed(wire485), {wire487, wire480}} ?
                      $signed((wire486 + reg494)) : wire484) ?
                  (+(reg489[(3'h4):(3'h4)] != (~&(7'h43)))) : (^{$signed(wire483)})) ?
              $signed(({(-wire483)} + $unsigned($unsigned(wire480)))) : (&reg490[(2'h2):(1'h1)])))
            begin
              reg495 <= reg490;
              reg496 <= ($unsigned((((+reg493) ~^ (reg490 & (8'ha8))) || $signed((~&wire487)))) ^~ ((wire485[(4'h9):(3'h5)] ?
                      ((wire488 == wire488) ?
                          (wire482 ?
                              wire483 : wire484) : wire485[(2'h2):(2'h2)]) : reg490) ?
                  ((~^wire482) ?
                      $unsigned((&(8'ha6))) : (&$signed(reg494))) : (~|$unsigned((&wire484)))));
              reg497 <= wire481;
              reg498 <= (wire483 ?
                  (wire486 >> $unsigned($signed({(8'ha7)}))) : (wire480 | ((wire480 ?
                      (wire484 ?
                          (8'h9c) : reg493) : (8'hbb)) > $unsigned(((8'ha8) < reg490)))));
            end
          else
            begin
              reg495 <= reg494;
            end
        end
      else
        begin
          reg489 <= $signed($unsigned((~&((^~(8'h9f)) ?
              $signed(reg493) : (-(8'hbb))))));
        end
      reg499 <= reg498;
      reg500 <= $signed($unsigned(reg499));
      reg501 <= ($signed((+(&wire488))) >>> ($signed($signed(wire482)) ?
          (~($unsigned(wire480) ~^ wire484)) : (~^{wire482[(4'hc):(3'h4)]})));
      if ((|(reg499 ?
          wire481 : $signed($unsigned((reg498 ? reg491 : reg497))))))
        begin
          if (reg494)
            begin
              reg502 <= (wire486[(2'h3):(1'h1)] ?
                  reg496[(3'h4):(1'h0)] : {reg489, (reg499 << reg492)});
            end
          else
            begin
              reg502 <= reg491;
              reg503 <= $unsigned($signed((wire483 * {$unsigned(reg493),
                  $unsigned(wire487)})));
              reg504 <= (~^$signed(wire487[(5'h15):(4'hb)]));
            end
          if ($unsigned(wire486))
            begin
              reg505 <= $unsigned(($signed((~((8'ha3) <= wire486))) ?
                  ($signed((8'h9f)) ?
                      reg493[(3'h4):(2'h2)] : (reg492[(3'h7):(3'h6)] + reg499[(4'hc):(1'h0)])) : ($unsigned($signed(reg496)) ?
                      $unsigned($unsigned((8'hab))) : $signed((~(8'ha4))))));
              reg506 <= ($signed(wire480) ? $signed((&reg497)) : wire486);
              reg507 <= reg500;
            end
          else
            begin
              reg505 <= (((8'hb2) ?
                      (($unsigned(wire482) & $signed(wire488)) <<< (((7'h43) ?
                          wire488 : wire480) ^~ wire483)) : wire487) ?
                  (8'ha2) : (((~$signed((7'h42))) ?
                          $signed($signed(wire483)) : reg491) ?
                      $unsigned((8'hb1)) : (reg499 * reg497[(1'h1):(1'h0)])));
              reg506 <= (~((~^reg502[(1'h0):(1'h0)]) || (^~{wire485[(1'h0):(1'h0)],
                  reg497[(2'h3):(1'h1)]})));
              reg507 <= reg503;
              reg508 <= reg490;
              reg509 <= ((((-reg493[(3'h4):(2'h3)]) | {(8'hb8),
                  {wire485, wire482}}) ~^ ($signed((reg499 ?
                      (8'ha4) : wire487)) ?
                  (|reg499) : wire488)) ^ ($signed({reg504,
                      $unsigned(reg496)}) ?
                  reg507[(4'he):(2'h2)] : (^reg507[(4'he):(3'h6)])));
            end
          if ($signed(wire483))
            begin
              reg510 <= ({reg493, reg498[(3'h5):(3'h4)]} ?
                  $signed(wire481) : ({reg509[(4'hb):(3'h7)]} ?
                      reg501[(2'h3):(2'h3)] : $signed($signed($unsigned(reg495)))));
              reg511 <= $unsigned(({$unsigned($signed(reg510))} * $unsigned({reg501})));
              reg512 <= (((~&reg497) ?
                  reg504 : (wire487 <= (^$signed(reg503)))) != {(((7'h43) ?
                      $signed(reg510) : $unsigned(reg504)) && {(reg508 ?
                          reg503 : reg489)})});
              reg513 <= reg496;
              reg514 <= $unsigned((!({reg506[(1'h0):(1'h0)]} ~^ ($unsigned(wire482) ?
                  reg491 : (wire486 ? wire483 : reg506)))));
            end
          else
            begin
              reg510 <= (reg512 ?
                  (wire487 ?
                      reg506 : {reg512,
                          reg514[(2'h2):(1'h1)]}) : $signed(((reg493[(1'h1):(1'h1)] ?
                          (reg489 || reg512) : wire480) ?
                      $signed((^~reg502)) : reg500)));
              reg511 <= (((^~(~|(reg505 <<< reg489))) >= (($unsigned(reg509) ?
                          reg502[(2'h3):(2'h3)] : (reg503 | (8'ha5))) ?
                      $unsigned($signed(wire485)) : reg492[(4'h9):(3'h4)])) ?
                  $signed($unsigned($signed((~^reg493)))) : reg504[(2'h3):(1'h1)]);
            end
          if ((~|({$unsigned((reg497 ? reg508 : reg513))} ?
              {($signed(wire484) ? $unsigned(reg490) : $signed(reg502)),
                  reg499} : ((&$signed(reg513)) ?
                  $signed((wire482 ?
                      reg506 : wire481)) : {$unsigned((8'hb4))}))))
            begin
              reg515 <= reg492;
              reg516 <= $unsigned(($signed($signed($unsigned(reg510))) - $unsigned({(+reg493)})));
              reg517 <= reg509[(4'hf):(2'h2)];
              reg518 <= $signed({((!reg514) * reg502), (~|$unsigned(reg505))});
            end
          else
            begin
              reg515 <= (reg512[(4'ha):(3'h5)] - (((8'ha8) ?
                      $unsigned($signed((8'ha1))) : reg499) ?
                  reg501[(2'h2):(1'h1)] : reg500));
              reg516 <= reg490;
              reg517 <= (+wire480);
              reg518 <= $signed(reg516);
            end
          reg519 <= reg515;
        end
      else
        begin
          if ((~^(8'hab)))
            begin
              reg502 <= wire487[(4'hb):(4'h9)];
              reg503 <= $unsigned(reg511[(4'he):(1'h0)]);
            end
          else
            begin
              reg502 <= (((~^(reg495 ?
                      {reg517, wire483} : reg489[(2'h2):(2'h2)])) & reg502) ?
                  $signed(({reg494[(4'hc):(1'h0)]} ?
                      $signed(wire483[(3'h5):(2'h2)]) : reg498[(3'h6):(2'h3)])) : ($signed(reg508[(1'h0):(1'h0)]) ?
                      (reg499 ?
                          $signed(reg506[(1'h1):(1'h1)]) : $unsigned(reg506)) : wire482[(5'h15):(4'hc)]));
              reg503 <= reg506;
              reg504 <= reg506[(1'h0):(1'h0)];
            end
        end
    end
  assign wire520 = $signed(((reg499[(3'h7):(1'h0)] ?
                       wire481[(4'ha):(1'h0)] : $unsigned($signed(reg517))) && ((^~$signed((8'ha7))) ?
                       ($signed(wire482) <= reg514) : ((+reg509) ?
                           $signed(reg491) : (8'hb6)))));
  assign wire521 = {{((wire480[(3'h4):(3'h4)] ?
                                   $unsigned(reg513) : $signed(wire482)) ?
                               ((-wire480) ?
                                   ((7'h44) + reg504) : (~|(8'haa))) : (~|(reg519 || reg507))),
                           (8'ha3)},
                       ($unsigned(reg499) >= $unsigned((~&reg518)))};
  always
    @(posedge clk) begin
      if ($unsigned($unsigned((reg490[(4'ha):(4'h8)] | wire483[(3'h4):(3'h4)]))))
        begin
          reg522 <= $signed($signed((8'hba)));
          if ((({wire482,
                      ((reg491 ? wire488 : reg522) ?
                          $signed(reg496) : reg522[(2'h3):(1'h0)])} ?
                  (+(reg502 ? {reg511, wire481} : (~&wire521))) : reg501) ?
              (&$unsigned($unsigned((~|wire487)))) : reg502[(2'h3):(1'h0)]))
            begin
              reg523 <= $unsigned($signed($signed($signed((reg490 ?
                  reg507 : wire488)))));
              reg524 <= (wire480 <<< ({((-wire482) ~^ (~reg501)),
                  {{(8'ha0), reg507},
                      (reg513 << (8'ha2))}} <<< (((reg506 || (8'ha4)) == $unsigned(reg506)) != ((-(8'haa)) ?
                  (reg514 ? reg493 : wire482) : $unsigned(reg490)))));
            end
          else
            begin
              reg523 <= wire488;
              reg524 <= reg518[(4'h9):(3'h6)];
              reg525 <= ($signed($signed(reg498[(4'h8):(3'h4)])) ?
                  (7'h40) : $signed({(reg498[(1'h0):(1'h0)] ?
                          $unsigned(wire480) : (reg499 ? reg498 : reg518))}));
            end
          reg526 <= (((((|reg489) ? reg503 : wire486[(1'h0):(1'h0)]) ^ (reg505 ?
                  (~^reg524) : (reg494 ?
                      reg515 : reg504))) < $signed(wire483[(3'h4):(1'h1)])) ?
              ($unsigned($signed($unsigned(reg508))) ?
                  reg525 : (!($unsigned(reg502) | reg523[(1'h0):(1'h0)]))) : $signed(((~$unsigned(reg523)) * reg498)));
        end
      else
        begin
          reg522 <= reg490[(2'h3):(2'h3)];
          if ((!(8'hbf)))
            begin
              reg523 <= $unsigned(wire482);
              reg524 <= $signed($unsigned(($unsigned($signed(reg497)) ?
                  {reg507, reg525[(4'ha):(4'ha)]} : (7'h42))));
              reg525 <= $unsigned({wire480[(2'h2):(2'h2)],
                  (+(reg513 ? (wire480 ~^ wire483) : $unsigned(wire487)))});
            end
          else
            begin
              reg523 <= (!reg497);
              reg524 <= ($signed(reg505[(4'h9):(2'h3)]) ~^ $signed({($signed(wire520) ?
                      (reg506 ? reg496 : reg526) : wire482),
                  (~|wire487[(5'h13):(5'h11)])}));
            end
          reg526 <= (&(-reg507));
          if (((7'h44) << {((~(&reg508)) << {reg489,
                  (reg494 ? reg503 : reg501)})}))
            begin
              reg527 <= reg498[(4'hd):(4'hb)];
              reg528 <= $signed({$signed({{reg514, reg517}}),
                  $unsigned($unsigned($signed((8'hb1))))});
            end
          else
            begin
              reg527 <= $unsigned(reg499);
              reg528 <= $unsigned($signed((^~$signed($unsigned(reg493)))));
              reg529 <= ((|(&$unsigned((8'ha4)))) >> (8'ha8));
              reg530 <= {wire485};
            end
        end
      reg531 <= reg508[(1'h0):(1'h0)];
      reg532 <= $signed((reg523 && $unsigned({(~^wire520),
          (reg500 ^ reg514)})));
      if (reg501)
        begin
          reg533 <= reg494;
          reg534 <= (&wire483);
        end
      else
        begin
          reg533 <= wire484;
          reg534 <= $unsigned((reg505[(4'h8):(3'h6)] > reg507));
          if ((8'ha6))
            begin
              reg535 <= {$signed($signed($signed((-(7'h43)))))};
              reg536 <= ($signed((!(reg517[(3'h5):(1'h1)] ?
                  (reg535 < reg528) : (reg529 && wire485)))) > (~&reg528));
            end
          else
            begin
              reg535 <= $unsigned(reg523);
              reg536 <= reg490;
              reg537 <= $unsigned($signed((~&(reg531[(2'h3):(1'h1)] ?
                  $unsigned(reg493) : (reg490 ? wire482 : reg496)))));
            end
        end
      reg538 <= $unsigned(reg515[(4'hd):(4'hd)]);
    end
  assign wire539 = {$unsigned(reg538[(5'h11):(2'h3)])};
  assign wire540 = $signed(($unsigned(reg529) || {$signed($signed(reg518))}));
  always
    @(posedge clk) begin
      reg541 <= reg492;
      reg542 <= (($unsigned(((!reg529) >>> $unsigned(reg541))) != $signed((+$signed(wire484)))) ?
          reg497[(1'h0):(1'h0)] : reg512[(5'h13):(4'ha)]);
      reg543 <= reg542;
    end
  assign wire544 = $signed((reg523[(3'h5):(2'h2)] <= (wire481[(3'h7):(2'h3)] ?
                       {reg514[(3'h6):(3'h4)]} : $unsigned(wire481[(2'h2):(1'h0)]))));
  assign wire545 = {(8'hb1)};
  assign wire546 = $signed({$unsigned($signed($unsigned((8'hb3)))),
                       reg508[(2'h2):(2'h2)]});
  assign wire547 = $signed($unsigned(((8'haa) ?
                       $signed($unsigned(wire486)) : $signed((reg501 ?
                           (8'haa) : reg531)))));
  assign wire548 = {reg489};
  assign wire549 = {$signed($unsigned($unsigned((8'hb2))))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module663
#( parameter param672 = {{((((8'hb0) || (8'haf)) >> {(8'hb2)}) & (((8'ha5) - (8'had)) ? ((8'h9f) || (8'ha6)) : (8'hbc)))}}
, parameter param673 = (^~(((param672 ? (param672 ? param672 : param672) : ((8'h9e) - param672)) ? {(param672 ? param672 : param672), (param672 ? param672 : param672)} : param672) > param672)) )
(y, clk, wire667, wire666, wire665, wire664);
  output wire [(32'h33):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire667;
  input wire [(4'hb):(1'h0)] wire666;
  input wire signed [(2'h2):(1'h0)] wire665;
  input wire [(5'h13):(1'h0)] wire664;
  wire [(2'h2):(1'h0)] wire671;
  wire signed [(4'hf):(1'h0)] wire670;
  wire signed [(5'h11):(1'h0)] wire669;
  wire signed [(5'h10):(1'h0)] wire668;
  assign y = {wire671, wire670, wire669, wire668, (1'h0)};
  assign wire668 = (wire664[(4'ha):(4'ha)] && ((8'hab) ?
                       ($signed($unsigned((8'ha2))) >> {wire667}) : wire667[(3'h7):(3'h7)]));
  assign wire669 = (|($signed((8'hb5)) | (($unsigned(wire665) & $unsigned(wire667)) ^ wire667)));
  assign wire670 = $signed(wire669[(5'h11):(4'hb)]);
  assign wire671 = wire665;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module871  (y, clk, wire875, wire874, wire873, wire872);
  output wire [(32'h41):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire875;
  input wire signed [(3'h6):(1'h0)] wire874;
  input wire signed [(4'hc):(1'h0)] wire873;
  input wire signed [(5'h10):(1'h0)] wire872;
  wire signed [(4'hf):(1'h0)] wire879;
  wire signed [(5'h15):(1'h0)] wire878;
  wire signed [(5'h11):(1'h0)] wire877;
  wire signed [(4'hb):(1'h0)] wire876;
  assign y = {wire879, wire878, wire877, wire876, (1'h0)};
  assign wire876 = (!$unsigned((&{wire873, wire872[(4'hd):(1'h0)]})));
  assign wire877 = wire872;
  assign wire878 = $unsigned(((7'h42) ?
                       wire873[(2'h3):(2'h2)] : ((+(wire876 << wire875)) ?
                           (8'ha8) : $signed($unsigned(wire877)))));
  assign wire879 = wire874;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module701
#( parameter param866 = {({(((8'haa) ? (8'hae) : (8'hab)) ? (~^(8'hb9)) : (~(8'ha1)))} <= (8'hb4))}
, parameter param867 = (|(~&(({param866} > (param866 <= param866)) >= (^~(&param866))))) )
(y, clk, wire705, wire704, wire703, wire702);
  output wire [(32'hf5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire705;
  input wire signed [(5'h13):(1'h0)] wire704;
  input wire signed [(5'h14):(1'h0)] wire703;
  input wire signed [(5'h15):(1'h0)] wire702;
  wire [(4'hb):(1'h0)] wire865;
  wire [(4'h9):(1'h0)] wire864;
  wire signed [(5'h10):(1'h0)] wire863;
  wire signed [(2'h3):(1'h0)] wire862;
  wire signed [(3'h5):(1'h0)] wire861;
  wire [(3'h4):(1'h0)] wire860;
  wire [(4'h8):(1'h0)] wire858;
  wire [(4'he):(1'h0)] wire833;
  wire [(4'h9):(1'h0)] wire832;
  reg signed [(4'hc):(1'h0)] reg831 = (1'h0);
  reg [(3'h6):(1'h0)] reg830 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg829 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg828 = (1'h0);
  reg [(3'h4):(1'h0)] reg827 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg826 = (1'h0);
  wire [(5'h15):(1'h0)] wire825;
  wire signed [(5'h11):(1'h0)] wire824;
  wire [(3'h5):(1'h0)] wire823;
  wire signed [(4'hd):(1'h0)] wire787;
  wire signed [(5'h14):(1'h0)] wire749;
  reg signed [(5'h13):(1'h0)] reg707 = (1'h0);
  wire [(4'hd):(1'h0)] wire706;
  wire signed [(4'hc):(1'h0)] wire821;
  assign y = {wire865,
                 wire864,
                 wire863,
                 wire862,
                 wire861,
                 wire860,
                 wire858,
                 wire833,
                 wire832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 reg827,
                 reg826,
                 wire825,
                 wire824,
                 wire823,
                 wire787,
                 wire749,
                 reg707,
                 wire706,
                 wire821,
                 (1'h0)};
  assign wire706 = wire703[(3'h7):(3'h6)];
  always
    @(posedge clk) begin
      reg707 <= (wire702[(1'h0):(1'h0)] < {(^~wire703[(4'hc):(4'ha)])});
    end
  module708 modinst750 (.clk(clk), .wire712(wire706), .y(wire749), .wire709(wire702), .wire711(wire704), .wire710(reg707));
  module751 modinst788 (wire787, clk, wire706, wire702, wire704, wire749, wire705);
  module789 modinst822 (.wire793(wire704), .y(wire821), .wire790(wire706), .wire792(wire705), .wire791(reg707), .clk(clk), .wire794(wire787));
  assign wire823 = wire703;
  assign wire824 = (8'hbf);
  assign wire825 = wire705;
  always
    @(posedge clk) begin
      if ($signed((({(&wire705)} ^ wire706) ?
          (-$signed({wire706, wire705})) : (&(wire824 > (~&wire825))))))
        begin
          reg826 <= $signed({(-$unsigned(wire704[(1'h1):(1'h0)]))});
        end
      else
        begin
          reg826 <= $unsigned({(($unsigned(wire787) || wire704[(4'hd):(4'h9)]) <= ($signed((8'ha6)) ?
                  (wire703 ? wire706 : wire703) : wire706)),
              ($signed($unsigned((7'h42))) >> {(wire706 ?
                      (8'hbf) : wire703)})});
          if (wire706[(3'h6):(3'h6)])
            begin
              reg827 <= reg826;
            end
          else
            begin
              reg827 <= wire702;
              reg828 <= (&((wire821 < (~|(~|wire821))) ?
                  $signed($signed((wire702 ?
                      wire703 : (8'hbd)))) : (($unsigned(wire821) * (-wire703)) << wire825[(3'h6):(3'h5)])));
              reg829 <= (~$unsigned(wire825[(4'he):(4'ha)]));
              reg830 <= ((wire825[(5'h14):(1'h1)] ?
                  $unsigned((~&((8'ha0) >> reg829))) : (wire821[(1'h1):(1'h0)] ?
                      $unsigned((wire705 != reg829)) : (+wire787[(3'h6):(3'h6)]))) ^ wire702);
              reg831 <= (~(8'hb1));
            end
        end
    end
  assign wire832 = (~^wire704);
  assign wire833 = wire832;
  module834 modinst859 (wire858, clk, wire703, wire702, reg830, wire706);
  assign wire860 = wire749;
  assign wire861 = $unsigned(((-(~^(8'ha0))) ?
                       $signed((~^(^~wire702))) : (wire860 & $signed((reg830 ?
                           reg830 : reg831)))));
  assign wire862 = wire825;
  assign wire863 = (wire787[(4'h9):(1'h0)] ?
                       wire833 : {(|{$signed((8'h9e)), $signed(reg826)})});
  assign wire864 = wire705;
  assign wire865 = $unsigned(wire824);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module834
#( parameter param856 = (-({(-(^(8'hae)))} >> (({(8'h9e), (8'hac)} ? ((8'h9f) - (8'ha4)) : ((8'ha1) ? (8'hbd) : (8'ha5))) ? (((7'h41) ? (7'h42) : (8'hb9)) ~^ ((8'ha5) != (8'hb5))) : (!(8'hb4)))))
, parameter param857 = param856 )
(y, clk, wire838, wire837, wire836, wire835);
  output wire [(32'hc8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire838;
  input wire [(4'h9):(1'h0)] wire837;
  input wire signed [(3'h6):(1'h0)] wire836;
  input wire [(2'h2):(1'h0)] wire835;
  wire signed [(5'h15):(1'h0)] wire855;
  wire [(3'h4):(1'h0)] wire854;
  wire signed [(4'hc):(1'h0)] wire853;
  wire [(4'ha):(1'h0)] wire852;
  wire signed [(3'h7):(1'h0)] wire851;
  reg [(2'h2):(1'h0)] reg850 = (1'h0);
  reg [(5'h12):(1'h0)] reg849 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire848;
  wire [(4'hc):(1'h0)] wire847;
  wire [(2'h3):(1'h0)] wire846;
  wire [(4'hb):(1'h0)] wire845;
  wire signed [(4'he):(1'h0)] wire844;
  wire [(5'h15):(1'h0)] wire843;
  wire [(4'hb):(1'h0)] wire842;
  reg signed [(5'h14):(1'h0)] reg841 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg840 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire839;
  assign y = {wire855,
                 wire854,
                 wire853,
                 wire852,
                 wire851,
                 reg850,
                 reg849,
                 wire848,
                 wire847,
                 wire846,
                 wire845,
                 wire844,
                 wire843,
                 wire842,
                 reg841,
                 reg840,
                 wire839,
                 (1'h0)};
  assign wire839 = $signed({(((+(8'ha7)) ? {wire836, wire837} : (~^wire836)) ?
                           wire838[(4'h8):(1'h0)] : ((~wire837) ?
                               $signed(wire838) : $signed(wire838))),
                       wire836[(2'h2):(1'h1)]});
  always
    @(posedge clk) begin
      reg840 <= (wire836[(2'h3):(1'h1)] || (!wire835[(1'h1):(1'h0)]));
      reg841 <= $signed({((-((8'hbb) == wire837)) ?
              $unsigned(wire837) : ($signed((8'hb3)) ?
                  $unsigned(wire837) : (&wire838)))});
    end
  assign wire842 = $unsigned({$signed($unsigned(((8'ha5) & wire839))),
                       (reg840 ?
                           ((wire836 ?
                               wire836 : wire837) - {wire837}) : (~wire837[(3'h7):(3'h6)]))});
  assign wire843 = $unsigned(wire836);
  assign wire844 = ($signed(reg840) & ($unsigned(wire836) ?
                       ($signed(wire838) >> wire835) : ((8'hba) ?
                           $signed($signed(wire835)) : (((8'ha0) + wire843) ~^ wire839))));
  assign wire845 = ($unsigned($unsigned($unsigned($signed(wire836)))) | {(-(~^$signed(wire835))),
                       wire836[(2'h3):(2'h2)]});
  assign wire846 = wire844;
  assign wire847 = wire844[(3'h7):(3'h4)];
  assign wire848 = wire847[(4'ha):(2'h2)];
  always
    @(posedge clk) begin
      reg849 <= (^(~^($unsigned((wire837 ?
          wire838 : wire837)) ~^ wire844[(3'h4):(1'h1)])));
      reg850 <= (wire843 > $unsigned(($unsigned((+wire845)) ?
          wire847[(4'hc):(2'h3)] : reg841)));
    end
  assign wire851 = $signed(($signed($unsigned($unsigned((8'hb2)))) ?
                       wire843[(3'h7):(3'h7)] : (|(&(wire845 & wire847)))));
  assign wire852 = wire837[(1'h1):(1'h1)];
  assign wire853 = wire847;
  assign wire854 = (+$signed((wire847[(3'h6):(3'h4)] >>> {wire839[(1'h0):(1'h0)]})));
  assign wire855 = $signed(((!((-wire853) ?
                       (wire846 ~^ wire845) : wire839)) == $signed((8'ha5))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module789
#( parameter param819 = ((((((8'hb7) ? (8'ha3) : (8'hbf)) ? (8'haa) : {(8'h9d), (7'h43)}) ? (((8'ha7) ^~ (8'hb3)) ^ (&(8'hae))) : (((8'hb8) ? (8'h9d) : (8'hbc)) ~^ {(8'hb1)})) ? ((((8'h9d) ? (8'ha6) : (8'ha3)) ? ((8'ha8) * (8'ha3)) : ((8'h9d) ? (8'ha3) : (8'ha1))) ? (((8'hba) <<< (8'ha2)) ^ ((8'h9c) != (8'hac))) : (~|(~|(8'ha4)))) : (((^~(8'ha4)) ? ((8'hab) ? (8'hb0) : (8'hb2)) : ((7'h44) ? (8'hab) : (8'ha2))) ? {(-(7'h43)), (&(8'h9d))} : (|(~^(8'hbb))))) ? (((-(~(8'hb4))) ? (((8'ha5) ? (8'ha5) : (8'ha3)) << (~(8'hba))) : {{(8'hba), (8'h9f)}}) ? (8'hb1) : ((((7'h41) ? (8'had) : (8'hb7)) || {(8'hb7), (8'hae)}) ^ (!(-(8'hb3))))) : ({((^(8'hab)) * (|(8'hb2)))} ? (-((+(8'ha6)) ? {(8'hbe), (8'hb9)} : ((8'hb8) + (8'h9e)))) : (~(((8'hb2) ? (8'hb3) : (8'ha2)) <= (+(8'ha5))))))
, parameter param820 = (!(param819 + param819)) )
(y, clk, wire794, wire793, wire792, wire791, wire790);
  output wire [(32'h113):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire794;
  input wire signed [(4'hd):(1'h0)] wire793;
  input wire [(2'h2):(1'h0)] wire792;
  input wire [(5'h13):(1'h0)] wire791;
  input wire signed [(3'h4):(1'h0)] wire790;
  wire [(4'hc):(1'h0)] wire818;
  wire [(5'h13):(1'h0)] wire817;
  wire [(4'he):(1'h0)] wire816;
  wire [(4'he):(1'h0)] wire815;
  wire signed [(3'h7):(1'h0)] wire814;
  wire [(4'h9):(1'h0)] wire813;
  reg [(5'h10):(1'h0)] reg812 = (1'h0);
  reg [(4'hc):(1'h0)] reg811 = (1'h0);
  reg [(5'h11):(1'h0)] reg810 = (1'h0);
  wire signed [(4'he):(1'h0)] wire809;
  reg [(4'hc):(1'h0)] reg808 = (1'h0);
  reg [(4'h9):(1'h0)] reg807 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg806 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg805 = (1'h0);
  reg [(4'hd):(1'h0)] reg804 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg803 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg802 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg801 = (1'h0);
  reg [(4'hd):(1'h0)] reg800 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg799 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg798 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire797;
  wire signed [(3'h7):(1'h0)] wire796;
  reg signed [(4'ha):(1'h0)] reg795 = (1'h0);
  assign y = {wire818,
                 wire817,
                 wire816,
                 wire815,
                 wire814,
                 wire813,
                 reg812,
                 reg811,
                 reg810,
                 wire809,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg802,
                 reg801,
                 reg800,
                 reg799,
                 reg798,
                 wire797,
                 wire796,
                 reg795,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg795 <= (^~(($unsigned({wire791,
          wire791}) == (~|wire790[(2'h3):(1'h0)])) | wire791));
    end
  assign wire796 = $unsigned($signed({$unsigned($signed(wire792)), (8'hae)}));
  assign wire797 = {(wire790 ? wire794[(1'h1):(1'h0)] : $unsigned(wire790))};
  always
    @(posedge clk) begin
      reg798 <= (wire794[(2'h3):(1'h1)] ?
          $unsigned(wire790) : {{$unsigned((8'hbc)),
                  ((wire793 ? (8'ha7) : wire794) | reg795)},
              ($signed(wire793[(1'h0):(1'h0)]) ?
                  (!{(7'h44)}) : wire790[(1'h0):(1'h0)])});
      reg799 <= $signed(reg798[(3'h5):(1'h1)]);
      if ((~|$signed(wire796)))
        begin
          reg800 <= {$signed((8'hb7)), wire793[(4'hc):(4'h9)]};
          reg801 <= $signed(reg795[(2'h2):(2'h2)]);
        end
      else
        begin
          reg800 <= ((8'ha0) ?
              $unsigned($unsigned($unsigned($unsigned(wire797)))) : (!$unsigned(($signed(reg801) != (reg798 ?
                  reg795 : reg799)))));
          if (wire790)
            begin
              reg801 <= (7'h40);
            end
          else
            begin
              reg801 <= ((^~(^~wire793[(3'h5):(1'h1)])) ?
                  {wire792} : $unsigned({($unsigned((8'hae)) ?
                          reg798 : (wire796 ~^ wire790)),
                      $unsigned((reg800 != reg798))}));
              reg802 <= wire791[(4'hb):(4'h8)];
              reg803 <= (-$unsigned((~^wire797)));
              reg804 <= reg800[(4'h8):(2'h3)];
            end
          reg805 <= (((reg798 ?
                  (&$signed(wire790)) : ((|wire793) ?
                      $unsigned(reg801) : (wire794 ^~ wire791))) - ($signed($signed((8'hbf))) & ($signed(reg801) >= (wire793 ?
                  reg801 : wire790)))) ?
              (~($unsigned($unsigned(reg804)) || $unsigned((reg800 ?
                  (8'ha5) : (7'h43))))) : ($unsigned(reg800) > (&$unsigned((reg795 > wire794)))));
          reg806 <= $unsigned((~&(~&((!wire792) <= {reg803, wire797}))));
          reg807 <= reg806[(1'h1):(1'h0)];
        end
      reg808 <= reg799;
    end
  assign wire809 = wire793[(4'hb):(2'h2)];
  always
    @(posedge clk) begin
      reg810 <= $signed($signed(wire797));
      reg811 <= wire809[(4'h9):(1'h0)];
      reg812 <= $signed((8'hb7));
    end
  assign wire813 = $signed({reg805});
  assign wire814 = ($signed($signed((wire792 ?
                           wire793[(4'hd):(4'h9)] : (-reg799)))) ?
                       $signed($signed($unsigned(reg803[(2'h2):(1'h1)]))) : (~&$unsigned(reg799[(1'h0):(1'h0)])));
  assign wire815 = $signed(wire790[(1'h1):(1'h0)]);
  assign wire816 = (reg799 ?
                       {(reg810[(3'h4):(2'h2)] + $signed((^(8'ha4))))} : wire813[(1'h0):(1'h0)]);
  assign wire817 = wire792[(1'h1):(1'h1)];
  assign wire818 = wire797[(2'h2):(2'h2)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module751  (y, clk, wire756, wire755, wire754, wire753, wire752);
  output wire [(32'h166):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire756;
  input wire [(4'h8):(1'h0)] wire755;
  input wire signed [(5'h11):(1'h0)] wire754;
  input wire signed [(5'h13):(1'h0)] wire753;
  input wire signed [(5'h11):(1'h0)] wire752;
  reg [(5'h14):(1'h0)] reg786 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg785 = (1'h0);
  reg [(4'hc):(1'h0)] reg784 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg783 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg782 = (1'h0);
  reg [(4'hb):(1'h0)] reg781 = (1'h0);
  reg [(5'h14):(1'h0)] reg780 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg779 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg778 = (1'h0);
  reg [(4'h9):(1'h0)] reg777 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg776 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg775 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg774 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg773 = (1'h0);
  reg [(5'h14):(1'h0)] reg772 = (1'h0);
  reg [(4'hd):(1'h0)] reg771 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg770 = (1'h0);
  reg [(5'h12):(1'h0)] reg769 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg768 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire767;
  wire [(4'hd):(1'h0)] wire766;
  wire [(4'hc):(1'h0)] wire765;
  wire signed [(5'h15):(1'h0)] wire764;
  wire signed [(2'h2):(1'h0)] wire763;
  wire [(4'hf):(1'h0)] wire762;
  wire signed [(5'h15):(1'h0)] wire761;
  wire signed [(4'h9):(1'h0)] wire760;
  wire signed [(2'h2):(1'h0)] wire759;
  wire signed [(4'h9):(1'h0)] wire758;
  wire [(4'hc):(1'h0)] wire757;
  assign y = {reg786,
                 reg785,
                 reg784,
                 reg783,
                 reg782,
                 reg781,
                 reg780,
                 reg779,
                 reg778,
                 reg777,
                 reg776,
                 reg775,
                 reg774,
                 reg773,
                 reg772,
                 reg771,
                 reg770,
                 reg769,
                 reg768,
                 wire767,
                 wire766,
                 wire765,
                 wire764,
                 wire763,
                 wire762,
                 wire761,
                 wire760,
                 wire759,
                 wire758,
                 wire757,
                 (1'h0)};
  assign wire757 = ((wire754 ^~ wire753[(3'h6):(1'h0)]) ?
                       (8'haa) : ({((^~wire753) ~^ (~&wire752)), wire754} ?
                           $signed(wire755) : (((wire755 ?
                                   wire755 : (8'ha6)) || $unsigned(wire754)) ?
                               ((wire754 ? wire754 : wire755) ?
                                   (&wire752) : $unsigned((8'ha6))) : $signed(wire752))));
  assign wire758 = wire755[(1'h1):(1'h1)];
  assign wire759 = $signed(wire755[(3'h6):(1'h0)]);
  assign wire760 = (wire755 ? wire752 : wire759);
  assign wire761 = ({(((wire752 ?
                               wire759 : wire760) >> $signed((8'haa))) == wire756),
                           (-wire758[(2'h2):(2'h2)])} ?
                       wire754[(3'h4):(2'h3)] : $signed(wire753));
  assign wire762 = wire755[(2'h3):(1'h1)];
  assign wire763 = {wire755[(1'h1):(1'h1)], wire761[(1'h1):(1'h0)]};
  assign wire764 = ({{wire752, ((wire755 & wire757) << {(8'hbe), wire753})},
                       $signed(($signed(wire754) >>> $unsigned(wire757)))} >>> ($signed(($signed(wire756) ?
                       (wire756 ? wire758 : (8'hba)) : {(8'ha3)})) ^ wire757));
  assign wire765 = (wire763 ?
                       ($signed((wire755 >= (wire761 != (8'haa)))) ?
                           wire764[(4'ha):(3'h6)] : ((wire760 ?
                                   wire762 : wire761) ?
                               wire752[(4'ha):(4'h8)] : wire763[(1'h0):(1'h0)])) : wire752);
  assign wire766 = ($signed(wire755[(3'h5):(2'h3)]) && (wire762[(4'hd):(1'h1)] ?
                       (($signed(wire761) ?
                           (~^wire759) : (wire761 <= (7'h40))) < wire763[(1'h0):(1'h0)]) : $signed($signed(wire752))));
  assign wire767 = (~wire755[(1'h1):(1'h0)]);
  always
    @(posedge clk) begin
      reg768 <= ((($signed((+wire752)) ?
              wire752 : {(~wire755)}) - (wire755[(3'h4):(3'h4)] ?
              wire760 : $unsigned($signed((8'hb7))))) ?
          $unsigned((((wire764 <= wire752) ?
              (+wire753) : (^wire759)) | ((wire764 ? wire753 : (7'h42)) ?
              (^(8'hbb)) : ((7'h44) ?
                  wire761 : (8'hb2))))) : (wire754[(3'h5):(3'h5)] && $unsigned($unsigned(wire757))));
      reg769 <= (wire759 || (^~reg768[(3'h5):(2'h3)]));
      if ($signed((((!wire763) ?
              $unsigned((wire764 ?
                  wire752 : wire758)) : (wire763[(1'h1):(1'h0)] ?
                  (wire758 ~^ (8'haa)) : wire767)) ?
          (wire765[(3'h4):(1'h0)] ?
              wire761[(4'hc):(3'h6)] : (!$unsigned(wire758))) : (^($signed((8'hb9)) ?
              {wire753, wire761} : {wire760, wire753})))))
        begin
          reg770 <= wire755;
          reg771 <= ((wire754[(4'h8):(4'h8)] ?
                  reg768 : $signed($signed((wire753 & wire764)))) ?
              $signed(((^~wire756) ?
                  $signed(reg769) : wire757)) : $signed((^~$unsigned(wire754))));
          reg772 <= (^~$signed(reg770[(4'hb):(3'h7)]));
        end
      else
        begin
          reg770 <= (wire764 ?
              $unsigned({reg771,
                  ((wire758 ? wire755 : wire758) ?
                      {(7'h41), wire766} : {reg770, wire756})}) : (~^(8'hba)));
          if (wire766[(4'hc):(4'h8)])
            begin
              reg771 <= $signed(wire752[(4'he):(2'h2)]);
              reg772 <= (8'ha9);
              reg773 <= $signed(wire764);
              reg774 <= $signed($unsigned(reg773));
            end
          else
            begin
              reg771 <= {wire758, wire759[(1'h1):(1'h0)]};
              reg772 <= (8'ha6);
            end
          reg775 <= {wire752};
        end
      if (wire757[(1'h0):(1'h0)])
        begin
          if ({wire757[(4'hb):(2'h2)]})
            begin
              reg776 <= {$signed($unsigned(({wire756, (8'had)} ?
                      $signed(reg769) : wire764))),
                  reg775[(1'h0):(1'h0)]};
              reg777 <= (((|wire758[(4'h8):(1'h1)]) >>> (($signed(wire752) ?
                          ((8'h9d) ? reg773 : wire759) : (reg769 > reg776)) ?
                      (^$unsigned(wire764)) : {{reg768, wire761}})) ?
                  $signed((-{wire766[(4'h8):(1'h1)],
                      $unsigned((8'hae))})) : (wire767 ?
                      ($unsigned($unsigned(wire758)) ^~ ((reg770 <= (8'hab)) ?
                          (~&reg771) : wire755[(1'h1):(1'h0)])) : ((-{wire755,
                          wire760}) | wire765)));
              reg778 <= wire752[(1'h1):(1'h1)];
              reg779 <= {{$signed($unsigned((~wire764))),
                      $unsigned((~|((8'ha0) ? reg772 : wire759)))},
                  wire752[(3'h7):(1'h0)]};
            end
          else
            begin
              reg776 <= $signed((&(wire753 ?
                  ($unsigned(wire758) ?
                      (8'hbb) : wire756[(2'h3):(1'h0)]) : ((wire756 != wire763) ?
                      wire757 : $unsigned(reg773)))));
              reg777 <= reg773[(3'h4):(2'h3)];
              reg778 <= wire765[(2'h2):(1'h1)];
              reg779 <= ({({$unsigned(wire756),
                          ((8'hab) ?
                              wire764 : wire754)} < (reg771[(3'h4):(1'h0)] ?
                          (wire758 ? (7'h44) : wire757) : reg779))} ?
                  $signed((wire765[(3'h7):(3'h5)] ?
                      ($signed(reg777) - reg772) : {$signed(reg770),
                          reg772})) : {{(~(wire758 ? wire761 : wire762))},
                      reg768});
            end
          if ($signed({reg774, {reg770[(4'he):(3'h7)]}}))
            begin
              reg780 <= {($unsigned($signed(wire763[(2'h2):(1'h0)])) * (reg775 ?
                      (~|$unsigned(wire753)) : ((wire764 <= wire764) >>> reg778)))};
              reg781 <= {($unsigned(((wire756 < reg770) != reg775[(1'h0):(1'h0)])) + wire753[(4'h8):(3'h7)])};
              reg782 <= wire755[(3'h4):(1'h1)];
              reg783 <= $signed(reg773);
            end
          else
            begin
              reg780 <= reg777[(2'h3):(2'h2)];
              reg781 <= ($unsigned((+$unsigned((reg776 ^~ wire763)))) ^~ $unsigned((wire756[(1'h0):(1'h0)] ?
                  reg773[(1'h0):(1'h0)] : reg769[(4'hc):(4'hc)])));
              reg782 <= (+(((^~$signed(wire752)) ?
                  {(^~reg780),
                      (wire757 - reg770)} : (wire754[(2'h3):(1'h1)] + reg780)) + reg783));
            end
          reg784 <= (wire767[(3'h5):(2'h2)] > reg781[(3'h7):(1'h1)]);
          reg785 <= wire759;
          reg786 <= $unsigned({(~^{(^~reg772)})});
        end
      else
        begin
          reg776 <= $unsigned($signed((($unsigned(reg778) >>> reg772) - (~(reg783 <= wire752)))));
          reg777 <= $signed(((!$signed((wire754 ? wire752 : wire757))) ?
              $signed(wire761) : ($unsigned(wire758) ?
                  $signed(((7'h41) - reg776)) : ((~^(8'hbb)) <= (reg775 ?
                      reg777 : wire757)))));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module708
#( parameter param748 = (~&((((7'h44) ? {(8'haa), (8'h9c)} : (~^(8'hb6))) ? (~((8'hab) < (7'h42))) : (((8'ha1) ? (8'hb8) : (8'hb5)) ? (7'h41) : ((8'hbf) ~^ (8'hb2)))) <<< ((((8'h9c) | (8'ha0)) != (~^(8'hbc))) ? (((7'h41) ? (8'hbc) : (8'ha7)) && (^~(8'ha7))) : {(~|(8'ha6))}))) )
(y, clk, wire712, wire711, wire710, wire709);
  output wire [(32'h198):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire712;
  input wire [(5'h13):(1'h0)] wire711;
  input wire signed [(3'h7):(1'h0)] wire710;
  input wire signed [(5'h14):(1'h0)] wire709;
  reg signed [(5'h10):(1'h0)] reg747 = (1'h0);
  reg [(4'he):(1'h0)] reg746 = (1'h0);
  reg signed [(4'he):(1'h0)] reg745 = (1'h0);
  reg [(4'hc):(1'h0)] reg744 = (1'h0);
  reg [(5'h12):(1'h0)] reg743 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg742 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg741 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg740 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg739 = (1'h0);
  reg [(5'h15):(1'h0)] reg738 = (1'h0);
  reg [(2'h2):(1'h0)] reg737 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg736 = (1'h0);
  reg [(5'h13):(1'h0)] reg735 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg734 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg733 = (1'h0);
  reg [(5'h13):(1'h0)] reg732 = (1'h0);
  reg [(3'h7):(1'h0)] reg731 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire730;
  wire [(4'h9):(1'h0)] wire729;
  reg [(4'he):(1'h0)] reg728 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg727 = (1'h0);
  reg [(2'h3):(1'h0)] reg726 = (1'h0);
  reg [(5'h12):(1'h0)] reg725 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg724 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg723 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg722 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg721 = (1'h0);
  reg [(5'h14):(1'h0)] reg720 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg719 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg718 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg717 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg716 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg715 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg714 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire713;
  assign y = {reg747,
                 reg746,
                 reg745,
                 reg744,
                 reg743,
                 reg742,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 wire730,
                 wire729,
                 reg728,
                 reg727,
                 reg726,
                 reg725,
                 reg724,
                 reg723,
                 reg722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 wire713,
                 (1'h0)};
  assign wire713 = $signed($signed((({wire709} ?
                           wire709[(1'h0):(1'h0)] : $unsigned(wire709)) ?
                       $signed((wire712 ? wire710 : wire711)) : wire712)));
  always
    @(posedge clk) begin
      reg714 <= wire709[(4'h9):(3'h6)];
      reg715 <= $signed(wire712[(1'h1):(1'h1)]);
      reg716 <= (wire710[(3'h4):(2'h2)] ?
          $signed(wire710) : $unsigned(reg714[(1'h1):(1'h0)]));
      if (wire713[(1'h0):(1'h0)])
        begin
          reg717 <= reg716;
          reg718 <= $unsigned(reg714);
          reg719 <= ((wire713 >>> ((&$unsigned(reg715)) ?
              wire712 : (8'hac))) || $signed(($signed((^reg716)) * (|reg716[(1'h0):(1'h0)]))));
        end
      else
        begin
          if ({(~^{reg719[(3'h7):(2'h2)], $unsigned(reg718)}), wire711})
            begin
              reg717 <= $signed(((wire713[(1'h1):(1'h1)] ^ $unsigned(((8'ha7) ?
                  reg715 : (8'ha7)))) == reg714[(1'h0):(1'h0)]));
              reg718 <= $unsigned(wire710);
              reg719 <= (($signed(reg714) >> $unsigned(($signed(wire712) ?
                  reg719[(3'h5):(1'h1)] : $unsigned(wire711)))) + $unsigned(reg718));
            end
          else
            begin
              reg717 <= $signed(wire713[(2'h2):(1'h1)]);
              reg718 <= ($signed({(wire713[(1'h0):(1'h0)] - wire711[(1'h1):(1'h0)]),
                      $signed({wire712})}) ?
                  (&(($unsigned(wire710) ?
                          (wire711 <= reg717) : reg716[(2'h3):(1'h1)]) ?
                      $signed((reg715 != wire711)) : $unsigned(wire712))) : reg719);
              reg719 <= reg714[(2'h3):(1'h1)];
              reg720 <= $signed((wire713 * ($unsigned((reg716 < reg714)) ?
                  ((reg715 << wire709) ?
                      (8'haa) : $unsigned(wire709)) : ({reg714} ?
                      (reg718 ? reg717 : reg716) : wire711))));
              reg721 <= (|reg718);
            end
          reg722 <= wire713[(1'h0):(1'h0)];
          reg723 <= (reg719[(3'h4):(1'h1)] * reg714[(2'h2):(1'h1)]);
          if ($signed(($signed((^wire710)) - $unsigned($unsigned($signed(reg716))))))
            begin
              reg724 <= ($unsigned($signed($unsigned($unsigned(wire711)))) >>> (wire713[(1'h0):(1'h0)] ?
                  reg714 : (~&wire711[(1'h0):(1'h0)])));
              reg725 <= (wire713[(2'h3):(1'h1)] ?
                  (^~($unsigned($signed(reg724)) << reg720[(1'h0):(1'h0)])) : (+(-wire712[(4'ha):(3'h5)])));
            end
          else
            begin
              reg724 <= (~({$signed({reg722, reg724}),
                  wire709[(4'h8):(3'h4)]} * (reg719[(3'h6):(3'h6)] ?
                  $unsigned(((8'ha9) ?
                      wire710 : reg723)) : wire710[(3'h6):(3'h6)])));
              reg725 <= $unsigned(((reg714 ?
                      {reg715} : ((~reg718) ?
                          (wire711 ? reg717 : wire712) : $signed(reg722))) ?
                  ($unsigned($unsigned((8'ha5))) ?
                      ($unsigned(reg721) ?
                          $signed(reg723) : (wire711 | (8'hae))) : (wire709 ?
                          reg714[(2'h2):(1'h0)] : $unsigned(reg723))) : wire712[(3'h5):(1'h1)]));
              reg726 <= ($unsigned({$unsigned($unsigned(reg721))}) ^ $unsigned((|(^~$signed(wire713)))));
              reg727 <= (+$signed(((~^reg716) ?
                  {wire710[(3'h4):(2'h2)]} : ($unsigned(reg724) & $unsigned(reg720)))));
            end
        end
      reg728 <= wire713;
    end
  assign wire729 = reg722[(1'h0):(1'h0)];
  assign wire730 = $signed(reg719[(1'h1):(1'h0)]);
  always
    @(posedge clk) begin
      reg731 <= {reg715[(3'h5):(3'h5)]};
      if ((8'h9d))
        begin
          if ($unsigned(({(&(reg725 >>> reg720))} && {$signed(((8'h9f) >> reg727))})))
            begin
              reg732 <= $unsigned((reg726 & $unsigned($signed($signed(reg724)))));
              reg733 <= (~wire712[(4'hc):(3'h5)]);
              reg734 <= (reg715[(1'h0):(1'h0)] >> $signed($signed({(reg727 < (8'hb9)),
                  (^~reg720)})));
            end
          else
            begin
              reg732 <= wire709;
              reg733 <= $signed(reg714);
              reg734 <= reg714;
              reg735 <= {$signed(reg724)};
              reg736 <= ((^~(~^({wire729} > (|reg733)))) ?
                  reg734 : $unsigned((((reg718 + reg734) ^~ ((7'h44) && reg726)) ?
                      {{reg722, (8'hb9)}} : (~|reg725[(3'h7):(3'h6)]))));
            end
          reg737 <= {(reg720 ?
                  reg724[(2'h2):(1'h0)] : ($signed(reg721) >= {(8'hb9)}))};
        end
      else
        begin
          reg732 <= reg735[(5'h11):(4'hd)];
          if (($signed(reg726) ?
              {$signed($signed(wire710)),
                  {$unsigned((reg715 ?
                          reg734 : reg721))}} : (|$signed(reg724[(2'h3):(2'h3)]))))
            begin
              reg733 <= wire730[(4'hb):(2'h3)];
              reg734 <= (~&reg733[(2'h3):(2'h3)]);
              reg735 <= (+((8'hbb) ? reg733[(1'h1):(1'h1)] : (8'hbe)));
              reg736 <= (|(+{($signed(wire730) ?
                      ((7'h42) ? (8'hb8) : reg717) : $unsigned((8'hbf)))}));
            end
          else
            begin
              reg733 <= reg725[(4'he):(4'hb)];
              reg734 <= (~^wire713);
            end
          reg737 <= (~|(reg720 ?
              $signed(((^~reg719) ?
                  (reg737 > reg724) : (~&(8'haf)))) : (~|{reg728[(1'h1):(1'h0)],
                  wire730[(3'h6):(2'h2)]})));
        end
      reg738 <= (!reg720);
      if ((^~(((8'ha1) ~^ ((~^reg721) - (reg738 ?
          (8'ha4) : wire711))) | reg736[(3'h5):(1'h1)])))
        begin
          reg739 <= reg735[(5'h13):(5'h11)];
          reg740 <= (reg714[(1'h1):(1'h0)] ?
              wire729[(4'h9):(2'h3)] : reg738[(3'h4):(1'h1)]);
          if (reg722)
            begin
              reg741 <= $unsigned($signed((($signed(reg723) << $signed(reg736)) ?
                  ((~reg732) >= wire711) : $signed((^(8'ha9))))));
              reg742 <= (^reg714);
              reg743 <= ((~|((reg741 != (reg722 || reg714)) >= {$signed(reg725),
                  reg735})) + (wire730 ? reg716 : $signed(reg720)));
              reg744 <= wire711[(2'h3):(1'h0)];
            end
          else
            begin
              reg741 <= reg732;
              reg742 <= reg739[(4'h8):(4'h8)];
            end
        end
      else
        begin
          if (reg720)
            begin
              reg739 <= (~(^~(8'h9f)));
              reg740 <= $unsigned(wire711[(4'h9):(1'h0)]);
              reg741 <= {wire729[(4'h9):(2'h2)],
                  $unsigned($signed($signed((wire711 ? reg720 : reg717))))};
              reg742 <= (~$unsigned(reg743[(2'h2):(1'h0)]));
              reg743 <= $signed(reg722[(3'h5):(2'h2)]);
            end
          else
            begin
              reg739 <= reg714;
              reg740 <= (8'ha0);
              reg741 <= reg731[(2'h3):(1'h1)];
              reg742 <= (&(({reg725,
                      (reg714 >= reg719)} >> $unsigned((reg726 & reg715))) ?
                  (+(~&reg734[(4'hf):(1'h1)])) : {wire730}));
            end
          if (wire711)
            begin
              reg744 <= (reg718[(4'hf):(3'h5)] ?
                  reg728 : wire710[(3'h4):(2'h3)]);
              reg745 <= (reg719 >> reg737[(2'h2):(1'h1)]);
              reg746 <= (8'ha9);
            end
          else
            begin
              reg744 <= ((~$signed($signed($signed((8'hb2))))) ^~ (~|reg716[(1'h0):(1'h0)]));
              reg745 <= $signed((reg725 ?
                  ((reg724 > $unsigned(reg746)) ?
                      ((reg742 ? reg737 : wire730) ?
                          $unsigned(reg727) : reg741[(4'hb):(3'h7)]) : $signed(wire710[(3'h6):(2'h3)])) : (~($signed((8'hb9)) >> wire729))));
              reg746 <= $signed(reg715[(1'h0):(1'h0)]);
            end
          reg747 <= {$signed({(reg741[(3'h4):(1'h1)] ?
                      $signed(reg743) : (reg719 ? reg719 : wire711)),
                  (^~$unsigned(reg714))}),
              {$signed(wire712)}};
        end
    end
endmodule