(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h13d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire4;
  input wire [(5'h15):(1'h0)] wire3;
  input wire [(5'h15):(1'h0)] wire2;
  input wire signed [(5'h15):(1'h0)] wire1;
  input wire [(5'h14):(1'h0)] wire0;
  wire [(4'h8):(1'h0)] wire1938;
  wire [(5'h13):(1'h0)] wire724;
  wire signed [(5'h11):(1'h0)] wire1940;
  wire signed [(5'h13):(1'h0)] wire1941;
  wire [(4'hb):(1'h0)] wire1942;
  wire signed [(4'h9):(1'h0)] wire1943;
  wire signed [(2'h3):(1'h0)] wire1945;
  reg [(4'he):(1'h0)] reg1946 = (1'h0);
  reg [(5'h14):(1'h0)] reg1947 = (1'h0);
  reg [(3'h7):(1'h0)] reg1948 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1949 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1950 = (1'h0);
  reg [(4'hb):(1'h0)] reg1951 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1952 = (1'h0);
  wire [(5'h11):(1'h0)] wire1953;
  wire signed [(5'h13):(1'h0)] wire1954;
  wire signed [(5'h12):(1'h0)] wire1955;
  wire [(3'h7):(1'h0)] wire1957;
  wire [(4'h8):(1'h0)] wire1959;
  wire [(5'h11):(1'h0)] wire1960;
  wire signed [(3'h7):(1'h0)] wire1961;
  wire signed [(5'h10):(1'h0)] wire1962;
  wire signed [(4'hb):(1'h0)] wire1963;
  assign y = {wire1938,
                 wire724,
                 wire1940,
                 wire1941,
                 wire1942,
                 wire1943,
                 wire1945,
                 reg1946,
                 reg1947,
                 reg1948,
                 reg1949,
                 reg1950,
                 reg1951,
                 reg1952,
                 wire1953,
                 wire1954,
                 wire1955,
                 wire1957,
                 wire1959,
                 wire1960,
                 wire1961,
                 wire1962,
                 wire1963,
                 (1'h0)};
  module5 modinst725 (.wire6(wire4), .wire7(wire1), .wire8(wire2), .y(wire724), .clk(clk), .wire9(wire3));
  module726 modinst1939 (wire1938, clk, wire2, wire3, wire1, wire724, wire0);
  assign wire1940 = wire724[(4'h9):(3'h7)];
  assign wire1941 = wire4;
  assign wire1942 = ((-(8'h9e)) ?
                        {$unsigned($unsigned(wire1938[(1'h0):(1'h0)]))} : $signed((((wire724 ?
                            wire1 : wire3) != $signed(wire3)) ^~ ((wire3 ~^ wire0) > $unsigned(wire2)))));
  module514 modinst1944 (.clk(clk), .wire516(wire1), .y(wire1943), .wire517(wire4), .wire518(wire0), .wire515(wire724));
  assign wire1945 = (-wire1938);
  always
    @(posedge clk) begin
      if (wire1943[(2'h2):(1'h0)])
        begin
          if (wire1942)
            begin
              reg1946 <= $signed(wire724);
            end
          else
            begin
              reg1946 <= (wire3 ?
                  (^~wire1941[(3'h6):(3'h6)]) : $signed({(wire1945 + (^reg1946)),
                      (^(-wire1942))}));
              reg1947 <= {((~(+(~(8'hbb)))) ?
                      (~^$unsigned(wire4[(4'h9):(2'h2)])) : ($signed($signed(wire1943)) ?
                          $unsigned(wire1942) : $unsigned((!wire724)))),
                  (wire2 ? wire1940 : (!$signed((wire1 >= (8'hb1)))))};
              reg1948 <= wire1945;
              reg1949 <= (wire1941 >>> $signed($signed((((8'hb4) && wire1942) ?
                  wire1942 : $unsigned(wire724)))));
              reg1950 <= {(8'hab)};
            end
          reg1951 <= wire1945[(2'h3):(2'h2)];
          reg1952 <= reg1949;
        end
      else
        begin
          reg1946 <= (~&((($unsigned(wire1) <= $signed(wire1940)) ?
              $signed((reg1949 ? (8'hae) : wire3)) : reg1950) ~^ reg1946));
          if ((8'ha0))
            begin
              reg1947 <= $signed({((reg1949[(4'he):(4'hc)] ?
                      $unsigned(reg1950) : (+wire1940)) && {(wire1 ?
                          reg1950 : wire1943)}),
                  {({wire2} + (wire1945 - wire2))}});
              reg1948 <= (+{(~(-(^~(8'h9d)))), (-$unsigned((~&(8'hae))))});
              reg1949 <= $unsigned(wire1940[(4'h8):(3'h7)]);
              reg1950 <= (wire1941[(4'h9):(3'h4)] != wire1938[(1'h1):(1'h1)]);
            end
          else
            begin
              reg1947 <= wire724;
              reg1948 <= ($signed(wire3[(4'h9):(3'h4)]) ?
                  $unsigned((-wire1943)) : ((reg1951[(1'h1):(1'h0)] * ((!(8'hb9)) >> {(8'h9f),
                      wire1941})) ^ $unsigned($unsigned($unsigned(wire1938)))));
              reg1949 <= {wire0, (&wire724[(4'h8):(2'h2)])};
            end
        end
    end
  assign wire1953 = $signed(wire1945[(1'h0):(1'h0)]);
  assign wire1954 = {wire2, $unsigned($signed(reg1949[(3'h7):(3'h4)]))};
  module218 modinst1956 (wire1955, clk, reg1950, wire1954, wire724, wire1941);
  module514 modinst1958 (.y(wire1957), .wire518(wire0), .clk(clk), .wire515(reg1950), .wire517(wire1953), .wire516(reg1947));
  assign wire1959 = wire0;
  assign wire1960 = reg1950;
  assign wire1961 = {$signed($signed(wire1953[(3'h6):(3'h4)]))};
  assign wire1962 = wire1941[(5'h11):(4'hc)];
  module759 modinst1964 (.wire764(wire1940), .clk(clk), .wire761(wire1938), .wire760(wire1943), .wire762(wire1955), .y(wire1963), .wire763(reg1951));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module726
#( parameter param1937 = (~&({({(8'hbb)} != (8'ha9))} ? (^~(((8'hbd) ? (8'ha3) : (8'hb0)) | (^~(8'hbf)))) : ({(~&(8'hb4)), ((8'ha8) ? (8'hbf) : (8'h9e))} > (((8'hb4) & (8'h9c)) ? ((8'hb1) ? (8'hb8) : (8'ha5)) : ((8'ha4) ? (8'ha0) : (8'ha9)))))) )
(y, clk, wire731, wire730, wire729, wire728, wire727);
  output wire [(32'hd5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire731;
  input wire signed [(5'h15):(1'h0)] wire730;
  input wire signed [(5'h15):(1'h0)] wire729;
  input wire [(5'h10):(1'h0)] wire728;
  input wire signed [(5'h10):(1'h0)] wire727;
  reg signed [(4'h9):(1'h0)] reg1936 = (1'h0);
  reg [(4'he):(1'h0)] reg1935 = (1'h0);
  reg [(4'h9):(1'h0)] reg1934 = (1'h0);
  reg [(3'h5):(1'h0)] reg1933 = (1'h0);
  reg [(4'he):(1'h0)] reg1932 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1931 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1930 = (1'h0);
  reg [(5'h10):(1'h0)] reg1929 = (1'h0);
  reg [(4'hf):(1'h0)] reg1928 = (1'h0);
  reg [(3'h4):(1'h0)] reg1927 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1926 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1925 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire1924;
  wire signed [(5'h10):(1'h0)] wire1923;
  wire signed [(5'h13):(1'h0)] wire1915;
  wire signed [(5'h15):(1'h0)] wire732;
  wire signed [(4'ha):(1'h0)] wire1917;
  wire signed [(2'h2):(1'h0)] wire1918;
  wire [(5'h11):(1'h0)] wire1919;
  wire signed [(2'h3):(1'h0)] wire1921;
  assign y = {reg1936,
                 reg1935,
                 reg1934,
                 reg1933,
                 reg1932,
                 reg1931,
                 reg1930,
                 reg1929,
                 reg1928,
                 reg1927,
                 reg1926,
                 reg1925,
                 wire1924,
                 wire1923,
                 wire1915,
                 wire732,
                 wire1917,
                 wire1918,
                 wire1919,
                 wire1921,
                 (1'h0)};
  assign wire732 = ((-wire728[(4'h8):(3'h4)]) ?
                       $signed((wire731[(1'h0):(1'h0)] ?
                           $signed((wire729 + wire727)) : ((-wire730) ^~ (wire729 || (8'haa))))) : ((wire729[(3'h7):(2'h2)] < wire729) ?
                           $signed({$unsigned((8'hba)),
                               {wire731}}) : (wire729[(4'he):(4'ha)] << $signed((~^wire729)))));
  module733 modinst1916 (wire1915, clk, wire727, wire732, wire730, wire729, wire731);
  assign wire1917 = wire732;
  assign wire1918 = {$signed((&(|{(8'haa)})))};
  module1445 modinst1920 (wire1919, clk, wire732, wire1917, wire728, wire727);
  module950 modinst1922 (wire1921, clk, wire728, wire732, wire729, wire1919, wire727);
  assign wire1923 = wire1917;
  assign wire1924 = (({wire728[(4'hb):(4'hb)]} - $unsigned($unsigned($signed((8'hba))))) ?
                        $signed((~&$signed((wire731 * wire727)))) : $signed({{$unsigned(wire730)}}));
  always
    @(posedge clk) begin
      if (wire727[(4'he):(2'h2)])
        begin
          reg1925 <= $unsigned(wire728);
          reg1926 <= wire1919;
        end
      else
        begin
          reg1925 <= wire1923[(2'h2):(2'h2)];
          reg1926 <= $unsigned((wire1915 != (!$signed((wire731 ?
              wire730 : wire1923)))));
        end
      if (($unsigned(wire1921) ~^ ($unsigned(wire727[(3'h4):(2'h2)]) * $unsigned(wire732))))
        begin
          if (((reg1926[(2'h2):(1'h1)] ^~ ((wire730 * (~^wire1923)) << (!(wire1918 != wire729)))) ?
              reg1925[(4'h8):(3'h7)] : (((wire1918[(2'h2):(2'h2)] | $signed(reg1925)) <= {(&wire1921),
                      wire1915[(4'hf):(4'hd)]}) ?
                  {((&wire730) == (wire729 - wire1924))} : (^~$unsigned((reg1925 ?
                      (8'hb6) : wire1919))))))
            begin
              reg1927 <= ((|wire730) == wire1924);
              reg1928 <= wire1917;
              reg1929 <= (~^(^~wire1921));
              reg1930 <= wire732[(4'he):(4'ha)];
              reg1931 <= wire730;
            end
          else
            begin
              reg1927 <= (~|(-(reg1929 ^ {(reg1929 ? (8'hbb) : wire1915)})));
              reg1928 <= (8'ha3);
            end
          if (($signed(($unsigned((wire730 ?
              wire1921 : (8'ha0))) & $unsigned($unsigned(wire1921)))) ~^ wire727[(4'hf):(4'hc)]))
            begin
              reg1932 <= wire1918[(1'h1):(1'h0)];
            end
          else
            begin
              reg1932 <= $signed(reg1929[(3'h7):(3'h5)]);
              reg1933 <= $unsigned((8'ha7));
              reg1934 <= wire731;
              reg1935 <= ($signed($unsigned($signed(wire729[(3'h4):(1'h1)]))) ?
                  wire1923[(4'hb):(3'h7)] : $unsigned($signed((-((8'hba) ^ wire730)))));
              reg1936 <= ($unsigned(wire728[(4'he):(4'h9)]) >>> reg1929[(2'h3):(1'h0)]);
            end
        end
      else
        begin
          reg1927 <= ($unsigned(reg1929[(4'he):(3'h4)]) >> (wire1917 >>> $unsigned($unsigned((reg1929 - wire1919)))));
          reg1928 <= {reg1935, (&wire1917)};
          reg1929 <= wire1915;
          if ($unsigned($signed((($unsigned(reg1935) || (&wire1915)) >>> $unsigned(reg1934[(1'h0):(1'h0)])))))
            begin
              reg1930 <= (~|($unsigned($signed(reg1933)) ?
                  $signed((wire732[(3'h4):(1'h0)] - {wire728,
                      reg1935})) : ($unsigned(reg1929) ?
                      $signed((^~(8'hb7))) : ($signed(reg1933) ^~ reg1928))));
            end
          else
            begin
              reg1930 <= $signed($signed($unsigned({wire728[(1'h0):(1'h0)]})));
              reg1931 <= (reg1929 * ($signed($signed($unsigned(reg1928))) ?
                  $unsigned((wire1923 >> wire727)) : $unsigned(reg1930[(4'h9):(3'h5)])));
              reg1932 <= (wire1923 ?
                  {$unsigned(wire731)} : ($unsigned(reg1929[(4'hb):(3'h4)]) ?
                      (wire1919 ?
                          ((wire731 >>> wire731) ?
                              (reg1926 >= wire1918) : ((8'hb4) ?
                                  reg1933 : reg1927)) : ($signed((8'ha7)) ?
                              wire730 : wire729[(4'h8):(3'h5)])) : wire730));
              reg1933 <= wire1919[(1'h0):(1'h0)];
              reg1934 <= $signed((reg1931[(1'h0):(1'h0)] || reg1928));
            end
          if ((reg1929 * ((~&$signed((^reg1925))) >> (wire1918 == $signed(wire1924[(2'h3):(1'h1)])))))
            begin
              reg1935 <= (((($unsigned(wire1919) ~^ wire730) - (+wire1923[(4'hf):(4'ha)])) ?
                      {({(8'hb1)} > (wire1917 << (8'ha7))),
                          reg1927[(2'h3):(1'h0)]} : {reg1933}) ?
                  wire1923 : ({($signed(reg1925) ?
                              (reg1927 * reg1926) : $signed(wire728))} ?
                      {reg1933[(1'h0):(1'h0)],
                          wire1915} : (!reg1926[(2'h3):(2'h3)])));
              reg1936 <= ((reg1930 ?
                      (wire1918[(1'h0):(1'h0)] ?
                          (+$unsigned(wire728)) : reg1936[(4'h9):(2'h2)]) : wire730) ?
                  (-(|(^((7'h43) >>> (8'hac))))) : $unsigned((reg1933 ?
                      {(^~wire1915),
                          $signed(wire1921)} : wire729[(5'h10):(4'ha)])));
            end
          else
            begin
              reg1935 <= (wire1919 <= {(7'h40)});
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module5
#( parameter param723 = (~&(({(7'h44)} <<< ((|(8'haf)) >= {(8'h9c)})) ? {(^~(~|(7'h43))), (~|((8'ha5) ? (7'h40) : (8'hae)))} : ((~((8'ha5) <= (8'ha6))) | ({(8'hbd)} ^~ {(8'ha5)})))) )
(y, clk, wire9, wire8, wire7, wire6);
  output wire [(32'h68):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire9;
  input wire [(5'h15):(1'h0)] wire8;
  input wire [(5'h13):(1'h0)] wire7;
  input wire [(4'ha):(1'h0)] wire6;
  reg signed [(5'h14):(1'h0)] reg722 = (1'h0);
  reg [(5'h14):(1'h0)] reg721 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg720 = (1'h0);
  reg [(3'h4):(1'h0)] reg719 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg718 = (1'h0);
  reg [(3'h5):(1'h0)] reg717 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg716 = (1'h0);
  wire [(2'h2):(1'h0)] wire715;
  wire signed [(4'hd):(1'h0)] wire713;
  wire [(4'hd):(1'h0)] wire10;
  assign y = {reg722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 reg716,
                 wire715,
                 wire713,
                 wire10,
                 (1'h0)};
  assign wire10 = $signed((wire8 ^ wire7));
  module11 modinst714 (wire713, clk, wire7, wire9, wire6, wire8);
  assign wire715 = $signed(wire9[(5'h13):(2'h2)]);
  always
    @(posedge clk) begin
      reg716 <= ($unsigned((~^wire713[(1'h1):(1'h0)])) <= $unsigned((wire10[(3'h6):(3'h6)] || ((wire715 ?
          wire6 : wire10) >>> (wire9 ? wire6 : wire715)))));
      if ($signed(((-wire713) << ((!$unsigned(wire7)) << (+(&wire8))))))
        begin
          reg717 <= (^$unsigned(($signed(wire10) ?
              ($signed((8'ha2)) ~^ (reg716 && wire8)) : ($unsigned((8'hae)) ?
                  wire10[(4'hc):(4'hc)] : {wire713}))));
          reg718 <= $signed(wire8[(5'h12):(4'hf)]);
          reg719 <= $unsigned(reg716);
          reg720 <= $unsigned($unsigned(((+$signed(wire7)) ?
              (wire6[(4'ha):(1'h1)] ?
                  $unsigned(reg719) : wire6) : $signed($signed(reg717)))));
          reg721 <= (~&wire713[(4'hb):(3'h5)]);
        end
      else
        begin
          reg717 <= (8'ha3);
          if ((^wire713))
            begin
              reg718 <= ($unsigned($signed(reg716[(2'h3):(1'h0)])) ?
                  (wire9[(4'hb):(2'h3)] ?
                      wire7 : wire8[(1'h0):(1'h0)]) : (reg718 ?
                      $unsigned((7'h41)) : $signed(reg716[(1'h0):(1'h0)])));
              reg719 <= ($unsigned((((~&reg721) ?
                      reg721[(5'h10):(4'h8)] : $unsigned((8'hbd))) <= {(+reg721)})) ?
                  (&($unsigned($signed(reg716)) << reg719)) : (7'h43));
              reg720 <= (&(reg717[(2'h3):(2'h2)] != {reg716,
                  wire9[(3'h6):(2'h3)]}));
              reg721 <= {{{$unsigned($unsigned(reg716)),
                          wire7[(3'h5):(1'h0)]}}};
              reg722 <= $signed($signed(((reg718[(2'h2):(2'h2)] * $signed(reg721)) ?
                  wire10 : {(reg717 ~^ wire8), ((8'had) & reg716)})));
            end
          else
            begin
              reg718 <= $signed((+$unsigned({reg721[(1'h0):(1'h0)]})));
              reg719 <= $unsigned((!(-$signed($signed(wire6)))));
              reg720 <= (reg718[(1'h1):(1'h0)] && $unsigned(wire713[(4'hb):(4'h8)]));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module11
#( parameter param711 = ({({(&(8'had))} ? (((8'h9f) ? (8'hb5) : (8'haa)) >= ((7'h41) > (8'hb6))) : {{(8'ha2)}})} && (-((((8'hb2) ? (8'ha3) : (8'hbd)) >> (8'hbd)) ? (((8'hb2) && (8'hba)) ? ((7'h43) ^ (8'hba)) : (&(7'h43))) : (^~((8'hab) || (8'hb3))))))
, parameter param712 = {{param711, param711}} )
(y, clk, wire15, wire14, wire13, wire12);
  output wire [(32'h187):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire15;
  input wire signed [(5'h14):(1'h0)] wire14;
  input wire signed [(2'h2):(1'h0)] wire13;
  input wire [(4'ha):(1'h0)] wire12;
  wire signed [(5'h11):(1'h0)] wire710;
  wire signed [(2'h2):(1'h0)] wire709;
  wire [(3'h6):(1'h0)] wire708;
  wire signed [(4'h9):(1'h0)] wire707;
  reg signed [(4'he):(1'h0)] reg706 = (1'h0);
  reg [(2'h3):(1'h0)] reg705 = (1'h0);
  reg [(5'h10):(1'h0)] reg704 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg703 = (1'h0);
  reg [(5'h13):(1'h0)] reg702 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg701 = (1'h0);
  reg [(4'hd):(1'h0)] reg700 = (1'h0);
  reg [(4'ha):(1'h0)] reg699 = (1'h0);
  wire [(4'ha):(1'h0)] wire697;
  wire signed [(5'h15):(1'h0)] wire435;
  wire signed [(3'h4):(1'h0)] wire433;
  reg signed [(5'h15):(1'h0)] reg308 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg307 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire306;
  wire signed [(5'h10):(1'h0)] wire305;
  wire [(5'h13):(1'h0)] wire304;
  wire [(5'h14):(1'h0)] wire303;
  wire signed [(4'ha):(1'h0)] wire302;
  wire signed [(3'h5):(1'h0)] wire301;
  wire signed [(5'h13):(1'h0)] wire300;
  reg [(5'h13):(1'h0)] reg299 = (1'h0);
  wire [(5'h14):(1'h0)] wire298;
  wire [(5'h10):(1'h0)] wire296;
  wire signed [(4'ha):(1'h0)] wire18;
  wire signed [(5'h15):(1'h0)] wire17;
  wire signed [(3'h6):(1'h0)] wire16;
  assign y = {wire710,
                 wire709,
                 wire708,
                 wire707,
                 reg706,
                 reg705,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 reg699,
                 wire697,
                 wire435,
                 wire433,
                 reg308,
                 reg307,
                 wire306,
                 wire305,
                 wire304,
                 wire303,
                 wire302,
                 wire301,
                 wire300,
                 reg299,
                 wire298,
                 wire296,
                 wire18,
                 wire17,
                 wire16,
                 (1'h0)};
  assign wire16 = (8'had);
  assign wire17 = (-$signed((|(wire15[(2'h3):(1'h1)] > $signed(wire15)))));
  assign wire18 = (~$unsigned(((wire14[(1'h1):(1'h0)] ?
                      wire12 : $unsigned((8'hb5))) ~^ $signed(wire15[(1'h1):(1'h1)]))));
  module19 modinst297 (wire296, clk, wire18, wire14, wire15, wire16);
  assign wire298 = wire13[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg299 <= (wire16[(2'h2):(1'h1)] < wire17);
    end
  assign wire300 = reg299;
  assign wire301 = $signed((&(+wire18)));
  assign wire302 = wire18[(1'h1):(1'h1)];
  assign wire303 = wire300[(4'hc):(2'h3)];
  assign wire304 = wire302[(2'h3):(2'h3)];
  assign wire305 = ($signed({wire12[(3'h6):(2'h3)], {wire13[(1'h1):(1'h0)]}}) ?
                       $signed(wire303[(1'h0):(1'h0)]) : ($signed(wire302[(2'h2):(1'h0)]) ?
                           (^((^~wire303) ?
                               $signed(wire302) : wire15[(5'h10):(4'he)])) : $unsigned($signed($unsigned(wire17)))));
  assign wire306 = (~&(~^$signed($signed(wire16))));
  always
    @(posedge clk) begin
      reg307 <= wire18[(4'h8):(3'h5)];
      reg308 <= {($unsigned((!reg307[(2'h3):(2'h3)])) ^ ((-(wire300 ?
              wire298 : wire305)) * (~|(reg307 == wire12)))),
          $signed($signed($unsigned((wire304 * wire306))))};
    end
  module309 modinst434 (wire433, clk, wire14, wire303, wire304, reg308);
  assign wire435 = $unsigned(wire304[(2'h3):(2'h2)]);
  module436 modinst698 (wire697, clk, wire304, reg308, reg299, wire296);
  always
    @(posedge clk) begin
      reg699 <= (|$signed($unsigned(((wire14 ? wire296 : wire298) ?
          $unsigned(reg299) : $unsigned(wire303)))));
      if ($unsigned($unsigned(reg699)))
        begin
          if (wire296[(4'ha):(1'h0)])
            begin
              reg700 <= (~{wire13});
              reg701 <= wire296[(2'h2):(1'h0)];
              reg702 <= {(^~$signed($signed((!wire14)))), $unsigned(wire300)};
            end
          else
            begin
              reg700 <= (~$signed((wire12 ?
                  wire433[(2'h3):(1'h1)] : $signed($signed(wire16)))));
            end
          reg703 <= (+reg699[(4'h9):(3'h4)]);
          reg704 <= reg307[(4'hb):(3'h6)];
          reg705 <= $signed(wire300[(4'ha):(1'h0)]);
        end
      else
        begin
          reg700 <= reg704[(2'h2):(2'h2)];
          reg701 <= reg702[(4'ha):(3'h4)];
        end
      reg706 <= (~((8'ha2) > wire15[(4'ha):(3'h6)]));
    end
  assign wire707 = $unsigned((({{wire304, (8'ha3)}, wire435[(1'h1):(1'h1)]} ?
                       {((8'ha8) << (8'hbd))} : wire305[(2'h2):(1'h1)]) != {($unsigned(reg701) ^ $signed(reg700))}));
  assign wire708 = $signed(({$unsigned(wire306),
                           (reg705[(1'h1):(1'h1)] ?
                               $signed(wire300) : (8'ha4))} ?
                       (((reg699 == (8'ha5)) ? wire435 : {wire303, wire435}) ?
                           {$signed((8'ha5)),
                               $signed(wire15)} : $signed(wire306)) : $signed($signed($unsigned(wire12)))));
  assign wire709 = ($unsigned((reg705 == ((wire305 && reg702) ?
                       $unsigned(reg701) : (reg700 - wire16)))) & reg706);
  assign wire710 = $signed(($unsigned(wire16) + $signed(($signed(wire707) ?
                       (reg299 && reg699) : reg700[(4'hc):(3'h7)]))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module436  (y, clk, wire440, wire439, wire438, wire437);
  output wire [(32'h249):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire440;
  input wire signed [(4'hd):(1'h0)] wire439;
  input wire signed [(5'h13):(1'h0)] wire438;
  input wire [(4'hf):(1'h0)] wire437;
  reg signed [(5'h10):(1'h0)] reg696 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg695 = (1'h0);
  reg [(4'h9):(1'h0)] reg694 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg693 = (1'h0);
  reg [(4'h9):(1'h0)] reg692 = (1'h0);
  wire [(3'h5):(1'h0)] wire691;
  wire signed [(4'h8):(1'h0)] wire690;
  reg signed [(5'h15):(1'h0)] reg689 = (1'h0);
  reg [(4'hb):(1'h0)] reg688 = (1'h0);
  reg [(5'h10):(1'h0)] reg687 = (1'h0);
  wire [(4'h9):(1'h0)] wire685;
  reg signed [(5'h11):(1'h0)] reg476 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg475 = (1'h0);
  reg [(5'h15):(1'h0)] reg474 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg473 = (1'h0);
  reg [(4'hf):(1'h0)] reg472 = (1'h0);
  reg [(3'h6):(1'h0)] reg471 = (1'h0);
  reg [(5'h13):(1'h0)] reg470 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg469 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg468 = (1'h0);
  reg [(5'h13):(1'h0)] reg467 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg466 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire465;
  wire signed [(4'h9):(1'h0)] wire464;
  reg signed [(3'h6):(1'h0)] reg463 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg462 = (1'h0);
  reg [(4'hf):(1'h0)] reg461 = (1'h0);
  reg [(3'h4):(1'h0)] reg460 = (1'h0);
  reg [(5'h11):(1'h0)] reg459 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg457 = (1'h0);
  reg signed [(4'he):(1'h0)] reg456 = (1'h0);
  reg [(3'h6):(1'h0)] reg455 = (1'h0);
  reg [(2'h3):(1'h0)] reg454 = (1'h0);
  reg [(4'hf):(1'h0)] reg453 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg452 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg451 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg450 = (1'h0);
  wire [(4'hc):(1'h0)] wire449;
  wire signed [(5'h15):(1'h0)] wire448;
  wire signed [(5'h12):(1'h0)] wire447;
  wire [(4'hf):(1'h0)] wire446;
  wire [(4'ha):(1'h0)] wire445;
  reg signed [(5'h12):(1'h0)] reg444 = (1'h0);
  reg [(5'h12):(1'h0)] reg443 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire442;
  wire signed [(4'h8):(1'h0)] wire441;
  assign y = {reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 wire691,
                 wire690,
                 reg689,
                 reg688,
                 reg687,
                 wire685,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 wire465,
                 wire464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 wire449,
                 wire448,
                 wire447,
                 wire446,
                 wire445,
                 reg444,
                 reg443,
                 wire442,
                 wire441,
                 (1'h0)};
  assign wire441 = {$signed($signed($unsigned(wire440[(1'h1):(1'h0)]))),
                       $unsigned($unsigned($unsigned(wire440)))};
  assign wire442 = ((&($unsigned($signed((8'ha8))) ?
                           wire439[(4'h8):(1'h1)] : $signed(((8'h9e) ?
                               wire440 : wire437)))) ?
                       wire437[(4'hf):(3'h4)] : $unsigned($signed($unsigned($unsigned(wire439)))));
  always
    @(posedge clk) begin
      reg443 <= ($signed((~^wire440[(2'h3):(1'h1)])) & (&(($unsigned((8'h9d)) < wire440) ^~ $signed((wire438 ?
          wire439 : wire438)))));
    end
  always
    @(posedge clk) begin
      reg444 <= (|(|$signed($unsigned($unsigned(wire439)))));
    end
  assign wire445 = (8'haf);
  assign wire446 = ($unsigned(({{wire437}} * {wire441[(1'h1):(1'h0)],
                           wire442})) ?
                       $signed($unsigned(((wire440 <<< reg444) || {wire445,
                           reg444}))) : reg444[(4'hc):(3'h5)]);
  assign wire447 = $unsigned(((wire438[(2'h2):(1'h1)] ?
                           wire438 : {$unsigned(reg444), wire439}) ?
                       $unsigned($unsigned({wire442})) : $signed($unsigned((wire442 - wire440)))));
  assign wire448 = wire442[(1'h0):(1'h0)];
  assign wire449 = (reg443[(3'h5):(1'h0)] << $signed((^(reg444[(1'h1):(1'h0)] ?
                       wire446 : (wire446 << wire437)))));
  always
    @(posedge clk) begin
      if (wire439[(1'h0):(1'h0)])
        begin
          reg450 <= reg443[(4'he):(2'h3)];
          reg451 <= $signed($signed({(wire439 ~^ reg450[(1'h0):(1'h0)])}));
          reg452 <= $unsigned(wire448[(2'h2):(1'h1)]);
          if ($signed(((!reg452) ?
              ((^reg452) ?
                  wire445 : (wire449[(2'h2):(1'h1)] ?
                      (wire445 ? wire447 : wire448) : (wire441 ?
                          wire448 : wire448))) : $signed((~&wire439)))))
            begin
              reg453 <= $unsigned((+(^($unsigned(wire437) < (wire441 ?
                  wire438 : reg443)))));
              reg454 <= ({((wire439 && (~reg453)) > {(8'hba)})} == (~&$signed($signed(wire442))));
              reg455 <= (~($signed((((8'hbe) < (8'hbd)) != ((8'hab) ?
                      wire445 : reg450))) ?
                  ($unsigned({wire449}) | (~|wire446[(1'h1):(1'h0)])) : wire437));
              reg456 <= $signed($unsigned(wire438));
              reg457 <= {reg451[(2'h3):(1'h0)]};
            end
          else
            begin
              reg453 <= (wire445 ?
                  (|wire437) : $signed($signed(reg450[(4'hc):(3'h5)])));
              reg454 <= (wire441 ?
                  {{wire438[(2'h2):(2'h2)],
                          wire441}} : (&$unsigned(($unsigned(reg450) ?
                      $signed(wire445) : (reg443 <= reg452)))));
              reg455 <= wire449;
              reg456 <= $signed((reg453 ? reg444 : wire448));
              reg457 <= (($signed(($unsigned(wire448) > (wire439 ?
                      reg454 : reg456))) ?
                  ($unsigned((reg453 ?
                      reg443 : wire437)) - {$signed(wire440)}) : {{(~|(7'h40))}}) == (reg452 ?
                  $unsigned(reg443) : wire449));
            end
        end
      else
        begin
          reg450 <= wire438[(3'h5):(2'h2)];
          reg451 <= (wire447 ?
              $signed(reg443[(1'h1):(1'h1)]) : wire442[(3'h4):(2'h2)]);
        end
      if (wire439)
        begin
          if (((^~{wire449[(4'hc):(1'h1)],
              $signed(wire449)}) << ((|{$signed(reg450)}) ?
              $signed(reg443[(4'hd):(1'h1)]) : $signed($signed($unsigned(reg452))))))
            begin
              reg458 <= (|$unsigned($signed({reg456[(2'h2):(1'h1)],
                  (reg443 ? wire445 : reg457)})));
              reg459 <= (~&(reg455[(1'h1):(1'h1)] ?
                  wire449[(3'h7):(3'h7)] : $unsigned({$signed(reg454)})));
              reg460 <= ($signed((-reg458)) ?
                  reg443 : ((&(|reg450[(3'h6):(2'h2)])) ?
                      (((7'h42) > reg444[(5'h12):(2'h3)]) && $unsigned($signed(wire445))) : $unsigned($unsigned((wire441 - reg451)))));
              reg461 <= $unsigned(wire437);
              reg462 <= reg459;
            end
          else
            begin
              reg458 <= (|reg459);
              reg459 <= ((^{(reg451[(1'h1):(1'h0)] ?
                          reg450[(5'h10):(2'h2)] : reg458[(3'h4):(1'h0)])}) ?
                  {$signed((wire441[(3'h5):(2'h3)] ?
                          (wire440 >= (8'hb2)) : (+reg459)))} : (7'h42));
              reg460 <= reg458;
              reg461 <= ((reg450[(4'hd):(3'h6)] - wire449) < ($signed({(8'hb4)}) ?
                  wire448 : ((wire445 >= ((8'hb6) >> reg459)) && {$signed(wire445),
                      (reg455 == reg455)})));
              reg462 <= (((8'hbe) ?
                      (wire438 || {reg444}) : $signed($unsigned((8'hae)))) ?
                  (^~((~^$signed(reg444)) << wire447[(4'hc):(4'ha)])) : $signed($signed(reg456)));
            end
        end
      else
        begin
          if ($signed({(($signed((8'hb4)) ^~ reg454[(2'h2):(1'h0)]) ?
                  {(reg450 ? wire438 : (8'hbb))} : reg458)}))
            begin
              reg458 <= reg457[(5'h11):(5'h11)];
              reg459 <= wire446;
              reg460 <= (~&(wire440 ^ $signed($signed(((8'h9d) == reg462)))));
              reg461 <= $signed(reg460[(3'h4):(3'h4)]);
            end
          else
            begin
              reg458 <= $signed(((~^reg456[(2'h2):(1'h0)]) ?
                  ($unsigned($unsigned(wire449)) <<< ($signed(reg454) > $unsigned(reg444))) : reg444));
              reg459 <= $unsigned(((-(!(~|reg451))) ?
                  reg461 : $signed((7'h44))));
            end
          if ($signed(reg454[(1'h1):(1'h0)]))
            begin
              reg462 <= $signed(wire448);
            end
          else
            begin
              reg462 <= $signed($signed($signed($signed(wire438))));
            end
          reg463 <= $unsigned(reg462[(4'he):(3'h5)]);
        end
    end
  assign wire464 = $signed(reg461);
  assign wire465 = $unsigned(reg459);
  always
    @(posedge clk) begin
      if (wire441)
        begin
          reg466 <= $signed(((8'ha0) ?
              (wire445 ?
                  $signed((^(8'ha1))) : $signed(((7'h40) ?
                      wire446 : wire447))) : $signed((^$unsigned((8'haa))))));
        end
      else
        begin
          if ((($signed(wire438[(2'h3):(2'h3)]) ?
              ((^~wire448) & $signed((~|wire464))) : ($signed(reg461[(4'hf):(3'h6)]) ?
                  {(reg463 - reg463)} : {$unsigned(wire442),
                      $signed(reg461)})) - wire440))
            begin
              reg466 <= $signed(((+wire448) >>> ($unsigned((wire437 ?
                  wire445 : wire441)) < $signed((|reg456)))));
            end
          else
            begin
              reg466 <= $signed($signed($unsigned(reg463[(2'h2):(1'h0)])));
              reg467 <= reg459[(1'h1):(1'h1)];
              reg468 <= $unsigned($unsigned(reg467[(4'h9):(3'h4)]));
              reg469 <= (~&$signed($signed((reg454 ?
                  (~&(8'hb4)) : (reg453 ? (8'ha7) : (8'hbf))))));
            end
          if (($signed(reg452) ?
              reg453 : ((((+wire465) <= (~reg460)) ?
                  ((reg458 < wire448) || (reg451 == (8'ha5))) : $unsigned($unsigned(reg454))) ^ {$signed(reg469[(3'h4):(2'h3)])})))
            begin
              reg470 <= reg462[(1'h0):(1'h0)];
              reg471 <= $signed(reg451[(3'h6):(2'h2)]);
            end
          else
            begin
              reg470 <= wire445[(2'h2):(1'h1)];
              reg471 <= reg454;
              reg472 <= {((reg451 ?
                      $unsigned($unsigned(reg459)) : (((8'ha1) ?
                              wire446 : reg459) ?
                          (reg451 || wire438) : $signed(wire449))) == ({reg471[(1'h1):(1'h0)],
                      reg461} << reg463)),
                  {reg452}};
              reg473 <= (|$unsigned(reg460));
            end
          reg474 <= $signed((^reg471));
          reg475 <= $signed((8'hb4));
        end
      reg476 <= $signed({(~^wire448)});
    end
  module477 modinst686 (wire685, clk, wire438, reg466, wire440, reg450);
  always
    @(posedge clk) begin
      reg687 <= wire442;
      reg688 <= reg458[(2'h2):(1'h0)];
      reg689 <= $signed((~|wire464[(3'h4):(2'h2)]));
    end
  assign wire690 = $signed(((((reg470 ^ reg472) && ((8'hb3) * reg462)) ?
                           reg461 : (~&$unsigned(reg467))) ?
                       {$unsigned($signed(reg453)),
                           $unsigned(reg475[(1'h1):(1'h0)])} : ($signed({(8'ha7),
                               reg687}) ?
                           ((wire441 ? wire448 : reg454) ?
                               (wire465 ?
                                   wire447 : reg455) : (reg450 ^ reg458)) : $unsigned((reg453 << reg462)))));
  assign wire691 = reg460[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg692 <= $unsigned({$unsigned((~&(wire464 ? reg444 : reg450)))});
      reg693 <= ({((wire690 ? reg472 : (reg466 >= (7'h43))) ?
                  (wire690[(3'h6):(2'h3)] ?
                      reg474[(4'hd):(3'h4)] : ((8'had) ?
                          reg466 : reg459)) : reg475[(4'h8):(3'h7)]),
              wire437} ?
          reg469[(2'h2):(1'h0)] : $unsigned($unsigned(wire442)));
      reg694 <= reg454;
      reg695 <= reg473;
      reg696 <= (~|({({reg458, reg454} ?
              $unsigned(reg472) : reg466)} ^ wire445));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module309
#( parameter param431 = (~{{(7'h44)}, {({(8'haa)} ? (+(8'hb3)) : ((8'hae) ? (8'h9c) : (7'h42)))}})
, parameter param432 = (((param431 <<< (+param431)) & (|(!param431))) ? (param431 ? param431 : (((8'ha5) - (param431 ? param431 : param431)) >>> (~^(param431 ? param431 : param431)))) : param431) )
(y, clk, wire313, wire312, wire311, wire310);
  output wire [(32'hc3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire313;
  input wire [(5'h14):(1'h0)] wire312;
  input wire [(5'h13):(1'h0)] wire311;
  input wire [(5'h15):(1'h0)] wire310;
  wire signed [(5'h11):(1'h0)] wire430;
  wire signed [(4'hc):(1'h0)] wire429;
  wire signed [(4'h9):(1'h0)] wire428;
  wire [(5'h15):(1'h0)] wire427;
  reg signed [(3'h6):(1'h0)] reg426 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg425 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg424 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg423 = (1'h0);
  reg [(3'h6):(1'h0)] reg422 = (1'h0);
  reg [(5'h12):(1'h0)] reg421 = (1'h0);
  reg [(4'h9):(1'h0)] reg420 = (1'h0);
  reg [(5'h14):(1'h0)] reg419 = (1'h0);
  reg [(4'ha):(1'h0)] reg418 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg417 = (1'h0);
  wire [(4'hc):(1'h0)] wire415;
  assign y = {wire430,
                 wire429,
                 wire428,
                 wire427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 wire415,
                 (1'h0)};
  module314 modinst416 (.wire318(wire310), .wire315(wire312), .wire317(wire311), .clk(clk), .wire316(wire313), .wire319((8'hb4)), .y(wire415));
  always
    @(posedge clk) begin
      reg417 <= (wire311[(2'h2):(1'h1)] ?
          $signed(wire415) : ({$signed(wire312),
                  $signed((wire310 ? wire313 : wire313))} ?
              ((~&(8'ha0)) << $signed(wire310)) : (~|wire313)));
      if (($signed((wire310[(1'h0):(1'h0)] && {$unsigned((8'haa))})) > $signed($unsigned({(~^wire310)}))))
        begin
          reg418 <= (7'h43);
          reg419 <= {$signed((-{(wire415 ? wire415 : wire313), reg418})),
              {(wire415 ? (^~reg417) : $signed((^~wire312)))}};
          reg420 <= (^~(($signed((^wire311)) ^~ {reg419}) <= (^wire313[(4'h9):(2'h2)])));
        end
      else
        begin
          if (reg417)
            begin
              reg418 <= ($signed($signed(wire415[(4'hc):(3'h6)])) | wire313);
              reg419 <= ((reg420 ^~ (^~((&(8'ha1)) + $signed(wire311)))) ?
                  $unsigned({reg417,
                      $unsigned(wire312)}) : $unsigned((reg418 + (wire312[(2'h2):(1'h1)] ^ $signed(wire313)))));
            end
          else
            begin
              reg418 <= $unsigned(wire415);
              reg419 <= wire311;
              reg420 <= $signed((~$unsigned(($unsigned(wire310) & $signed(wire415)))));
            end
          reg421 <= reg417[(3'h5):(3'h5)];
          reg422 <= {($signed(((~|reg418) ?
                  $unsigned((8'hb0)) : (wire311 ?
                      wire313 : wire312))) ~^ (reg421[(5'h10):(2'h2)] ~^ (^$signed(reg417)))),
              {(!(~^((8'hb4) ? reg419 : reg420)))}};
          if (reg418[(2'h2):(1'h0)])
            begin
              reg423 <= (8'ha8);
              reg424 <= reg418[(4'h8):(3'h4)];
            end
          else
            begin
              reg423 <= reg424;
            end
          reg425 <= {wire313, (wire311 ^ $signed((&reg424)))};
        end
      reg426 <= $unsigned(wire415[(4'hb):(4'h9)]);
    end
  assign wire427 = $signed(reg424);
  assign wire428 = $signed($signed(reg420[(3'h4):(2'h2)]));
  assign wire429 = $signed(((-$unsigned(wire313)) ?
                       $unsigned(((~&wire415) ^ reg417[(3'h7):(2'h2)])) : ({(+wire428),
                               wire428[(1'h0):(1'h0)]} ?
                           wire313 : reg420[(4'h9):(4'h9)])));
  assign wire430 = (wire428[(4'h8):(2'h3)] ^ wire313[(5'h13):(5'h11)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module19  (y, clk, wire20, wire21, wire22, wire23);
  output wire [(32'h417):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire20;
  input wire [(4'hf):(1'h0)] wire21;
  input wire [(5'h13):(1'h0)] wire22;
  input wire signed [(3'h6):(1'h0)] wire23;
  reg signed [(3'h5):(1'h0)] reg295 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg294 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg293 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire291;
  wire [(4'hb):(1'h0)] wire217;
  wire signed [(5'h11):(1'h0)] wire216;
  wire signed [(2'h3):(1'h0)] wire215;
  wire [(2'h3):(1'h0)] wire214;
  wire signed [(4'h8):(1'h0)] wire213;
  wire [(3'h4):(1'h0)] wire212;
  wire signed [(5'h14):(1'h0)] wire211;
  wire [(2'h3):(1'h0)] wire210;
  wire [(5'h12):(1'h0)] wire209;
  wire signed [(4'h9):(1'h0)] wire208;
  reg [(4'hb):(1'h0)] reg207 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg206 = (1'h0);
  reg [(3'h5):(1'h0)] reg205 = (1'h0);
  reg [(5'h13):(1'h0)] reg204 = (1'h0);
  reg [(3'h5):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg202 = (1'h0);
  reg [(2'h2):(1'h0)] reg201 = (1'h0);
  reg [(2'h2):(1'h0)] reg200 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire199;
  wire [(4'hd):(1'h0)] wire198;
  reg signed [(4'hc):(1'h0)] reg197 = (1'h0);
  reg [(3'h6):(1'h0)] reg196 = (1'h0);
  reg [(4'hf):(1'h0)] reg195 = (1'h0);
  reg [(4'hf):(1'h0)] reg194 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg24 = (1'h0);
  reg [(3'h4):(1'h0)] reg25 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg26 = (1'h0);
  reg [(3'h7):(1'h0)] reg27 = (1'h0);
  reg [(5'h15):(1'h0)] reg28 = (1'h0);
  reg [(4'h8):(1'h0)] reg29 = (1'h0);
  reg [(5'h15):(1'h0)] reg30 = (1'h0);
  reg [(4'hf):(1'h0)] reg31 = (1'h0);
  reg [(4'hf):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg33 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg34 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg35 = (1'h0);
  reg [(5'h10):(1'h0)] reg36 = (1'h0);
  reg [(4'hf):(1'h0)] reg37 = (1'h0);
  reg [(5'h15):(1'h0)] reg38 = (1'h0);
  reg [(4'he):(1'h0)] reg39 = (1'h0);
  reg [(4'h9):(1'h0)] reg40 = (1'h0);
  reg [(5'h14):(1'h0)] reg41 = (1'h0);
  reg [(5'h10):(1'h0)] reg42 = (1'h0);
  reg [(5'h13):(1'h0)] reg43 = (1'h0);
  reg [(5'h11):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg46 = (1'h0);
  reg signed [(4'he):(1'h0)] reg47 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg48 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg49 = (1'h0);
  reg [(5'h12):(1'h0)] reg50 = (1'h0);
  reg [(5'h12):(1'h0)] reg51 = (1'h0);
  reg [(5'h12):(1'h0)] reg52 = (1'h0);
  reg [(4'hc):(1'h0)] reg53 = (1'h0);
  wire [(5'h10):(1'h0)] wire54;
  wire [(4'h9):(1'h0)] wire55;
  reg signed [(4'h9):(1'h0)] reg56 = (1'h0);
  reg [(2'h2):(1'h0)] reg57 = (1'h0);
  reg [(5'h15):(1'h0)] reg58 = (1'h0);
  reg [(5'h13):(1'h0)] reg59 = (1'h0);
  reg [(5'h13):(1'h0)] reg60 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg61 = (1'h0);
  reg [(5'h12):(1'h0)] reg62 = (1'h0);
  reg [(4'h9):(1'h0)] reg63 = (1'h0);
  reg signed [(4'he):(1'h0)] reg64 = (1'h0);
  reg [(5'h15):(1'h0)] reg65 = (1'h0);
  reg [(5'h15):(1'h0)] reg66 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg67 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg68 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg69 = (1'h0);
  reg [(2'h3):(1'h0)] reg70 = (1'h0);
  reg [(3'h4):(1'h0)] reg71 = (1'h0);
  reg [(4'ha):(1'h0)] reg72 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg73 = (1'h0);
  reg [(4'ha):(1'h0)] reg74 = (1'h0);
  reg [(4'hb):(1'h0)] reg75 = (1'h0);
  reg [(4'ha):(1'h0)] reg76 = (1'h0);
  wire [(3'h7):(1'h0)] wire77;
  wire signed [(5'h11):(1'h0)] wire78;
  wire [(3'h4):(1'h0)] wire192;
  assign y = {reg295,
                 reg294,
                 reg293,
                 wire291,
                 wire217,
                 wire216,
                 wire215,
                 wire214,
                 wire213,
                 wire212,
                 wire211,
                 wire210,
                 wire209,
                 wire208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 wire199,
                 wire198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 reg28,
                 reg29,
                 reg30,
                 reg31,
                 reg32,
                 reg33,
                 reg34,
                 reg35,
                 reg36,
                 reg37,
                 reg38,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 reg44,
                 reg45,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 reg50,
                 reg51,
                 reg52,
                 reg53,
                 wire54,
                 wire55,
                 reg56,
                 reg57,
                 reg58,
                 reg59,
                 reg60,
                 reg61,
                 reg62,
                 reg63,
                 reg64,
                 reg65,
                 reg66,
                 reg67,
                 reg68,
                 reg69,
                 reg70,
                 reg71,
                 reg72,
                 reg73,
                 reg74,
                 reg75,
                 reg76,
                 wire77,
                 wire78,
                 wire192,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((($unsigned((&(wire23 + wire20))) ?
          (((!wire20) ? $unsigned(wire23) : wire20) ?
              ({(7'h42), wire20} ?
                  wire23[(1'h0):(1'h0)] : wire21[(2'h2):(2'h2)]) : wire20[(4'ha):(2'h3)]) : $unsigned(($unsigned(wire21) ?
              (-wire21) : ((8'ha7) ?
                  wire21 : wire23)))) || $signed({(wire20[(3'h7):(1'h0)] ?
              $signed(wire22) : {wire20}),
          (-(wire20 ? wire21 : (8'hb4)))})))
        begin
          if ($signed(wire21))
            begin
              reg24 <= ((|wire21[(4'h8):(2'h3)]) ?
                  $signed((8'ha8)) : $signed($unsigned($unsigned((-(8'hb8))))));
              reg25 <= (~&$signed(((~|wire23) <<< $signed((~^wire23)))));
              reg26 <= $signed($signed((wire22 ?
                  {reg24[(4'hd):(4'hc)]} : {$signed(wire22)})));
              reg27 <= (8'h9e);
              reg28 <= wire23[(2'h2):(1'h1)];
            end
          else
            begin
              reg24 <= $unsigned($signed($signed(($signed(wire22) * reg28))));
              reg25 <= $unsigned($unsigned({$unsigned($signed(reg27))}));
            end
          reg29 <= (8'hb4);
          reg30 <= {{(^((|(8'hb7)) ? (!reg29) : $signed(wire21))),
                  (!reg29[(2'h3):(1'h0)])},
              (^(8'h9d))};
          if ((wire20[(3'h4):(2'h3)] ?
              $signed(reg28[(4'hf):(4'hd)]) : $unsigned((($signed(reg26) & (wire20 ?
                      reg30 : wire23)) ?
                  reg24 : $signed(reg25)))))
            begin
              reg31 <= (~^(($signed({(7'h44)}) || reg24) && $unsigned(reg26[(1'h0):(1'h0)])));
              reg32 <= (-reg29[(3'h6):(3'h6)]);
              reg33 <= ({{wire20, $unsigned((|(8'hba)))}} ?
                  (reg28[(4'hd):(1'h0)] ?
                      wire20 : (~&$signed((|reg24)))) : (-$signed(reg25)));
            end
          else
            begin
              reg31 <= (wire20 ?
                  reg26 : $unsigned($unsigned(reg32[(4'hb):(3'h6)])));
              reg32 <= (-(8'hab));
              reg33 <= reg30[(2'h2):(2'h2)];
            end
          reg34 <= reg28[(5'h11):(2'h2)];
        end
      else
        begin
          if ($unsigned($signed($signed(reg24[(5'h12):(3'h5)]))))
            begin
              reg24 <= reg24[(4'h8):(3'h7)];
              reg25 <= reg26[(1'h1):(1'h1)];
              reg26 <= wire21;
              reg27 <= (((|$signed({(8'ha6), reg24})) ?
                  (&reg24[(5'h10):(3'h4)]) : ((8'hba) ?
                      reg25[(2'h3):(1'h1)] : reg28[(1'h0):(1'h0)])) | ($unsigned(wire23) ?
                  reg26 : $signed((wire21 || wire20[(3'h4):(2'h3)]))));
              reg28 <= {($signed($signed($unsigned(reg32))) ?
                      reg32 : ($signed({wire21, wire23}) ?
                          {(reg25 ? wire23 : reg26),
                              $signed(reg32)} : wire21[(3'h4):(2'h3)]))};
            end
          else
            begin
              reg24 <= ($unsigned({(!(reg30 ? reg28 : reg27)),
                  reg33[(4'hc):(1'h1)]}) * ((+{$unsigned(reg29)}) * {reg34[(4'h8):(3'h4)]}));
              reg25 <= $signed({($unsigned($unsigned(reg33)) ^ $unsigned(reg27[(3'h4):(3'h4)])),
                  (+wire23[(1'h0):(1'h0)])});
            end
          reg29 <= (reg32[(4'hf):(4'hf)] && (~^(8'hb8)));
          reg30 <= reg27;
        end
      if ((~|wire23))
        begin
          reg35 <= $unsigned(reg29[(3'h6):(1'h1)]);
          reg36 <= ($signed({reg27[(3'h7):(2'h3)], (8'ha0)}) ?
              wire22 : (~^reg33));
          reg37 <= wire20;
          reg38 <= (|{$unsigned({(wire21 ? reg24 : reg24), $signed(reg30)})});
        end
      else
        begin
          if (reg29[(1'h0):(1'h0)])
            begin
              reg35 <= $unsigned($signed($signed($signed($signed(reg36)))));
              reg36 <= ((wire22 ?
                  $unsigned(reg27) : (reg28 >= wire20[(3'h4):(2'h2)])) + $signed(({(!(8'ha7)),
                  $unsigned((8'ha5))} + wire20[(3'h5):(1'h0)])));
              reg37 <= ($unsigned($unsigned(reg33)) >>> $unsigned($signed(((^(8'hb3)) * $unsigned(reg34)))));
              reg38 <= $unsigned(reg25);
              reg39 <= {($signed(reg33[(1'h1):(1'h1)]) ?
                      $signed($unsigned({(8'h9c), reg27})) : wire23),
                  reg26};
            end
          else
            begin
              reg35 <= reg31;
              reg36 <= reg30[(2'h3):(2'h2)];
              reg37 <= $unsigned($unsigned(($unsigned(reg37) <<< (reg28 >> {reg27}))));
            end
          if ({$signed($signed($signed((reg28 ? reg25 : reg25)))),
              wire21[(1'h0):(1'h0)]})
            begin
              reg40 <= ((~^(~$unsigned(reg34))) ?
                  wire21[(3'h7):(3'h4)] : wire20);
              reg41 <= {reg28,
                  {($unsigned((reg24 <<< reg40)) ? (^~(!wire21)) : wire23)}};
              reg42 <= $signed(reg34);
              reg43 <= (!(reg29 < {$signed($signed(reg41)), $signed({reg28})}));
              reg44 <= (&$signed($signed($signed(reg37[(4'ha):(3'h5)]))));
            end
          else
            begin
              reg40 <= (~|wire21);
              reg41 <= ($signed({($signed((8'ha0)) ^~ $unsigned(reg40))}) == reg41);
              reg42 <= ({(~|{$unsigned(reg30)}),
                      ($signed($unsigned(reg32)) & {reg36, $signed(reg42)})} ?
                  $unsigned($unsigned(({reg32, (8'hb0)} ?
                      $unsigned(reg37) : wire23[(3'h5):(1'h0)]))) : $signed((!$unsigned((reg33 & reg32)))));
              reg43 <= (reg42 ? reg43 : wire20[(4'h9):(4'h9)]);
              reg44 <= (^$unsigned((($signed((8'haa)) != reg38[(4'ha):(3'h6)]) >= (8'ha1))));
            end
          if ((~($unsigned((wire23 ?
              (^~(8'h9d)) : reg35[(1'h0):(1'h0)])) & {reg32[(3'h4):(1'h1)]})))
            begin
              reg45 <= reg25;
              reg46 <= reg28;
              reg47 <= $unsigned(reg25);
              reg48 <= reg38;
              reg49 <= ({(((&reg37) ?
                          $unsigned((8'hb9)) : reg35[(3'h4):(1'h0)]) ?
                      $signed((-reg42)) : ({reg33} ?
                          ((8'hbb) ? reg44 : (8'hb2)) : (reg45 < reg35))),
                  (reg34 ?
                      ((reg26 < reg33) ?
                          reg25 : (~^wire21)) : reg48)} - (&(reg46[(5'h13):(3'h5)] ?
                  $signed((reg43 - reg25)) : $signed({wire22, reg24}))));
            end
          else
            begin
              reg45 <= (~&{($unsigned((reg44 < reg29)) || (~&(-wire23))),
                  {$signed($unsigned(reg24)), $unsigned(reg49)}});
              reg46 <= (reg26[(2'h2):(1'h0)] ?
                  $signed(reg43) : ({(wire23[(3'h5):(1'h1)] ?
                              wire20[(1'h1):(1'h1)] : $unsigned(reg33)),
                          ((reg27 >= (8'hab)) & reg42)} ?
                      ((~&{reg45, (8'hba)}) < ({(8'hb3)} && (reg49 ?
                          reg29 : reg30))) : $unsigned((~&(reg40 ^ reg35)))));
              reg47 <= $signed($signed(((reg45 ?
                      $signed(reg38) : {reg24, (8'ha7)}) ?
                  reg31 : reg36[(3'h4):(2'h3)])));
            end
          reg50 <= (&(reg34[(1'h0):(1'h0)] ?
              (~&$signed((reg32 ?
                  reg43 : reg25))) : $unsigned($unsigned($unsigned(reg37)))));
          if ((^~reg46[(3'h7):(2'h3)]))
            begin
              reg51 <= {$unsigned($unsigned(reg36[(3'h5):(1'h1)])),
                  (+(-((reg27 ? reg25 : (8'hb7)) < {wire23, reg30})))};
              reg52 <= $signed(reg24[(2'h2):(1'h0)]);
            end
          else
            begin
              reg51 <= (($signed((reg27[(1'h0):(1'h0)] ?
                          (&reg51) : wire20[(4'h8):(3'h5)])) ?
                      (wire23[(1'h1):(1'h1)] ?
                          ($unsigned(reg37) ?
                              (reg52 ?
                                  reg27 : reg40) : (^~reg29)) : reg26[(2'h3):(1'h1)]) : $signed(wire22[(4'hc):(2'h3)])) ?
                  ((($unsigned(reg30) ?
                      $signed(reg39) : reg26[(3'h5):(3'h4)]) | {(reg43 ?
                          reg36 : reg52)}) + $unsigned($unsigned((reg40 < (8'hbb))))) : {{reg24[(1'h1):(1'h1)],
                          (~&reg35)}});
              reg52 <= $unsigned({(!$unsigned((reg48 << reg29))),
                  (reg29 ?
                      $signed(reg44) : ((wire20 ?
                          reg30 : reg26) >> (^reg33)))});
              reg53 <= ((reg31[(4'ha):(4'h9)] ?
                      (reg49[(1'h0):(1'h0)] ?
                          $signed(reg27[(1'h1):(1'h0)]) : $signed((reg31 ?
                              reg42 : reg28))) : (^reg43[(4'ha):(2'h2)])) ?
                  reg52 : (~reg39));
            end
        end
    end
  assign wire54 = {((8'hbb) >> $signed((~|{reg38})))};
  assign wire55 = reg49[(3'h4):(1'h0)];
  always
    @(posedge clk) begin
      if ((8'h9c))
        begin
          if (({$unsigned({reg36[(3'h6):(2'h2)], $unsigned(reg25)}),
                  $unsigned((~{reg52, (7'h41)}))} ?
              $signed($signed($signed((wire20 ?
                  reg51 : reg40)))) : (wire22[(2'h2):(1'h1)] & reg35[(3'h4):(2'h3)])))
            begin
              reg56 <= (((~(~wire20)) * $signed($signed((^reg24)))) >> $unsigned($unsigned(reg49[(4'hc):(2'h3)])));
              reg57 <= reg41[(4'h8):(2'h3)];
              reg58 <= reg56;
              reg59 <= ($signed((+reg44)) << reg45);
            end
          else
            begin
              reg56 <= $signed((reg56[(4'h9):(1'h0)] && $unsigned(((~^reg25) ?
                  (reg40 || (8'hb7)) : (reg28 ? reg52 : wire20)))));
              reg57 <= reg50;
              reg58 <= reg30[(5'h12):(4'he)];
              reg59 <= reg25;
            end
          if ((^~$signed(reg39[(3'h7):(1'h0)])))
            begin
              reg60 <= ($signed({{((8'h9c) ? (8'hb3) : (7'h42)),
                      $unsigned(wire21)}}) != ($unsigned(((wire54 || reg40) ?
                      (wire22 ? (8'hb1) : reg27) : {reg40})) ?
                  (((~&reg58) >>> (reg36 ?
                      reg51 : reg45)) <= $unsigned($signed((8'ha7)))) : $unsigned($unsigned({reg53}))));
              reg61 <= reg30[(4'ha):(2'h2)];
              reg62 <= reg45;
              reg63 <= $signed((~^(((8'hb1) ? (~^reg59) : (+reg30)) ?
                  (^reg39) : ($unsigned(reg57) ? {wire23} : $signed(reg61)))));
              reg64 <= $signed(($signed($signed((!reg31))) ?
                  ($unsigned($signed(wire22)) ^ ((-reg44) & (reg36 || wire20))) : $unsigned($signed($signed((8'hac))))));
            end
          else
            begin
              reg60 <= (^(~&$signed(reg51[(4'hf):(3'h4)])));
              reg61 <= (^reg53);
              reg62 <= $signed($signed(reg27[(2'h3):(1'h1)]));
              reg63 <= (((|reg35[(4'hb):(3'h5)]) * $unsigned(($signed(reg31) ?
                  (reg62 == reg32) : (reg37 ?
                      reg36 : reg45)))) | reg50[(1'h1):(1'h1)]);
            end
          if (reg25[(1'h0):(1'h0)])
            begin
              reg65 <= (($unsigned($unsigned(reg34[(3'h4):(2'h3)])) << $unsigned((~$signed(reg25)))) && reg24);
              reg66 <= (!(+(((wire23 ? reg27 : reg58) ?
                      $unsigned(reg52) : reg40[(1'h1):(1'h1)]) ?
                  $unsigned(reg46) : $signed((reg62 ? reg45 : wire55)))));
              reg67 <= {((wire22[(4'ha):(3'h5)] >> (&reg47[(1'h1):(1'h1)])) ?
                      $signed((~(wire20 == reg37))) : (&(^(wire54 || wire23))))};
              reg68 <= ((((~&(8'hb6)) != (^~(reg60 ~^ reg58))) ?
                      (wire54 ?
                          $unsigned((&reg31)) : (~&reg49)) : reg65[(5'h12):(5'h11)]) ?
                  (($signed((wire23 ^ wire23)) ? (!(&reg42)) : reg30) ?
                      $unsigned(reg44) : reg31[(4'hf):(4'he)]) : ({$signed(reg52[(5'h12):(3'h5)]),
                      ($signed(reg38) ?
                          reg59[(4'he):(4'h8)] : ((8'hab) ?
                              reg29 : wire54))} * {({reg50} ?
                          (|reg42) : reg30)}));
            end
          else
            begin
              reg65 <= (((~&{(^~reg52)}) ?
                  $signed((!(reg30 >> (8'hb3)))) : reg35) >>> $signed((wire54[(4'hd):(3'h7)] ?
                  (8'hab) : reg62)));
              reg66 <= ($unsigned(({(-reg28), $unsigned(reg53)} ?
                  wire20 : ((reg61 ?
                      wire20 : reg26) >> reg45[(2'h3):(2'h2)]))) + ($unsigned(reg68) >>> ($signed((&reg33)) ^~ ((reg41 >= reg62) ?
                  wire54[(4'hb):(3'h7)] : (reg25 ? wire20 : reg47)))));
              reg67 <= reg63[(1'h1):(1'h0)];
              reg68 <= ((^{reg60, reg37}) ^ reg38);
            end
          reg69 <= reg36;
        end
      else
        begin
          if ((8'hbc))
            begin
              reg56 <= (reg29[(2'h2):(2'h2)] * {(-$unsigned($unsigned(reg48)))});
            end
          else
            begin
              reg56 <= {(reg26 & wire23), (8'ha1)};
            end
          if (reg59)
            begin
              reg57 <= (^~wire55[(1'h0):(1'h0)]);
              reg58 <= (((($unsigned(reg67) != (reg59 >= wire22)) <<< ($signed(reg24) ?
                          $signed(reg24) : $signed(reg37))) ?
                      reg35[(3'h7):(1'h1)] : $unsigned(reg60)) ?
                  (reg29 == $signed($signed((reg67 ?
                      reg47 : reg33)))) : $unsigned((~&(~(reg66 ?
                      wire23 : reg41)))));
            end
          else
            begin
              reg57 <= ((8'hb8) ?
                  {(~|(~&(&reg42))),
                      ({$signed(reg53), $unsigned(reg52)} ?
                          reg60 : (!(^~reg36)))} : (reg27[(3'h5):(3'h5)] ?
                      $unsigned(reg42) : reg60));
              reg58 <= ({(+$signed((^reg62)))} ?
                  (($signed($signed(reg27)) * {$unsigned(reg42),
                      (wire20 ?
                          reg52 : reg27)}) || reg59[(4'hb):(2'h2)]) : reg57[(2'h2):(2'h2)]);
              reg59 <= (~^reg50[(3'h6):(3'h5)]);
              reg60 <= reg46[(5'h15):(1'h1)];
            end
        end
      if (reg56[(2'h3):(2'h2)])
        begin
          reg70 <= reg31;
        end
      else
        begin
          reg70 <= (&(~|$unsigned({reg50[(4'hd):(2'h3)], (~^reg40)})));
        end
      reg71 <= reg46[(5'h10):(3'h5)];
      if ($unsigned(((^reg48) <= $unsigned(reg41[(3'h6):(3'h5)]))))
        begin
          reg72 <= ($signed(($signed((&reg38)) ?
                  $signed((reg71 ? wire21 : (8'hb6))) : ($unsigned(reg34) ?
                      $unsigned(reg42) : (reg41 ? reg45 : reg27)))) ?
              (!(|$signed({reg25}))) : (($signed(((8'ha1) ?
                      reg28 : reg29)) >> reg41[(5'h12):(4'hf)]) ?
                  $unsigned((reg69[(3'h7):(3'h5)] && ((8'hb1) ?
                      reg41 : reg31))) : (({reg67} >= (!reg25)) ?
                      ($signed(reg27) ?
                          (reg65 ?
                              reg47 : reg64) : (reg43 >>> reg39)) : (8'hb0))));
          reg73 <= (wire21 >> ($signed(({(8'hb5), reg42} > {reg53})) ?
              {reg26[(3'h5):(1'h1)],
                  ((reg68 ? reg36 : reg48) != (8'hb4))} : (reg69 ?
                  $unsigned($signed(reg64)) : (8'hb2))));
        end
      else
        begin
          reg72 <= ($signed({(reg28[(4'hd):(1'h0)] ? $signed(reg72) : (~reg72)),
                  reg56[(1'h0):(1'h0)]}) ?
              reg31[(4'hc):(4'h8)] : reg58[(3'h4):(3'h4)]);
          if ({(+$unsigned((~|reg40))),
              ((((+reg57) ^ (reg24 > (8'haa))) ^~ (reg44[(3'h4):(1'h0)] ?
                  $signed(wire54) : ((8'ha8) & wire23))) << {$signed($unsigned(reg35)),
                  $signed($signed(wire21))})})
            begin
              reg73 <= (wire22[(1'h0):(1'h0)] ~^ {(((reg37 ~^ reg52) ?
                      (&reg68) : $signed(reg38)) - ((+reg57) > (^reg26)))});
              reg74 <= reg29[(3'h7):(1'h1)];
              reg75 <= $signed($signed(((~&reg50[(4'hc):(3'h5)]) * reg71[(1'h1):(1'h0)])));
            end
          else
            begin
              reg73 <= reg67[(4'h8):(3'h6)];
              reg74 <= (~((^~reg31) & reg41));
            end
          reg76 <= ((reg75[(2'h2):(1'h0)] >>> {reg41[(5'h13):(4'ha)]}) ?
              (^~$signed((+$unsigned((7'h43))))) : reg43);
        end
    end
  assign wire77 = (~(((8'hb0) ?
                          (+(reg32 > (8'hba))) : $signed($signed((8'ha3)))) ?
                      (8'hb9) : (!$unsigned({reg61, reg69}))));
  assign wire78 = $unsigned((($signed({reg26}) >>> ((reg26 < reg36) == $signed(reg71))) << $unsigned(reg52)));
  module79 modinst193 (.y(wire192), .wire82(reg40), .clk(clk), .wire81(wire21), .wire80(reg62), .wire83(reg76), .wire84(reg67));
  always
    @(posedge clk) begin
      if ($unsigned((~|reg35)))
        begin
          if (reg46[(5'h10):(2'h3)])
            begin
              reg194 <= (reg36[(3'h7):(3'h5)] ?
                  $unsigned((|(~^$signed(reg25)))) : wire22);
            end
          else
            begin
              reg194 <= $signed((!$signed(($signed(reg33) ?
                  (8'hb3) : (wire21 >> reg33)))));
              reg195 <= wire20[(4'h9):(3'h5)];
              reg196 <= (+($signed($unsigned((~&(7'h43)))) == (~&reg25[(1'h1):(1'h1)])));
              reg197 <= reg64;
            end
        end
      else
        begin
          reg194 <= $signed(reg195);
        end
    end
  assign wire198 = $unsigned((reg59 >>> $unsigned((8'hbf))));
  assign wire199 = reg56[(2'h3):(2'h2)];
  always
    @(posedge clk) begin
      if ($unsigned(((($unsigned(wire199) ?
              $signed((8'hbb)) : reg49) <<< reg37[(1'h1):(1'h1)]) ?
          ((!$signed(reg64)) ?
              reg71[(1'h0):(1'h0)] : $signed(reg65[(5'h11):(3'h7)])) : (~reg40[(2'h2):(2'h2)]))))
        begin
          if (reg32)
            begin
              reg200 <= reg59[(5'h12):(1'h0)];
              reg201 <= (((~reg52) ~^ {$unsigned((^~(8'ha5)))}) ?
                  wire77 : $signed((~&(8'hbc))));
            end
          else
            begin
              reg200 <= $signed({(-(~$signed(reg46))), (|(-reg50))});
              reg201 <= ((^({(reg36 ? reg201 : wire199),
                      reg50} & reg29[(3'h5):(2'h3)])) ?
                  reg58[(4'hd):(1'h0)] : (reg32 ?
                      $unsigned(($unsigned(reg72) ?
                          (~reg44) : $signed(reg39))) : (|reg26)));
              reg202 <= {(7'h44), reg52};
              reg203 <= $unsigned($unsigned(reg32));
            end
        end
      else
        begin
          reg200 <= wire23[(3'h4):(1'h0)];
          reg201 <= {$signed(reg203[(1'h1):(1'h0)]),
              {$unsigned({reg67[(4'hb):(3'h5)], (reg25 ? reg51 : reg27)}),
                  {$unsigned(reg45), (wire198 >= (&reg195))}}};
          if (reg66)
            begin
              reg202 <= {(wire198 & ((~^(reg62 ?
                      reg67 : reg197)) & ((^~reg52) >> {reg47, reg52}))),
                  reg69};
              reg203 <= (-wire78[(4'h8):(2'h2)]);
            end
          else
            begin
              reg202 <= ($unsigned($unsigned(reg72[(3'h6):(2'h2)])) ?
                  $signed((~&(^~(reg47 | (8'ha0))))) : ((^{((8'haa) ?
                              reg59 : reg52)}) ?
                      {reg58} : $signed($unsigned($unsigned(reg195)))));
            end
        end
      reg204 <= (wire22[(4'ha):(3'h6)] * $unsigned(($unsigned(reg47[(3'h6):(3'h6)]) ?
          reg202[(2'h2):(2'h2)] : reg69[(1'h0):(1'h0)])));
      reg205 <= reg43;
      reg206 <= reg69;
      reg207 <= reg40;
    end
  assign wire208 = {reg70[(2'h2):(1'h0)],
                       ($unsigned(wire192[(1'h0):(1'h0)]) ?
                           $unsigned(($unsigned(reg70) ?
                               $unsigned(wire54) : wire21)) : (({(8'h9f),
                                   reg196} <= wire55[(2'h2):(2'h2)]) ?
                               ((wire199 != (7'h41)) >>> reg71[(1'h0):(1'h0)]) : wire20))};
  assign wire209 = reg34[(3'h4):(1'h1)];
  assign wire210 = $unsigned((($signed(reg195[(4'hd):(4'hc)]) ?
                       (reg67 == $unsigned((8'ha9))) : reg41) <<< reg206));
  assign wire211 = $signed($unsigned({((reg45 <= reg28) != {(8'hb9)}),
                       reg33[(2'h2):(1'h0)]}));
  assign wire212 = reg204;
  assign wire213 = (&((&((reg197 ? reg51 : reg25) || (~^reg203))) ~^ reg61));
  assign wire214 = (((wire213 ?
                           reg42[(2'h3):(1'h1)] : $unsigned($signed(reg35))) ?
                       ((^~reg63[(1'h0):(1'h0)]) ~^ ((~(8'hb3)) ~^ ((8'hbd) ?
                           (8'hb8) : reg42))) : (^$signed({reg196,
                           reg196}))) & ($signed((+(wire213 + reg200))) != $signed({(reg59 >= reg74),
                       (wire192 ? reg203 : reg207)})));
  assign wire215 = wire77;
  assign wire216 = {(^(reg66 ? {reg69[(4'h8):(3'h6)], reg69} : reg197))};
  assign wire217 = $signed((7'h40));
  module218 modinst292 (.wire220(reg60), .wire219(reg61), .clk(clk), .wire222(reg204), .wire221(wire22), .y(wire291));
  always
    @(posedge clk) begin
      reg293 <= $unsigned((($signed($unsigned(wire209)) ^ $unsigned((reg50 >>> reg200))) >> (~|$signed((~reg25)))));
      reg294 <= ($unsigned(reg68) ?
          reg205[(3'h5):(1'h1)] : (reg34 ?
              ((&(reg45 & wire77)) ?
                  (((7'h42) > reg62) ?
                      (reg74 ?
                          reg197 : reg202) : (8'hb0)) : $unsigned(reg194)) : reg201[(1'h0):(1'h0)]));
      reg295 <= (~{(((&wire55) ? (reg201 ? (8'hb3) : reg65) : $signed(reg66)) ?
              (!$unsigned((8'hbe))) : $signed(((8'ha0) ? reg43 : wire20)))});
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module218
#( parameter param289 = (+((^(!((8'h9c) > (8'ha9)))) << ((((8'hbb) ^~ (8'hb8)) ? {(8'hba), (8'h9d)} : ((8'ha5) ? (8'ha7) : (8'ha6))) ? (((8'hbb) <<< (8'h9e)) ^~ ((8'h9c) ? (8'hb6) : (8'h9e))) : ((8'ha8) ? (~&(8'hba)) : ((8'ha4) ? (8'hb5) : (8'hab))))))
, parameter param290 = param289 )
(y, clk, wire219, wire220, wire221, wire222);
  output wire [(32'h10f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire219;
  input wire signed [(5'h13):(1'h0)] wire220;
  input wire [(5'h12):(1'h0)] wire221;
  input wire [(5'h13):(1'h0)] wire222;
  wire signed [(5'h10):(1'h0)] wire288;
  wire [(2'h3):(1'h0)] wire287;
  wire [(4'ha):(1'h0)] wire286;
  wire [(4'hc):(1'h0)] wire284;
  reg signed [(5'h13):(1'h0)] reg272 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg271 = (1'h0);
  reg signed [(4'he):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg269 = (1'h0);
  reg [(3'h7):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg267 = (1'h0);
  reg [(5'h10):(1'h0)] reg266 = (1'h0);
  wire [(5'h11):(1'h0)] wire265;
  wire [(3'h7):(1'h0)] wire264;
  wire signed [(4'h9):(1'h0)] wire238;
  wire [(5'h15):(1'h0)] wire240;
  reg signed [(4'ha):(1'h0)] reg241 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg242 = (1'h0);
  reg [(4'hb):(1'h0)] reg243 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire244;
  wire [(3'h5):(1'h0)] wire245;
  wire signed [(5'h14):(1'h0)] wire262;
  assign y = {wire288,
                 wire287,
                 wire286,
                 wire284,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 wire265,
                 wire264,
                 wire238,
                 wire240,
                 reg241,
                 reg242,
                 reg243,
                 wire244,
                 wire245,
                 wire262,
                 (1'h0)};
  module223 modinst239 (wire238, clk, wire220, wire219, wire222, wire221);
  assign wire240 = wire222;
  always
    @(posedge clk) begin
      reg241 <= wire221[(5'h11):(4'h8)];
      reg242 <= $signed((^$signed(((reg241 ? wire221 : reg241) ?
          (8'hae) : $unsigned(wire240)))));
      reg243 <= (~^(wire219[(1'h1):(1'h1)] ?
          (^{wire240, (wire222 - reg242)}) : (({(8'hb0)} ?
              $signed((8'hb2)) : (wire219 || (8'hb0))) && $unsigned(wire219[(4'h9):(2'h3)]))));
    end
  assign wire244 = wire222[(4'h9):(3'h4)];
  assign wire245 = (wire222 ~^ (wire220[(3'h4):(1'h0)] ?
                       $signed($unsigned({wire244,
                           (8'hb3)})) : $unsigned(wire238[(4'h9):(4'h9)])));
  module246 modinst263 (.clk(clk), .wire249(wire219), .wire247(wire220), .wire250(wire221), .wire251(wire240), .y(wire262), .wire248(wire245));
  assign wire264 = wire221[(4'ha):(3'h7)];
  assign wire265 = (-$signed($unsigned(($unsigned(wire262) > (wire238 | (8'hbb))))));
  always
    @(posedge clk) begin
      reg266 <= (&$signed((wire264[(2'h3):(2'h3)] | ($signed(wire264) ?
          wire219 : (wire221 < wire238)))));
      reg267 <= $signed(($signed($signed($signed(wire264))) ?
          $unsigned((reg266[(4'hd):(3'h6)] + (8'h9e))) : (8'h9d)));
      if ($unsigned(((reg266 ?
          $signed(wire220[(2'h3):(1'h1)]) : ((~&wire244) & (7'h44))) << $signed((+$signed(wire219))))))
        begin
          reg268 <= ($signed($signed($unsigned((reg243 ?
              reg267 : wire245)))) && ({(wire262 ? (^~wire240) : wire221),
              wire240[(3'h7):(1'h1)]} < ($signed(reg266) ?
              ((wire264 ?
                  wire265 : wire244) ^ (wire222 <= wire220)) : (&(~^wire262)))));
          reg269 <= (+({$unsigned(reg242[(3'h4):(2'h3)])} ?
              (reg268 <<< ((wire244 ~^ reg242) ?
                  (wire240 ^ reg267) : {wire265,
                      wire219})) : (~&((wire264 ~^ wire222) <= (reg243 ?
                  wire240 : reg243)))));
          reg270 <= reg242;
          reg271 <= ((reg269[(5'h14):(4'ha)] & $unsigned((-reg243[(3'h6):(3'h5)]))) ^~ (~^(8'ha7)));
        end
      else
        begin
          reg268 <= (($unsigned(($unsigned(reg241) ?
                  (reg242 ? wire265 : (8'hae)) : (reg242 | wire244))) ?
              $signed(reg267[(2'h3):(2'h3)]) : $unsigned(({(8'ha7),
                  reg271} ^ {wire222}))) <= {wire245[(3'h5):(3'h4)]});
          reg269 <= $signed((^~((8'had) >= (7'h42))));
          reg270 <= (reg269[(4'hb):(3'h7)] || $unsigned(reg268[(3'h6):(3'h4)]));
        end
      reg272 <= (+$unsigned($signed(reg270)));
    end
  module273 modinst285 (wire284, clk, reg241, wire244, wire265, wire240);
  assign wire286 = ($unsigned(wire240[(5'h13):(4'ha)]) ?
                       (($signed(reg269) ?
                           ($signed(wire264) ?
                               (wire238 ? reg269 : (8'hb6)) : (wire220 ?
                                   wire284 : (8'hbd))) : wire221[(4'h8):(4'h8)]) * $signed((+(reg242 == wire262)))) : (8'hb7));
  assign wire287 = (&((reg269[(1'h0):(1'h0)] < reg241[(1'h0):(1'h0)]) && (($signed(wire220) ?
                           ((8'ha0) <<< reg241) : wire245[(2'h3):(1'h1)]) ?
                       $signed(reg272[(3'h7):(3'h6)]) : $unsigned((!(7'h40))))));
  assign wire288 = (~$unsigned(wire220));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module79
#( parameter param191 = (({(!{(8'hbc)})} ? {((!(8'ha2)) ? (|(7'h43)) : (~^(8'hb4))), {((7'h40) ? (8'ha1) : (8'had))}} : ({(!(8'hba)), ((8'hb7) ? (8'hb8) : (8'ha3))} > (((8'ha3) + (8'hb4)) ? {(8'hb5), (8'ha6)} : ((8'ha6) >> (8'h9c))))) ~^ ((^(^~((8'h9c) * (8'ha4)))) ^ (({(8'hb4)} ? ((8'hae) <= (8'hbd)) : (!(8'ha2))) ? (~|((8'hbe) ? (7'h44) : (8'hb5))) : (((8'hab) | (8'hb5)) ? ((8'haf) << (7'h43)) : (+(7'h43)))))) )
(y, clk, wire80, wire81, wire82, wire83, wire84);
  output wire [(32'h165):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire80;
  input wire signed [(4'hf):(1'h0)] wire81;
  input wire signed [(4'h9):(1'h0)] wire82;
  input wire [(4'ha):(1'h0)] wire83;
  input wire signed [(5'h15):(1'h0)] wire84;
  wire signed [(4'hb):(1'h0)] wire190;
  wire signed [(4'he):(1'h0)] wire189;
  wire [(5'h12):(1'h0)] wire188;
  wire [(5'h11):(1'h0)] wire187;
  wire [(3'h4):(1'h0)] wire186;
  wire [(4'he):(1'h0)] wire85;
  wire [(3'h7):(1'h0)] wire86;
  wire [(5'h10):(1'h0)] wire87;
  reg signed [(4'hf):(1'h0)] reg88 = (1'h0);
  reg [(5'h15):(1'h0)] reg89 = (1'h0);
  reg [(4'ha):(1'h0)] reg90 = (1'h0);
  wire [(5'h13):(1'h0)] wire91;
  wire signed [(4'h9):(1'h0)] wire92;
  wire [(5'h13):(1'h0)] wire93;
  wire signed [(5'h12):(1'h0)] wire94;
  reg signed [(5'h11):(1'h0)] reg95 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg96 = (1'h0);
  wire [(5'h15):(1'h0)] wire97;
  wire signed [(2'h3):(1'h0)] wire98;
  wire signed [(5'h10):(1'h0)] wire99;
  reg [(4'he):(1'h0)] reg100 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg101 = (1'h0);
  reg [(4'hd):(1'h0)] reg102 = (1'h0);
  reg [(4'h9):(1'h0)] reg103 = (1'h0);
  wire [(4'h9):(1'h0)] wire104;
  wire signed [(3'h5):(1'h0)] wire144;
  wire [(2'h2):(1'h0)] wire184;
  assign y = {wire190,
                 wire189,
                 wire188,
                 wire187,
                 wire186,
                 wire85,
                 wire86,
                 wire87,
                 reg88,
                 reg89,
                 reg90,
                 wire91,
                 wire92,
                 wire93,
                 wire94,
                 reg95,
                 reg96,
                 wire97,
                 wire98,
                 wire99,
                 reg100,
                 reg101,
                 reg102,
                 reg103,
                 wire104,
                 wire144,
                 wire184,
                 (1'h0)};
  assign wire85 = (~|wire80);
  assign wire86 = $unsigned(wire83);
  assign wire87 = wire81[(4'h9):(4'h8)];
  always
    @(posedge clk) begin
      reg88 <= (~&wire87);
      reg89 <= $signed(wire86);
      reg90 <= (8'hb9);
    end
  assign wire91 = ($signed((8'hb6)) * ($signed($signed(wire80[(2'h2):(2'h2)])) ?
                      {(+reg89)} : (!reg89)));
  assign wire92 = {$unsigned(($unsigned({(8'hae),
                          wire81}) ^ ($signed((8'hba)) <<< ((8'hbc) ~^ reg90)))),
                      (((!wire82) < wire82) ~^ (^$unsigned(wire91[(3'h6):(1'h1)])))};
  assign wire93 = $signed(((((8'ha1) ^~ (+wire86)) ?
                      $signed((~&reg90)) : $unsigned(wire80[(1'h1):(1'h1)])) <= (($signed(wire82) * $signed(wire87)) ?
                      wire86[(2'h2):(1'h0)] : (!$signed((8'h9c))))));
  assign wire94 = (wire87 ?
                      (&$unsigned($signed((reg88 == wire91)))) : ((reg89 <<< $unsigned({wire83})) ?
                          (wire92 ?
                              wire81 : reg88[(2'h2):(1'h1)]) : ((^(^(7'h41))) <= reg88)));
  always
    @(posedge clk) begin
      reg95 <= ((!((wire92 ?
          (wire81 > (8'hb4)) : {wire86}) ^~ wire83[(4'h8):(3'h6)])) <<< wire84[(2'h2):(1'h0)]);
      reg96 <= wire87;
    end
  assign wire97 = $unsigned(($signed($signed($signed(reg90))) ?
                      ({(8'ha3), ((7'h42) | wire92)} ?
                          wire93 : $signed(wire81)) : {($signed((8'hb3)) ?
                              ((8'hb4) << wire92) : $signed(reg96))}));
  assign wire98 = ($unsigned($signed(wire92)) + wire83[(1'h1):(1'h1)]);
  assign wire99 = (~&wire85[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      reg100 <= ((~^(wire82[(2'h3):(1'h1)] >= $signed((^~wire91)))) - (wire86[(3'h5):(1'h1)] && reg90));
    end
  always
    @(posedge clk) begin
      reg101 <= wire94;
      reg102 <= (wire92[(1'h0):(1'h0)] <= (8'haa));
    end
  always
    @(posedge clk) begin
      reg103 <= wire86[(3'h7):(1'h1)];
    end
  assign wire104 = reg90[(4'h9):(2'h2)];
  module105 modinst145 (.wire109(wire82), .wire107(wire91), .wire108(wire93), .clk(clk), .y(wire144), .wire106(reg102));
  module146 modinst185 (.clk(clk), .wire148(wire97), .wire149(wire144), .wire150(wire84), .wire147(reg100), .y(wire184), .wire151(wire87));
  assign wire186 = reg88;
  assign wire187 = ((wire80[(2'h3):(2'h2)] ?
                           $unsigned(reg89[(5'h11):(4'hf)]) : (^~((wire87 ?
                                   reg89 : reg95) ?
                               $unsigned(reg88) : (~reg90)))) ?
                       $signed(($signed($signed(reg101)) ?
                           $unsigned(wire92[(4'h9):(1'h0)]) : $signed($unsigned(wire99)))) : ((^~(^~wire184[(1'h1):(1'h0)])) ^~ wire104[(2'h3):(1'h1)]));
  assign wire188 = $signed($unsigned(wire104));
  assign wire189 = (~&wire144[(2'h2):(1'h1)]);
  assign wire190 = {$signed(reg102)};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module146
#( parameter param182 = (|(({(&(8'hb1))} <<< (((8'hb9) ? (7'h40) : (7'h44)) ~^ (&(8'ha2)))) || {((+(8'ha2)) ? (~|(8'hbb)) : ((7'h43) == (8'ha5)))}))
, parameter param183 = ((~^{(^~param182), ((8'hb5) ? (~param182) : (param182 ? param182 : param182))}) || ((+(param182 || {(8'hb3)})) ^~ (((-param182) ? (~&param182) : (~^(8'hbc))) ? param182 : ((~|param182) ? (param182 ? param182 : (8'haf)) : (-param182))))) )
(y, clk, wire151, wire150, wire149, wire148, wire147);
  output wire [(32'h150):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire151;
  input wire [(5'h10):(1'h0)] wire150;
  input wire [(3'h5):(1'h0)] wire149;
  input wire [(4'hc):(1'h0)] wire148;
  input wire [(4'he):(1'h0)] wire147;
  wire [(3'h6):(1'h0)] wire181;
  reg signed [(4'hb):(1'h0)] reg180 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg179 = (1'h0);
  reg [(4'hc):(1'h0)] reg178 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg177 = (1'h0);
  reg [(2'h3):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg175 = (1'h0);
  reg [(3'h5):(1'h0)] reg174 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg173 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg172 = (1'h0);
  reg [(4'hc):(1'h0)] reg171 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg170 = (1'h0);
  reg [(4'hd):(1'h0)] reg169 = (1'h0);
  reg [(5'h15):(1'h0)] reg168 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg167 = (1'h0);
  reg [(5'h13):(1'h0)] reg166 = (1'h0);
  reg [(4'he):(1'h0)] reg165 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg164 = (1'h0);
  reg [(4'h8):(1'h0)] reg163 = (1'h0);
  reg [(3'h6):(1'h0)] reg162 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg161 = (1'h0);
  reg [(3'h6):(1'h0)] reg160 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg159 = (1'h0);
  reg [(4'hf):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg157 = (1'h0);
  wire [(3'h4):(1'h0)] wire156;
  wire [(4'hf):(1'h0)] wire155;
  wire signed [(3'h4):(1'h0)] wire154;
  wire signed [(4'hf):(1'h0)] wire153;
  wire signed [(4'he):(1'h0)] wire152;
  assign y = {wire181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 wire156,
                 wire155,
                 wire154,
                 wire153,
                 wire152,
                 (1'h0)};
  assign wire152 = wire149[(3'h5):(3'h5)];
  assign wire153 = (^$signed($signed($signed((wire147 ? (8'hb2) : wire152)))));
  assign wire154 = (+($unsigned($unsigned($signed(wire151))) ?
                       $signed((wire153 ?
                           (7'h44) : wire147[(3'h4):(2'h3)])) : wire149));
  assign wire155 = wire152[(3'h4):(1'h0)];
  assign wire156 = $unsigned(wire154[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      if ($signed($unsigned($signed((+$unsigned(wire155))))))
        begin
          reg157 <= $unsigned($signed({((wire148 ?
                  (8'ha0) : wire153) + (7'h40)),
              wire149}));
        end
      else
        begin
          reg157 <= reg157;
          if (wire155)
            begin
              reg158 <= ((wire156[(2'h2):(1'h0)] >> wire155) ?
                  (+($signed($unsigned((8'h9d))) ?
                      (((8'hb4) ?
                          wire150 : wire155) || $signed(wire149)) : $unsigned((8'h9c)))) : $signed((((7'h42) ?
                      (wire147 ? wire148 : wire152) : (wire147 ?
                          reg157 : wire153)) <<< wire149[(2'h2):(1'h0)])));
              reg159 <= reg157;
              reg160 <= (wire155[(3'h5):(2'h3)] ?
                  reg158 : (&(wire152[(4'he):(1'h1)] | wire152)));
              reg161 <= wire152;
              reg162 <= wire148;
            end
          else
            begin
              reg158 <= wire152[(4'he):(4'h8)];
              reg159 <= {(~&(~wire154)), $unsigned(wire152[(3'h6):(1'h0)])};
              reg160 <= {wire152[(4'hb):(1'h0)]};
            end
          reg163 <= {wire156};
        end
      if (($signed(({reg160[(1'h0):(1'h0)],
              $unsigned(wire152)} < $signed(wire153))) ?
          {{{(8'hbd)},
                  ((wire147 ?
                      reg161 : wire151) >> reg158)}} : (wire147 >> $unsigned((reg160[(3'h6):(1'h1)] ?
              (reg161 ? wire148 : wire151) : $unsigned(reg157))))))
        begin
          reg164 <= {((-(~$unsigned(reg158))) ?
                  wire153[(4'he):(4'hd)] : $unsigned($unsigned(reg157[(3'h5):(3'h5)]))),
              (~&wire147)};
          if (($unsigned($signed(wire156[(1'h1):(1'h0)])) ~^ $unsigned(reg158[(4'h9):(3'h4)])))
            begin
              reg165 <= (^~wire154);
              reg166 <= wire152[(1'h0):(1'h0)];
              reg167 <= {{reg162[(1'h1):(1'h0)],
                      ($unsigned($unsigned(reg160)) ?
                          $unsigned(reg160[(3'h5):(3'h4)]) : $unsigned(reg162[(3'h5):(3'h4)]))}};
              reg168 <= ($signed(reg157) + (&{$signed($unsigned(reg158)),
                  $unsigned($signed((8'haa)))}));
              reg169 <= reg166;
            end
          else
            begin
              reg165 <= reg167;
              reg166 <= reg165[(3'h7):(3'h4)];
            end
          reg170 <= $unsigned(reg162[(3'h4):(1'h0)]);
        end
      else
        begin
          reg164 <= $signed($signed(wire147[(3'h4):(3'h4)]));
          reg165 <= (+(+($unsigned(((8'hbd) ? (8'ha0) : reg159)) ?
              (reg168[(4'hf):(4'h9)] && reg167) : $unsigned((reg163 ?
                  wire154 : (8'ha2))))));
          reg166 <= (wire150 == $signed($signed(({(8'ha6),
              reg158} ^ (reg158 & reg165)))));
          reg167 <= $signed(reg169[(4'hd):(4'hc)]);
          reg168 <= (($unsigned($signed(reg168)) <<< $signed(((reg157 ?
                      reg160 : (8'hbe)) ?
                  {reg169, wire147} : (reg165 >= reg161)))) ?
              $signed(reg169) : ((^~$signed((reg157 == wire152))) + wire149[(3'h5):(3'h4)]));
        end
      if ((reg157 ? reg158 : {reg165}))
        begin
          reg171 <= wire153;
          reg172 <= $signed((+$unsigned(((reg165 ?
              reg166 : wire151) | wire154))));
          if (wire155[(2'h2):(1'h0)])
            begin
              reg173 <= $unsigned(reg162);
              reg174 <= ((((^~(reg159 != wire149)) - {(reg172 | reg162)}) + ({reg164[(4'hf):(2'h2)],
                      reg172} ?
                  $unsigned({reg157,
                      reg161}) : $signed($unsigned(reg160)))) && reg157);
              reg175 <= wire148[(4'h9):(2'h3)];
              reg176 <= {$unsigned(wire150[(4'hb):(1'h1)]), (8'hb8)};
            end
          else
            begin
              reg173 <= $signed((~$signed($signed((reg163 - reg167)))));
            end
          reg177 <= (($signed(reg161[(3'h5):(3'h5)]) < reg174[(1'h0):(1'h0)]) ?
              (((!wire155) ^~ wire148[(1'h0):(1'h0)]) ?
                  {reg165,
                      $unsigned(wire147[(3'h5):(2'h2)])} : $signed(reg158[(3'h6):(3'h5)])) : $signed((wire154 ?
                  ($unsigned(reg163) ?
                      (reg173 >= reg165) : (8'ha4)) : ((reg164 ^~ (8'hbf)) ?
                      reg157[(3'h4):(3'h4)] : ((7'h41) ? wire154 : reg171)))));
          reg178 <= (($unsigned($signed((reg172 ? wire151 : (8'hb3)))) ?
                  {(|(&reg165)), (|(8'ha1))} : $signed((wire154[(1'h0):(1'h0)] ?
                      ((8'hbc) < reg162) : wire153[(4'hc):(4'h9)]))) ?
              $unsigned((^(reg173 + $signed(reg163)))) : ((|{(8'ha8)}) ^~ ((+(+reg168)) ?
                  reg170[(1'h1):(1'h1)] : (^(wire148 ? reg170 : reg161)))));
        end
      else
        begin
          reg171 <= $signed(((reg172[(1'h1):(1'h0)] ?
              wire148 : $signed({reg175})) < (~|wire156)));
          reg172 <= {(({{reg168, reg172},
                      (reg157 ?
                          wire147 : wire150)} <<< $unsigned($signed(reg160))) ?
                  (+(~|$signed(reg169))) : reg177[(4'h8):(3'h4)]),
              ({$signed($signed(reg167)),
                      (reg158[(4'h8):(3'h6)] + $unsigned(reg162))} ?
                  wire150 : (!({(8'hb2)} << reg157[(4'hf):(4'hc)])))};
          if ($signed($signed($unsigned(reg168[(2'h2):(1'h1)]))))
            begin
              reg173 <= (wire156[(2'h3):(2'h2)] ?
                  reg166[(3'h5):(1'h1)] : (-$unsigned(($signed(reg167) && (reg170 != wire149)))));
            end
          else
            begin
              reg173 <= ($signed(((^{(8'hbc)}) ?
                  ((wire150 ?
                      (8'ha0) : wire147) ^ (!reg176)) : ($signed(wire150) + (reg178 ?
                      wire152 : reg161)))) ^~ {{$unsigned((reg176 | reg177)),
                      wire155},
                  $signed($signed((reg177 || (8'h9f))))});
              reg174 <= (^(~(~|reg170[(2'h2):(2'h2)])));
              reg175 <= $signed(((~|{reg171, $unsigned(reg168)}) ?
                  ((^~reg167) - $signed({(8'ha6)})) : $signed($unsigned((wire151 >> (7'h44))))));
              reg176 <= reg159[(3'h4):(3'h4)];
            end
          reg177 <= reg170;
          if (reg171[(4'hc):(3'h4)])
            begin
              reg178 <= $unsigned($unsigned(reg178));
              reg179 <= {$unsigned(reg165[(1'h1):(1'h0)])};
              reg180 <= ({((-reg172[(4'h9):(1'h1)]) ?
                      $unsigned((wire155 | reg179)) : reg160[(3'h5):(1'h1)]),
                  ((~^(~|(8'hb1))) && reg167)} + $unsigned($unsigned(($unsigned((8'hb1)) ~^ $unsigned(reg162)))));
            end
          else
            begin
              reg178 <= (|$unsigned(reg163[(1'h1):(1'h1)]));
              reg179 <= ((!wire153) != wire155[(3'h6):(3'h6)]);
              reg180 <= (7'h41);
            end
        end
    end
  assign wire181 = {(~|$signed((8'hb3)))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module105
#( parameter param142 = (((-(~&((8'hb0) + (7'h44)))) < {(((7'h44) ? (8'ha2) : (8'hac)) - {(8'haa), (8'hae)}), (8'hab)}) ? (^~{{((8'ha1) ? (8'hb7) : (7'h43)), ((8'ha1) ^~ (8'haa))}}) : (8'ha7))
, parameter param143 = (~param142) )
(y, clk, wire109, wire108, wire107, wire106);
  output wire [(32'h18c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire109;
  input wire signed [(2'h3):(1'h0)] wire108;
  input wire signed [(3'h5):(1'h0)] wire107;
  input wire signed [(4'h9):(1'h0)] wire106;
  wire signed [(5'h12):(1'h0)] wire141;
  wire signed [(4'hb):(1'h0)] wire140;
  reg [(4'hc):(1'h0)] reg139 = (1'h0);
  reg [(5'h13):(1'h0)] reg138 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg137 = (1'h0);
  reg [(5'h10):(1'h0)] reg136 = (1'h0);
  reg [(4'h8):(1'h0)] reg135 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg134 = (1'h0);
  reg [(3'h5):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg132 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg131 = (1'h0);
  reg [(4'ha):(1'h0)] reg130 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg129 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg128 = (1'h0);
  reg [(3'h4):(1'h0)] reg127 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg126 = (1'h0);
  reg [(5'h15):(1'h0)] reg125 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg124 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg123 = (1'h0);
  reg [(3'h5):(1'h0)] reg122 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg121 = (1'h0);
  reg [(5'h14):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg119 = (1'h0);
  reg [(4'he):(1'h0)] reg118 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg117 = (1'h0);
  reg [(4'ha):(1'h0)] reg116 = (1'h0);
  reg [(5'h13):(1'h0)] reg115 = (1'h0);
  reg [(5'h13):(1'h0)] reg114 = (1'h0);
  reg [(4'he):(1'h0)] reg113 = (1'h0);
  reg [(5'h12):(1'h0)] reg112 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg111 = (1'h0);
  wire [(4'hd):(1'h0)] wire110;
  assign y = {wire141,
                 wire140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 wire110,
                 (1'h0)};
  assign wire110 = (~&wire106[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      if ($signed({(~wire107[(1'h1):(1'h0)])}))
        begin
          reg111 <= (({(wire106[(1'h0):(1'h0)] >> {(8'hb1)}),
                      {(^wire110), $signed((8'ha1))}} ?
                  ($unsigned((wire109 ^~ wire109)) != wire108[(1'h1):(1'h0)]) : (+{(+wire108),
                      wire107[(3'h4):(1'h1)]})) ?
              ((wire107 ?
                      ((wire107 < wire108) >> ((8'hb1) ?
                          wire106 : wire108)) : wire108[(1'h0):(1'h0)]) ?
                  (&wire108[(2'h3):(1'h1)]) : wire107) : (wire109[(3'h4):(3'h4)] ?
                  wire110 : (&(((8'ha8) ? wire107 : (8'hbc)) ?
                      wire109[(1'h1):(1'h1)] : (wire110 ?
                          wire108 : wire108)))));
          reg112 <= (reg111 + ({((~(8'ha7)) ?
                      reg111 : (wire109 ? reg111 : wire110)),
                  $signed((~wire107))} ?
              (wire108 ?
                  ({reg111} & (reg111 ?
                      wire110 : (8'hbe))) : (^~(8'h9c))) : $unsigned(((wire110 ?
                      wire110 : wire109) ?
                  (!wire107) : (wire109 ? wire108 : wire110)))));
          if ((8'hbf))
            begin
              reg113 <= reg111[(2'h2):(1'h1)];
              reg114 <= (((+(7'h44)) ?
                      (((wire110 ? (7'h43) : (7'h43)) ?
                              {wire108} : (&wire108)) ?
                          wire110 : ($unsigned(wire106) ?
                              $signed((8'hac)) : wire109)) : ((8'ha0) ^ wire110)) ?
                  reg112[(3'h7):(2'h3)] : $unsigned($unsigned(wire109[(2'h3):(1'h0)])));
            end
          else
            begin
              reg113 <= reg114[(1'h1):(1'h0)];
              reg114 <= (wire108 * ((reg114[(5'h10):(3'h4)] ?
                      {$signed(reg112)} : $signed(reg111[(2'h3):(1'h1)])) ?
                  $signed(wire109) : wire108));
              reg115 <= ((+(($unsigned(reg112) >= $signed(wire106)) ?
                      wire106[(1'h1):(1'h0)] : $unsigned(wire110))) ?
                  (wire109[(1'h1):(1'h0)] ?
                      (&reg112[(4'h9):(2'h3)]) : $unsigned(wire110)) : reg114);
              reg116 <= reg113[(4'hb):(3'h5)];
              reg117 <= {($unsigned(reg115) * wire108[(2'h3):(2'h3)])};
            end
          reg118 <= $signed($signed(wire106));
          reg119 <= reg112[(4'hf):(4'hf)];
        end
      else
        begin
          reg111 <= reg117;
          reg112 <= $unsigned(reg114);
        end
      if (wire106)
        begin
          if ((~&wire108[(2'h3):(1'h0)]))
            begin
              reg120 <= $unsigned((&(~^(^~$unsigned(wire107)))));
            end
          else
            begin
              reg120 <= ($unsigned({$unsigned(reg113[(4'hb):(3'h7)])}) ?
                  $signed((-(!reg119[(1'h0):(1'h0)]))) : (~^$unsigned({wire107[(1'h1):(1'h1)]})));
              reg121 <= ({(+(8'ha7)), ($signed({wire110, reg116}) > (8'ha5))} ?
                  wire106 : ((^~(reg113[(1'h1):(1'h0)] ?
                      $unsigned(reg120) : (!reg120))) ^~ (^~wire108)));
              reg122 <= {$unsigned($signed($unsigned(reg119[(3'h4):(1'h1)]))),
                  reg121[(3'h5):(2'h3)]};
            end
          reg123 <= {(^~(~((~^reg116) | (~&wire107)))),
              ((|reg119[(4'h8):(1'h1)]) < $signed(reg119[(3'h6):(1'h0)]))};
        end
      else
        begin
          if ($unsigned($signed((($unsigned((8'hb8)) + (^~reg115)) ?
              $unsigned(((7'h43) >>> (8'hb0))) : $unsigned(reg118[(4'h8):(4'h8)])))))
            begin
              reg120 <= {(8'hb9), wire108};
            end
          else
            begin
              reg120 <= wire108;
            end
        end
      reg124 <= $unsigned($unsigned(($unsigned((reg118 ? reg115 : reg117)) ?
          (reg122[(3'h4):(1'h0)] ?
              {reg123, (8'hab)} : $signed((7'h41))) : reg115)));
      reg125 <= ((^~wire107[(1'h1):(1'h0)]) != reg112[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg126 <= (-reg120[(4'h8):(1'h0)]);
      if ({((~|(7'h40)) ? (&(reg118 << (8'hb0))) : {$unsigned({reg118})}),
          (&$unsigned(($unsigned((8'h9d)) ?
              $unsigned(reg123) : (reg114 - reg122))))})
        begin
          reg127 <= reg112[(5'h12):(1'h1)];
          if ($unsigned($signed(reg122[(1'h1):(1'h1)])))
            begin
              reg128 <= $signed((reg127 - (~|reg116[(3'h4):(2'h3)])));
              reg129 <= {$unsigned((((reg123 != reg123) ?
                          $signed(reg111) : ((8'ha8) ^~ wire107)) ?
                      ((reg117 * reg119) ?
                          ((7'h44) | wire110) : {wire107}) : reg117[(4'hc):(4'ha)]))};
            end
          else
            begin
              reg128 <= ((^~(-reg118[(4'he):(3'h6)])) ?
                  (8'hac) : ($unsigned(reg119[(2'h3):(1'h1)]) ?
                      (^~(~|{reg123,
                          reg124})) : $signed($signed(reg129[(3'h6):(2'h2)]))));
            end
        end
      else
        begin
          reg127 <= {reg114[(4'hd):(4'hd)],
              ((($signed(wire109) ?
                  (!(8'ha1)) : (reg127 ?
                      reg119 : reg126)) << $unsigned({(8'hba)})) & $signed(reg126[(4'h9):(4'h8)]))};
          reg128 <= $unsigned(reg128);
          if ($unsigned((8'hae)))
            begin
              reg129 <= (reg119 ~^ wire108[(2'h2):(2'h2)]);
              reg130 <= {reg122, {(|($unsigned(reg129) < (7'h44)))}};
              reg131 <= $signed(((&(wire108 ?
                  $signed(reg122) : (reg111 <<< reg125))) | reg116[(2'h2):(1'h1)]));
              reg132 <= $unsigned($unsigned((($signed(reg128) > (wire106 <= (8'hb6))) ?
                  ((^~reg131) == (reg114 == reg130)) : {(reg126 <<< reg115),
                      reg129[(2'h2):(1'h1)]})));
              reg133 <= reg116[(3'h5):(1'h1)];
            end
          else
            begin
              reg129 <= $signed($unsigned(reg127[(3'h4):(2'h3)]));
              reg130 <= $signed(reg115[(1'h1):(1'h1)]);
              reg131 <= $unsigned(reg113);
            end
        end
      reg134 <= wire107[(1'h0):(1'h0)];
      if (reg123[(2'h2):(2'h2)])
        begin
          reg135 <= wire108;
          reg136 <= reg114;
          reg137 <= (8'ha0);
        end
      else
        begin
          reg135 <= $signed($unsigned($unsigned(wire110[(4'hc):(3'h5)])));
        end
      if ($unsigned(reg115))
        begin
          reg138 <= $signed($signed({reg119[(2'h3):(1'h1)],
              ($unsigned(reg137) ?
                  (wire106 ? reg122 : reg120) : ((8'hb7) != reg125))}));
          reg139 <= (8'hab);
        end
      else
        begin
          reg138 <= $unsigned($signed(wire106));
        end
    end
  assign wire140 = $unsigned($unsigned(reg116));
  assign wire141 = (7'h44);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module273
#( parameter param283 = {{((((8'ha9) ? (8'hb8) : (8'hb3)) ^~ {(8'ha0)}) && (((8'hb5) >> (8'h9d)) ? (~|(7'h42)) : (~^(7'h40)))), (+(((8'ha7) >>> (8'hb2)) ? ((8'had) ? (8'ha7) : (8'hb9)) : ((8'hb1) ? (8'h9c) : (8'hb9))))}} )
(y, clk, wire277, wire276, wire275, wire274);
  output wire [(32'h33):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire277;
  input wire signed [(2'h3):(1'h0)] wire276;
  input wire [(5'h11):(1'h0)] wire275;
  input wire [(5'h15):(1'h0)] wire274;
  wire signed [(4'hb):(1'h0)] wire282;
  wire [(4'hb):(1'h0)] wire281;
  wire [(4'h8):(1'h0)] wire280;
  wire [(4'hd):(1'h0)] wire279;
  wire [(3'h7):(1'h0)] wire278;
  assign y = {wire282, wire281, wire280, wire279, wire278, (1'h0)};
  assign wire278 = (&$unsigned({wire277, wire276[(2'h3):(2'h3)]}));
  assign wire279 = ($unsigned($signed(($unsigned(wire276) ^ $signed((8'had))))) * (wire275 > $signed(wire278)));
  assign wire280 = $unsigned(((^(~^(wire278 + wire277))) ?
                       {wire274[(5'h15):(4'hc)]} : (&((|(8'ha2)) ?
                           $unsigned(wire274) : $unsigned(wire274)))));
  assign wire281 = ($unsigned(((^(wire274 ? wire275 : wire275)) ?
                       (wire279[(4'hc):(3'h5)] ?
                           wire279[(1'h0):(1'h0)] : wire274) : ((&wire275) >> $signed((8'ha0))))) | $unsigned((wire275 >>> {(wire274 ?
                           wire280 : wire277),
                       (^~wire278)})));
  assign wire282 = (($signed(((~wire275) ?
                           $unsigned(wire281) : $signed((8'hb3)))) ?
                       (wire275[(4'h9):(1'h1)] ?
                           $unsigned(((7'h41) ?
                               wire275 : (8'hbd))) : ((|(8'hbb)) ?
                               wire279[(2'h3):(2'h3)] : wire278[(3'h5):(1'h1)])) : ((^wire277[(4'h9):(4'h8)]) ?
                           $unsigned(((8'ha0) ?
                               (8'ha4) : (8'ha4))) : (wire278[(3'h5):(3'h4)] >> wire274))) > ({{wire274},
                       $unsigned({wire280})} ~^ $unsigned($signed((wire280 ?
                       wire276 : wire275)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module246
#( parameter param260 = {(~(^(~((8'ha4) <<< (8'haa)))))}
, parameter param261 = ((param260 >= (param260 ? ((8'hac) ? ((8'hb2) >= param260) : (param260 >>> (8'h9c))) : ({param260, param260} ? {param260} : (param260 ? param260 : param260)))) ? ((^~param260) ^ param260) : {param260}) )
(y, clk, wire251, wire250, wire249, wire248, wire247);
  output wire [(32'h44):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire251;
  input wire [(4'hf):(1'h0)] wire250;
  input wire [(4'he):(1'h0)] wire249;
  input wire signed [(3'h5):(1'h0)] wire248;
  input wire signed [(5'h13):(1'h0)] wire247;
  wire [(4'hf):(1'h0)] wire259;
  wire signed [(3'h6):(1'h0)] wire258;
  wire signed [(3'h6):(1'h0)] wire257;
  wire signed [(3'h6):(1'h0)] wire256;
  reg signed [(3'h6):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg254 = (1'h0);
  wire [(4'h9):(1'h0)] wire253;
  wire [(2'h2):(1'h0)] wire252;
  assign y = {wire259,
                 wire258,
                 wire257,
                 wire256,
                 reg255,
                 reg254,
                 wire253,
                 wire252,
                 (1'h0)};
  assign wire252 = (7'h44);
  assign wire253 = (^wire250[(3'h7):(2'h2)]);
  always
    @(posedge clk) begin
      reg254 <= wire252[(2'h2):(1'h1)];
      reg255 <= ({$signed((wire249 ^ (wire247 | wire249)))} > wire253[(1'h1):(1'h1)]);
    end
  assign wire256 = reg254[(2'h2):(1'h1)];
  assign wire257 = wire248;
  assign wire258 = ((~^(~(wire247 ? (~|wire251) : wire251))) ?
                       $signed((((~^reg255) > $unsigned(wire247)) ?
                           $unsigned(wire250) : wire248)) : ((wire253 ?
                           (~$signed(reg254)) : (~&$signed(wire257))) >= {$unsigned((~^(8'hb6))),
                           (wire252 - ((8'haa) ^ reg254))}));
  assign wire259 = (~&wire258);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module223  (y, clk, wire227, wire226, wire225, wire224);
  output wire [(32'h7a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire227;
  input wire [(5'h10):(1'h0)] wire226;
  input wire signed [(4'ha):(1'h0)] wire225;
  input wire [(5'h12):(1'h0)] wire224;
  wire [(4'hc):(1'h0)] wire237;
  wire signed [(5'h11):(1'h0)] wire236;
  reg signed [(4'ha):(1'h0)] reg235 = (1'h0);
  wire [(4'hd):(1'h0)] wire234;
  wire signed [(5'h11):(1'h0)] wire233;
  wire signed [(4'ha):(1'h0)] wire232;
  wire signed [(4'hf):(1'h0)] wire231;
  wire signed [(4'h8):(1'h0)] wire230;
  wire signed [(4'ha):(1'h0)] wire229;
  wire [(4'h9):(1'h0)] wire228;
  assign y = {wire237,
                 wire236,
                 reg235,
                 wire234,
                 wire233,
                 wire232,
                 wire231,
                 wire230,
                 wire229,
                 wire228,
                 (1'h0)};
  assign wire228 = (&wire224[(4'h8):(3'h4)]);
  assign wire229 = (8'hba);
  assign wire230 = ((wire226 >= $unsigned($signed((8'hb9)))) ?
                       (+$unsigned(($unsigned(wire226) + wire226))) : wire224);
  assign wire231 = (wire225 >>> (~&(+wire228)));
  assign wire232 = wire226;
  assign wire233 = (wire231 <= (wire231[(4'he):(4'hb)] ^~ (7'h40)));
  assign wire234 = (~^(wire231[(2'h2):(1'h1)] ^~ {((wire231 ?
                               wire225 : wire230) ?
                           (wire231 ? (8'hab) : wire227) : wire224)}));
  always
    @(posedge clk) begin
      reg235 <= ((~^(^{wire232[(4'h9):(2'h2)], wire226[(4'hf):(4'hb)]})) ?
          wire227 : wire224);
    end
  assign wire236 = wire231[(3'h4):(1'h0)];
  assign wire237 = (8'hb5);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module314
#( parameter param413 = {({(!(8'hbd))} <= (~(((8'ha3) > (8'hae)) ? ((7'h44) ? (8'ha8) : (8'hab)) : (8'haf)))), (+{({(8'haa)} > (!(7'h40))), ((^(8'hbe)) ? ((8'hb0) ? (8'ha9) : (8'h9c)) : {(8'hb2), (8'hbf)})})}
, parameter param414 = ({(^(param413 ~^ {(8'hac), (8'hb2)}))} ? param413 : (|((~&(^param413)) ? (((8'hbf) << param413) ? (~&(8'hbc)) : (param413 ~^ param413)) : (&param413)))) )
(y, clk, wire315, wire316, wire317, wire318, wire319);
  output wire [(32'hed):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire315;
  input wire [(5'h14):(1'h0)] wire316;
  input wire signed [(5'h13):(1'h0)] wire317;
  input wire [(5'h11):(1'h0)] wire318;
  input wire signed [(4'h8):(1'h0)] wire319;
  wire signed [(5'h12):(1'h0)] wire412;
  reg [(5'h13):(1'h0)] reg411 = (1'h0);
  reg [(2'h3):(1'h0)] reg410 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg409 = (1'h0);
  reg [(5'h12):(1'h0)] reg408 = (1'h0);
  reg [(4'h8):(1'h0)] reg407 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg406 = (1'h0);
  reg [(4'ha):(1'h0)] reg405 = (1'h0);
  reg [(4'h9):(1'h0)] reg404 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg403 = (1'h0);
  reg [(4'hd):(1'h0)] reg402 = (1'h0);
  reg [(4'hf):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg400 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg399 = (1'h0);
  reg signed [(4'he):(1'h0)] reg398 = (1'h0);
  wire [(3'h4):(1'h0)] wire397;
  wire [(3'h7):(1'h0)] wire396;
  wire [(5'h13):(1'h0)] wire395;
  wire signed [(5'h10):(1'h0)] wire394;
  wire signed [(3'h4):(1'h0)] wire392;
  assign y = {wire412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 wire397,
                 wire396,
                 wire395,
                 wire394,
                 wire392,
                 (1'h0)};
  module320 modinst393 (.clk(clk), .wire325(wire317), .wire321(wire318), .wire322(wire316), .wire324(wire315), .wire323(wire319), .y(wire392));
  assign wire394 = (^wire315[(3'h4):(3'h4)]);
  assign wire395 = ({(({wire315, (8'haf)} ? wire394 : (wire315 < wire317)) ?
                               $signed((wire394 > (8'hb6))) : wire315[(4'h9):(2'h3)]),
                           (($unsigned((8'ha6)) - wire392) + (!$unsigned(wire392)))} ?
                       (wire319 ~^ ((wire318[(3'h7):(3'h6)] || (&(8'ha1))) == wire317[(4'h9):(1'h1)])) : {(+$unsigned(wire318))});
  assign wire396 = $signed((($unsigned((wire395 ^ wire392)) != (wire392[(1'h1):(1'h0)] ?
                           $unsigned((7'h44)) : {wire319, wire315})) ?
                       $signed($signed($signed(wire315))) : ($signed(wire317[(1'h0):(1'h0)]) << wire316[(5'h14):(5'h12)])));
  assign wire397 = ((+($signed((8'ha2)) >= $unsigned($unsigned(wire392)))) ?
                       ($unsigned((~&(wire318 * wire316))) ?
                           $unsigned(wire396[(2'h3):(2'h3)]) : (~&wire394)) : $signed(wire318));
  always
    @(posedge clk) begin
      reg398 <= ((wire395 ?
          $unsigned({(+wire316)}) : ((wire315 == $unsigned(wire317)) >>> wire397[(3'h4):(1'h1)])) ^~ $unsigned($unsigned((|(wire395 ?
          wire397 : (8'had))))));
      if (((((wire316 && (8'hac)) > ((wire392 ? wire397 : (8'hb1)) ?
          {(8'hb7)} : (~^reg398))) ^ $signed(($signed(reg398) ?
          (!wire392) : wire397[(2'h2):(1'h0)]))) > (~|wire396)))
        begin
          reg399 <= $unsigned($signed(wire318));
          reg400 <= $signed(wire316[(5'h14):(4'hd)]);
          reg401 <= wire318;
        end
      else
        begin
          reg399 <= (^$signed($signed($signed((wire317 + wire318)))));
          reg400 <= {$signed($signed($unsigned((-reg398)))),
              ({wire316} == ((^~reg401[(2'h3):(2'h2)]) <<< ($unsigned(wire319) ?
                  $unsigned(wire397) : (wire316 - wire317))))};
        end
      reg402 <= (7'h42);
      if (($signed($unsigned((!wire318))) ?
          (wire318[(4'hb):(1'h0)] >= wire397) : $signed((&$unsigned($signed(reg400))))))
        begin
          reg403 <= ((~|{$signed((wire318 ? wire316 : reg401))}) ?
              $signed(wire397) : $unsigned(($signed((wire392 ?
                  wire316 : wire318)) * wire318)));
          if ($signed({(&($unsigned((8'ha7)) ?
                  $signed(wire392) : $signed((8'hae)))),
              (reg401 && $signed((reg399 ^~ wire392)))}))
            begin
              reg404 <= $signed(({(+wire392),
                  (~|(^~wire315))} << reg400[(1'h0):(1'h0)]));
              reg405 <= $signed((wire394[(3'h7):(1'h0)] == $signed((~$unsigned(reg403)))));
              reg406 <= (+wire316);
            end
          else
            begin
              reg404 <= wire319;
            end
          if ($signed($signed(wire395)))
            begin
              reg407 <= reg406[(3'h6):(1'h0)];
              reg408 <= (~$unsigned({($unsigned(reg400) >> (wire318 << wire316))}));
              reg409 <= reg402[(4'hd):(4'hc)];
              reg410 <= {reg404[(3'h4):(2'h3)]};
              reg411 <= (^$signed((wire315 == reg398)));
            end
          else
            begin
              reg407 <= $unsigned($unsigned((reg399 ?
                  (!(~|reg403)) : $signed(wire395))));
              reg408 <= $signed((($unsigned(reg407[(1'h0):(1'h0)]) ?
                  $unsigned((wire318 ?
                      wire396 : wire395)) : (wire396[(2'h2):(1'h0)] ?
                      reg404 : $unsigned(reg404))) & $unsigned(((reg411 ?
                  reg405 : wire318) << (reg410 * wire315)))));
            end
        end
      else
        begin
          reg403 <= (+({$signed({(8'ha9), wire318})} ?
              ($signed((wire397 == reg408)) ?
                  reg400[(4'hd):(3'h5)] : ({reg402,
                      (8'hb2)} | ((8'hb6) ^ wire318))) : ((wire396[(2'h3):(2'h2)] ?
                  ((8'hac) < wire318) : wire318) ~^ ((reg407 ?
                  wire315 : reg411) && $signed(reg411)))));
          reg404 <= (-wire397[(1'h1):(1'h1)]);
        end
    end
  assign wire412 = $signed(reg404[(3'h7):(1'h0)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module320  (y, clk, wire325, wire324, wire323, wire322, wire321);
  output wire [(32'h2ed):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire325;
  input wire signed [(2'h2):(1'h0)] wire324;
  input wire signed [(4'h8):(1'h0)] wire323;
  input wire signed [(5'h14):(1'h0)] wire322;
  input wire signed [(5'h11):(1'h0)] wire321;
  wire [(4'hb):(1'h0)] wire391;
  reg signed [(5'h10):(1'h0)] reg390 = (1'h0);
  reg [(2'h2):(1'h0)] reg389 = (1'h0);
  reg [(3'h5):(1'h0)] reg388 = (1'h0);
  reg [(4'ha):(1'h0)] reg387 = (1'h0);
  reg [(5'h13):(1'h0)] reg386 = (1'h0);
  reg [(5'h11):(1'h0)] reg385 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg384 = (1'h0);
  reg [(4'hf):(1'h0)] reg383 = (1'h0);
  reg [(4'he):(1'h0)] reg382 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg381 = (1'h0);
  reg [(4'hb):(1'h0)] reg380 = (1'h0);
  reg [(5'h10):(1'h0)] reg379 = (1'h0);
  reg [(3'h6):(1'h0)] reg378 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg377 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg376 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg375 = (1'h0);
  reg signed [(4'he):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg373 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg372 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg371 = (1'h0);
  reg [(2'h3):(1'h0)] reg370 = (1'h0);
  reg [(5'h14):(1'h0)] reg369 = (1'h0);
  reg [(3'h7):(1'h0)] reg368 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg366 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg365 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg363 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg362 = (1'h0);
  reg [(5'h13):(1'h0)] reg361 = (1'h0);
  reg [(4'ha):(1'h0)] reg360 = (1'h0);
  reg [(4'hd):(1'h0)] reg359 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg358 = (1'h0);
  reg [(4'ha):(1'h0)] reg357 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg356 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg355 = (1'h0);
  wire [(5'h11):(1'h0)] wire354;
  wire [(5'h10):(1'h0)] wire353;
  wire signed [(4'hb):(1'h0)] wire352;
  reg signed [(4'hb):(1'h0)] reg351 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg350 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg349 = (1'h0);
  reg [(4'hc):(1'h0)] reg348 = (1'h0);
  reg [(4'h8):(1'h0)] reg347 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire346;
  wire signed [(4'h8):(1'h0)] wire345;
  wire [(2'h3):(1'h0)] wire344;
  wire [(3'h5):(1'h0)] wire343;
  reg [(4'hc):(1'h0)] reg342 = (1'h0);
  reg [(3'h5):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg340 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg339 = (1'h0);
  reg [(3'h7):(1'h0)] reg338 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg337 = (1'h0);
  reg [(5'h13):(1'h0)] reg336 = (1'h0);
  reg [(2'h2):(1'h0)] reg335 = (1'h0);
  reg [(5'h15):(1'h0)] reg334 = (1'h0);
  reg [(4'h8):(1'h0)] reg333 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg332 = (1'h0);
  reg [(3'h4):(1'h0)] reg331 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire330;
  wire [(4'hc):(1'h0)] wire329;
  wire signed [(4'he):(1'h0)] wire328;
  reg [(4'hf):(1'h0)] reg327 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg326 = (1'h0);
  assign y = {wire391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 wire354,
                 wire353,
                 wire352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 wire346,
                 wire345,
                 wire344,
                 wire343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 wire330,
                 wire329,
                 wire328,
                 reg327,
                 reg326,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg326 <= (^~($unsigned(wire324) - wire324));
      reg327 <= ((reg326[(3'h7):(3'h7)] << ($unsigned((|wire321)) - ((wire323 * reg326) == (wire324 || (8'hb5))))) & wire322);
    end
  assign wire328 = wire321;
  assign wire329 = {($signed((!$unsigned(wire322))) >>> ((~|wire323) ?
                           ((wire325 ?
                               wire321 : (8'hbb)) <<< (~^(8'ha5))) : wire325))};
  assign wire330 = $unsigned((reg326 < {((wire328 ?
                           wire328 : wire324) & ((8'hbb) ?
                           wire323 : wire325))}));
  always
    @(posedge clk) begin
      if (wire321)
        begin
          reg331 <= ((-wire328) ?
              (8'ha6) : {wire322[(4'hf):(3'h7)],
                  (((wire325 <<< reg326) >>> (reg327 > wire321)) ?
                      wire325[(4'h8):(3'h4)] : reg327[(4'hc):(4'ha)])});
          reg332 <= wire330;
          if (((^~wire321) ? (8'ha3) : wire330))
            begin
              reg333 <= (($signed({(^~reg326)}) ~^ (+{(wire323 >> wire322),
                  wire321})) == ((wire325[(4'hc):(3'h5)] ?
                  (~(wire324 ?
                      wire328 : wire321)) : $unsigned((reg326 == reg327))) >> {(7'h41)}));
              reg334 <= (~|$signed($signed((8'hbb))));
              reg335 <= (8'hbb);
            end
          else
            begin
              reg333 <= ((wire328 ?
                  ($unsigned({reg327,
                      wire324}) != $unsigned((wire330 <= wire321))) : ($signed($unsigned(wire328)) ~^ (reg333[(2'h3):(2'h3)] ?
                      $signed(reg334) : $signed(reg334)))) & wire328[(3'h5):(1'h0)]);
              reg334 <= ({(8'hb1),
                      ($signed($unsigned(wire328)) < (reg332 ~^ (+wire321)))} ?
                  ($unsigned(((8'hba) ?
                          $unsigned(reg332) : (wire324 == (8'hb2)))) ?
                      ({$signed(wire328)} != (~(reg332 ^ wire324))) : wire329[(1'h0):(1'h0)]) : {(8'ha4)});
            end
          reg336 <= reg333[(3'h6):(1'h0)];
          if (((8'hb6) * (+reg336[(4'hf):(4'hd)])))
            begin
              reg337 <= wire323[(2'h3):(1'h0)];
              reg338 <= (reg334 ?
                  $unsigned(((^~(reg335 ? reg331 : wire323)) ?
                      $signed($signed((8'hb3))) : $unsigned((reg326 ?
                          reg334 : wire322)))) : {$signed($unsigned((~(8'hbb))))});
              reg339 <= (&wire329[(1'h1):(1'h0)]);
              reg340 <= (|(reg331 ?
                  ({(wire321 ?
                          (7'h43) : wire325)} == wire324) : (wire321 + ((wire330 < (8'hb3)) != reg332))));
              reg341 <= $unsigned($signed($unsigned(($signed(wire323) ?
                  (wire321 ^~ wire322) : {wire328, reg339}))));
            end
          else
            begin
              reg337 <= wire325[(4'hf):(3'h5)];
              reg338 <= {($signed((^wire329)) ?
                      $signed(reg334[(2'h2):(2'h2)]) : reg326[(3'h6):(2'h2)])};
              reg339 <= wire322;
              reg340 <= $unsigned((reg338 < reg336));
            end
        end
      else
        begin
          reg331 <= ({wire325[(1'h0):(1'h0)]} ^ $signed($signed((wire324 << reg334))));
        end
      reg342 <= (~|reg341);
    end
  assign wire343 = (^$unsigned(reg331));
  assign wire344 = (~&$signed($signed(reg340[(4'he):(4'ha)])));
  assign wire345 = {$signed({reg331[(1'h0):(1'h0)]})};
  assign wire346 = wire343[(3'h4):(3'h4)];
  always
    @(posedge clk) begin
      reg347 <= ($signed($signed(reg331)) ? wire345 : wire325[(3'h5):(2'h2)]);
      reg348 <= reg332[(1'h0):(1'h0)];
      reg349 <= wire346[(3'h4):(1'h1)];
      reg350 <= (((-$unsigned((^reg327))) << reg339[(3'h5):(1'h1)]) ?
          (wire321[(5'h10):(4'ha)] != $signed($signed((wire328 ?
              reg334 : reg331)))) : (8'hba));
      reg351 <= (!($signed(wire322[(4'hd):(4'hb)]) ?
          $unsigned(reg338) : {$unsigned((&wire345))}));
    end
  assign wire352 = (~wire328);
  assign wire353 = reg341[(2'h3):(1'h0)];
  assign wire354 = (({$signed(reg336[(4'hd):(2'h3)]), ((8'hb4) | (^~wire330))} ?
                       (~&{(&(8'hb5)), reg339}) : (reg332 ?
                           {(wire329 ? reg339 : reg351),
                               (reg348 >>> wire321)} : wire346)) >> (+{(~^wire329[(2'h3):(1'h1)]),
                       ((|wire344) ? reg333 : (reg327 || reg348))}));
  always
    @(posedge clk) begin
      reg355 <= (^(~{(^~((8'h9f) && reg334)), $signed(reg348[(3'h4):(2'h3)])}));
      if ($signed($unsigned((&(~reg351[(3'h4):(2'h2)])))))
        begin
          reg356 <= (~|$signed((($signed(reg327) == (!wire345)) ^ ((reg331 ?
                  wire322 : wire321) ?
              ((8'hbb) ? reg341 : wire321) : reg350[(2'h3):(2'h3)]))));
          reg357 <= (|$unsigned((8'hbf)));
        end
      else
        begin
          reg356 <= wire343;
          reg357 <= (-$signed(((|$signed(wire330)) ?
              {(8'hb6), $unsigned(wire325)} : wire323[(1'h1):(1'h1)])));
          reg358 <= (^$unsigned((({(8'ha6), wire328} ?
              $unsigned(reg335) : (-wire324)) == wire322)));
          reg359 <= (!($signed(reg347[(3'h4):(1'h1)]) ^~ ((-(~reg355)) - {$signed(reg327),
              (reg349 | wire330)})));
        end
      reg360 <= $unsigned((~|$unsigned(wire329)));
      reg361 <= reg358;
    end
  always
    @(posedge clk) begin
      reg362 <= $signed((^~reg348));
      reg363 <= $signed(wire352[(4'h9):(3'h5)]);
      if ((!{$signed($unsigned($unsigned(wire329)))}))
        begin
          reg364 <= $signed(wire322);
          reg365 <= reg348[(1'h0):(1'h0)];
          reg366 <= $signed((($unsigned($signed(wire354)) ?
                  wire330[(3'h6):(3'h5)] : $unsigned($signed(reg340))) ?
              (~(reg364[(1'h0):(1'h0)] >> reg338)) : {(reg355[(4'ha):(3'h7)] ?
                      (|reg363) : wire321[(4'hf):(1'h1)]),
                  $unsigned((wire321 ? reg336 : reg333))}));
          reg367 <= {$unsigned((((wire324 ? reg338 : reg326) && (~&(8'hae))) ?
                  (reg347[(3'h6):(1'h0)] ?
                      (reg351 >> wire321) : (reg327 * reg350)) : ((wire323 ?
                          (8'ha9) : reg339) ?
                      wire346[(3'h5):(1'h0)] : reg356)))};
        end
      else
        begin
          if ({(({(!(8'ha2))} ?
                  (wire323 ?
                      (wire343 ?
                          reg365 : (8'hab)) : reg364[(3'h5):(2'h3)]) : reg340) <= $unsigned($signed((reg333 ?
                  wire354 : reg337)))),
              reg362[(4'h8):(1'h0)]})
            begin
              reg364 <= wire324[(1'h1):(1'h1)];
              reg365 <= (^reg367);
              reg366 <= ($unsigned(((reg365 ?
                  (wire345 ?
                      wire345 : (8'haa)) : wire328) & (|$unsigned(wire352)))) >= $unsigned((-{$signed(wire321),
                  $signed(wire353)})));
              reg367 <= $unsigned($unsigned(((!$signed(wire343)) > reg337)));
              reg368 <= (7'h41);
            end
          else
            begin
              reg364 <= {reg334};
              reg365 <= (^$signed(reg366[(1'h0):(1'h0)]));
            end
          reg369 <= reg348;
        end
      reg370 <= $signed(reg338[(1'h1):(1'h0)]);
      reg371 <= (8'hb9);
    end
  always
    @(posedge clk) begin
      if ($unsigned($unsigned(reg342[(4'hb):(4'h9)])))
        begin
          reg372 <= (~|{(wire354[(3'h6):(1'h1)] >>> ((8'hb7) <<< {reg365}))});
          if (($signed($unsigned(((^reg359) << ((8'ha3) ? (8'hb7) : reg337)))) ?
              ($signed(wire329) >>> $signed(((|reg356) ?
                  $signed(wire353) : (8'hb2)))) : ($signed((+$unsigned(wire353))) ?
                  reg340 : $signed($signed($signed(reg326))))))
            begin
              reg373 <= reg331;
              reg374 <= $unsigned((($signed($signed((7'h40))) ?
                      wire325 : (reg327 ? (|wire353) : $signed(wire344))) ?
                  $signed(reg331[(2'h3):(1'h1)]) : $unsigned(reg366)));
              reg375 <= $signed((~^$unsigned((&$unsigned((8'hac))))));
              reg376 <= reg356;
              reg377 <= $signed(wire330);
            end
          else
            begin
              reg373 <= {reg377[(5'h12):(5'h12)],
                  $signed($unsigned(wire325[(5'h12):(4'hc)]))};
            end
          reg378 <= (reg340[(3'h4):(3'h4)] & {reg334[(3'h4):(3'h4)],
              {((reg326 || wire343) >> (reg327 ^ reg372))}});
          reg379 <= reg371;
        end
      else
        begin
          reg372 <= {(|((-$signed(reg377)) + (wire330[(1'h1):(1'h1)] - (reg377 ?
                  reg331 : reg364)))),
              {(~&(reg350[(3'h5):(2'h2)] - (wire325 || reg332)))}};
        end
      if ({reg368[(3'h4):(2'h2)]})
        begin
          if (reg377[(4'hc):(1'h0)])
            begin
              reg380 <= reg360[(3'h7):(1'h0)];
              reg381 <= ($signed(({reg327,
                  $unsigned(reg364)} != wire323)) ^~ (((^$signed(reg326)) < reg333) | reg369[(5'h14):(4'hd)]));
            end
          else
            begin
              reg380 <= {reg362};
              reg381 <= (($unsigned(reg373) ?
                      reg380 : (^~$signed($signed(wire325)))) ?
                  {((((8'hb7) | (8'hbb)) >> (reg358 ?
                          reg326 : reg377)) | wire325[(4'hb):(4'ha)])} : (~|reg381));
              reg382 <= ($signed($unsigned((!reg381))) ?
                  wire325 : {reg350[(3'h4):(1'h1)],
                      $signed({$signed(reg375)})});
              reg383 <= {reg342, reg360[(3'h5):(2'h3)]};
            end
          if ($unsigned({{$signed({reg370}), reg360}, wire330}))
            begin
              reg384 <= ($unsigned(reg337) - wire343);
              reg385 <= reg334;
              reg386 <= $signed(((+(-{reg374})) ?
                  reg375[(3'h7):(3'h7)] : ((8'hb4) ?
                      (8'ha7) : ({reg384, (8'hae)} ~^ reg379[(2'h3):(2'h3)]))));
              reg387 <= ($unsigned(reg347[(3'h4):(1'h1)]) >> ($signed((&reg335)) && $unsigned(((reg381 ?
                      reg374 : (8'ha3)) ?
                  (wire324 ? wire328 : reg337) : reg371))));
              reg388 <= {{(~^reg366), $unsigned((~|wire330))},
                  wire330[(3'h4):(1'h1)]};
            end
          else
            begin
              reg384 <= ((reg355 << reg366[(2'h3):(2'h3)]) ~^ reg331);
            end
          reg389 <= reg384;
          reg390 <= (~$signed(reg377[(3'h6):(1'h0)]));
        end
      else
        begin
          if (wire324)
            begin
              reg380 <= $signed($signed({{(reg326 ? (8'h9d) : wire324),
                      (^reg340)}}));
              reg381 <= $unsigned($unsigned(reg375[(5'h10):(4'he)]));
              reg382 <= ((~&(~$unsigned($signed(reg372)))) != (~&(8'hbf)));
            end
          else
            begin
              reg380 <= reg382;
              reg381 <= reg337;
            end
          reg383 <= $signed(reg356[(2'h3):(1'h1)]);
          reg384 <= {(reg366 << reg327),
              $signed(($unsigned(((8'ha4) ^ wire344)) << (^{reg347,
                  (8'h9f)})))};
          reg385 <= reg357;
        end
    end
  assign wire391 = (reg327[(4'ha):(2'h2)] >>> ($signed(wire321[(4'hb):(4'h9)]) ?
                       ((+$signed(reg379)) ?
                           ((7'h40) ^ reg337[(3'h6):(1'h1)]) : {(wire343 ?
                                   reg386 : wire343),
                               $unsigned(reg361)}) : (&$signed(reg377))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module477  (y, clk, wire481, wire480, wire479, wire478);
  output wire [(32'h46d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire481;
  input wire signed [(5'h12):(1'h0)] wire480;
  input wire signed [(5'h11):(1'h0)] wire479;
  input wire [(3'h6):(1'h0)] wire478;
  wire [(4'ha):(1'h0)] wire683;
  wire signed [(5'h14):(1'h0)] wire649;
  reg [(5'h13):(1'h0)] reg648 = (1'h0);
  reg [(4'hb):(1'h0)] reg647 = (1'h0);
  reg [(4'hd):(1'h0)] reg646 = (1'h0);
  reg [(5'h11):(1'h0)] reg645 = (1'h0);
  reg [(4'he):(1'h0)] reg644 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg643 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg642 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg641 = (1'h0);
  reg [(4'hd):(1'h0)] reg640 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg639 = (1'h0);
  reg [(3'h5):(1'h0)] reg638 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg637 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg636 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg635 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg634 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg633 = (1'h0);
  reg signed [(4'he):(1'h0)] reg632 = (1'h0);
  reg [(4'hf):(1'h0)] reg631 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg630 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg629 = (1'h0);
  reg [(2'h3):(1'h0)] reg628 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg627 = (1'h0);
  reg [(4'hc):(1'h0)] reg626 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire625;
  reg signed [(3'h5):(1'h0)] reg624 = (1'h0);
  reg [(4'h9):(1'h0)] reg623 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg622 = (1'h0);
  reg [(4'h8):(1'h0)] reg621 = (1'h0);
  reg [(4'hc):(1'h0)] reg620 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire619;
  wire [(3'h4):(1'h0)] wire618;
  reg [(5'h15):(1'h0)] reg617 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg616 = (1'h0);
  reg [(4'hf):(1'h0)] reg615 = (1'h0);
  reg [(5'h15):(1'h0)] reg614 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg613 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg612 = (1'h0);
  reg [(4'hf):(1'h0)] reg611 = (1'h0);
  reg [(4'hc):(1'h0)] reg610 = (1'h0);
  reg [(5'h12):(1'h0)] reg609 = (1'h0);
  reg [(5'h10):(1'h0)] reg608 = (1'h0);
  reg [(2'h2):(1'h0)] reg607 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg606 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg605 = (1'h0);
  reg [(5'h15):(1'h0)] reg604 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg603 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg602 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg601 = (1'h0);
  reg [(4'h8):(1'h0)] reg600 = (1'h0);
  reg [(3'h6):(1'h0)] reg599 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg598 = (1'h0);
  reg [(4'h8):(1'h0)] reg597 = (1'h0);
  reg [(5'h13):(1'h0)] reg596 = (1'h0);
  reg [(4'hb):(1'h0)] reg595 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg594 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire592;
  wire [(4'h9):(1'h0)] wire550;
  wire [(5'h10):(1'h0)] wire548;
  reg signed [(2'h2):(1'h0)] reg513 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg512 = (1'h0);
  reg [(3'h4):(1'h0)] reg511 = (1'h0);
  reg [(5'h15):(1'h0)] reg510 = (1'h0);
  reg [(5'h14):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg508 = (1'h0);
  reg [(5'h14):(1'h0)] reg507 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg506 = (1'h0);
  reg [(4'ha):(1'h0)] reg505 = (1'h0);
  reg [(3'h6):(1'h0)] reg504 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg503 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg502 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg501 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg500 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg498 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg497 = (1'h0);
  reg [(5'h12):(1'h0)] reg496 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg495 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg494 = (1'h0);
  reg [(4'hf):(1'h0)] reg493 = (1'h0);
  reg [(4'he):(1'h0)] reg492 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg491 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg490 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg489 = (1'h0);
  reg [(5'h15):(1'h0)] reg488 = (1'h0);
  reg [(4'hb):(1'h0)] reg487 = (1'h0);
  reg [(4'ha):(1'h0)] reg486 = (1'h0);
  reg [(2'h2):(1'h0)] reg485 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg484 = (1'h0);
  reg [(4'hb):(1'h0)] reg483 = (1'h0);
  reg [(4'hb):(1'h0)] reg482 = (1'h0);
  assign y = {wire683,
                 wire649,
                 reg648,
                 reg647,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 reg642,
                 reg641,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 reg636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 wire625,
                 reg624,
                 reg623,
                 reg622,
                 reg621,
                 reg620,
                 wire619,
                 wire618,
                 reg617,
                 reg616,
                 reg615,
                 reg614,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 wire592,
                 wire550,
                 wire548,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 reg501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 reg491,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ({($unsigned({wire479,
              wire481[(1'h0):(1'h0)]}) & wire478[(3'h5):(3'h4)])})
        begin
          if (wire480[(3'h6):(3'h5)])
            begin
              reg482 <= (^~wire479[(1'h1):(1'h0)]);
              reg483 <= wire478;
            end
          else
            begin
              reg482 <= ($signed((^$unsigned($unsigned(wire481)))) >>> (wire480[(1'h0):(1'h0)] * (wire481 ?
                  (~(wire479 ? reg483 : (8'h9f))) : wire479)));
              reg483 <= ((8'h9e) ?
                  (8'hac) : {{reg482}, ((-reg482[(4'ha):(2'h3)]) == wire480)});
              reg484 <= ($signed(reg482[(4'h9):(3'h6)]) <<< ((($signed(wire478) * (wire478 ?
                  (8'hb2) : (8'hae))) >> wire480[(4'hc):(1'h1)]) >> {{(~^wire480)}}));
              reg485 <= (7'h43);
            end
          reg486 <= reg482[(1'h0):(1'h0)];
        end
      else
        begin
          reg482 <= $unsigned((reg483[(3'h7):(3'h7)] < ((~reg484[(1'h1):(1'h0)]) ?
              ({(7'h43), wire480} ?
                  $unsigned(reg485) : reg483) : reg482[(2'h2):(2'h2)])));
        end
      reg487 <= {(^~((|$signed(reg482)) ?
              ({wire481} ?
                  (wire480 ? reg486 : wire481) : (~|wire480)) : reg482))};
    end
  always
    @(posedge clk) begin
      reg488 <= (^({(wire481 ? wire481 : (reg486 ? reg482 : reg484))} ?
          ({$unsigned(reg484), (reg483 != wire478)} ?
              {(|wire481), wire481} : (7'h44)) : (8'hbf)));
      if ({$signed($signed((reg483 * (7'h42)))),
          (($signed(reg485) == $signed(reg483)) + wire480[(3'h6):(2'h2)])})
        begin
          if (reg486[(4'h8):(1'h0)])
            begin
              reg489 <= (~^{$unsigned((((8'hb5) ?
                      reg486 : reg488) > $signed(wire479))),
                  $signed(reg485)});
              reg490 <= $signed(reg484);
            end
          else
            begin
              reg489 <= {((8'hb8) && reg482[(3'h7):(2'h3)]),
                  {reg485, (+reg488)}};
              reg490 <= wire478;
            end
          reg491 <= {((^~(!wire480[(3'h7):(3'h4)])) ?
                  $unsigned($unsigned((reg487 | (8'ha5)))) : ((((8'hbe) ?
                          reg489 : wire479) ?
                      (wire480 && wire480) : $signed(reg489)) * ((^~(8'h9f)) ?
                      $unsigned(wire481) : (reg489 ? reg488 : wire481))))};
          reg492 <= reg491;
          reg493 <= $signed(reg490);
        end
      else
        begin
          reg489 <= $signed($unsigned((reg484 * $unsigned((reg487 ?
              reg488 : reg486)))));
          reg490 <= $unsigned((reg484 != $unsigned((reg493[(4'he):(4'h9)] - reg489))));
          if ((wire480 && $signed($unsigned(reg486))))
            begin
              reg491 <= $signed($unsigned($signed((!(~^(8'hb1))))));
              reg492 <= (~^($signed(reg488[(4'h8):(1'h1)]) < ($signed((~|wire478)) ?
                  $signed((reg484 ? reg487 : reg484)) : $signed((reg485 ?
                      wire480 : (8'hac))))));
            end
          else
            begin
              reg491 <= $signed(($signed($unsigned((wire478 <= reg484))) ?
                  $signed(reg489) : $unsigned(reg489)));
              reg492 <= ($unsigned($signed(reg483[(4'h9):(2'h2)])) ?
                  ({reg483, (wire481 || (~&reg489))} ?
                      $unsigned((~&{(8'haf),
                          reg489})) : {$unsigned($unsigned(reg487))}) : (reg488[(3'h5):(1'h1)] & $unsigned(reg485)));
              reg493 <= reg483;
              reg494 <= $unsigned(reg482);
              reg495 <= (+$signed($unsigned($signed($unsigned(reg482)))));
            end
          if ($signed($signed((8'had))))
            begin
              reg496 <= $signed($unsigned(($unsigned(wire480) == (^$signed(reg490)))));
              reg497 <= $signed(reg490[(2'h2):(2'h2)]);
              reg498 <= (reg494[(4'h8):(3'h4)] >= reg489[(4'hb):(1'h0)]);
            end
          else
            begin
              reg496 <= ($signed({(^~(&reg486)),
                      (-(reg497 ? wire478 : (8'h9f)))}) ?
                  ($signed((8'hb9)) ?
                      reg494[(3'h5):(3'h5)] : reg493[(4'hd):(3'h4)]) : ($unsigned(reg482[(4'ha):(3'h6)]) ?
                      ($unsigned((^reg489)) ?
                          ($unsigned((8'ha9)) >>> (reg494 ?
                              reg492 : reg498)) : $signed((&wire479))) : reg498));
              reg497 <= ((!(!$signed((wire478 ? reg493 : (8'ha6))))) ?
                  ($unsigned((^$signed(reg483))) >= $signed(reg497[(5'h10):(4'he)])) : ((((reg494 + reg488) <<< (reg493 ?
                          reg496 : reg487)) ?
                      reg496 : (reg495 ?
                          (reg490 >= reg495) : (&reg494))) >= {(|reg495[(3'h5):(1'h1)])}));
            end
        end
      reg499 <= (({$signed($signed(reg490)),
              $unsigned($unsigned(reg483))} == reg491) ?
          reg489 : $signed(reg485[(1'h1):(1'h0)]));
      if (($unsigned($signed({{(8'hac)}})) << (^reg487)))
        begin
          if (((+$signed(((reg488 > reg496) ?
                  (reg498 ^ wire481) : (reg499 ^ (8'hbf))))) ?
              $unsigned((!$signed(reg484[(1'h0):(1'h0)]))) : (!($unsigned($signed(reg484)) < (~&(reg486 ?
                  reg491 : wire479))))))
            begin
              reg500 <= reg489;
              reg501 <= $signed({reg500});
              reg502 <= (-reg486);
              reg503 <= (reg500[(4'hb):(4'hb)] ?
                  (^~(8'hb7)) : $unsigned(wire481));
            end
          else
            begin
              reg500 <= $signed(({reg492[(4'hb):(3'h7)],
                  {reg494,
                      $signed((8'hac))}} * (^~$signed(reg492[(2'h3):(1'h0)]))));
              reg501 <= ({reg503,
                      {(((8'ha1) ? reg486 : reg483) ^ $unsigned(reg485)),
                          reg483}} ?
                  $unsigned(reg482) : $unsigned(reg489));
            end
          reg504 <= reg494[(4'h8):(3'h6)];
          if (($unsigned($unsigned(reg487)) ?
              $unsigned(($unsigned((wire481 ?
                  reg498 : reg485)) << (~^reg490[(1'h1):(1'h0)]))) : (8'ha8)))
            begin
              reg505 <= reg488[(3'h5):(3'h5)];
            end
          else
            begin
              reg505 <= ((~&reg500[(5'h12):(3'h6)]) >= $signed((((wire481 ?
                      reg484 : reg505) < (reg490 ? reg496 : reg494)) ?
                  ((reg485 ? reg505 : reg490) ?
                      $signed(wire479) : {wire479,
                          reg486}) : $signed((!reg493)))));
              reg506 <= (+wire481);
              reg507 <= reg486;
              reg508 <= ($unsigned(reg491) - (~^wire478));
            end
          if ((+{{reg508[(1'h0):(1'h0)]}}))
            begin
              reg509 <= reg483[(4'hb):(4'ha)];
              reg510 <= {$signed(reg487[(1'h1):(1'h1)])};
              reg511 <= reg510[(5'h13):(1'h1)];
              reg512 <= $unsigned($unsigned($unsigned(($unsigned((8'ha3)) ?
                  reg491[(4'h9):(3'h6)] : reg485[(1'h1):(1'h1)]))));
              reg513 <= ($signed(reg489) >= ($unsigned((((8'hac) ?
                          reg495 : reg506) ?
                      $unsigned((8'hba)) : reg510[(3'h4):(3'h4)])) ?
                  $signed((reg495 & (^~reg485))) : (~&(((8'ha9) | (8'ha6)) * reg504[(1'h1):(1'h1)]))));
            end
          else
            begin
              reg509 <= ((reg498 ?
                  ($signed($unsigned(reg499)) ?
                      reg488 : reg491) : (^~(~$unsigned(reg508)))) >= {(~|$signed((reg506 ?
                      reg487 : wire481)))});
              reg510 <= $signed(((^~(~^$unsigned(reg499))) ?
                  reg513 : {(^~(reg502 + reg484)), (8'had)}));
              reg511 <= (~&reg487[(2'h3):(1'h1)]);
              reg512 <= reg497;
              reg513 <= (!$signed((^~reg488)));
            end
        end
      else
        begin
          reg500 <= $signed((^$signed((~^((8'ha9) && reg498)))));
          if (({((7'h42) <= reg504)} ?
              (-(+$signed((~&reg513)))) : $signed(wire480)))
            begin
              reg501 <= reg487;
            end
          else
            begin
              reg501 <= reg488;
              reg502 <= {($signed(($signed((8'hbf)) | reg500[(4'h9):(4'h8)])) >>> (~|reg513)),
                  ($signed((|(reg504 ? reg506 : reg488))) ?
                      (|(8'ha7)) : ($signed(reg501[(5'h11):(5'h10)]) >> $signed((!reg500))))};
            end
          reg503 <= $unsigned(reg485);
          reg504 <= reg507;
        end
    end
  module514 modinst549 (wire548, clk, reg489, reg498, reg507, wire481);
  assign wire550 = $unsigned($unsigned($unsigned((&(reg482 >>> reg487)))));
  module551 modinst593 (.y(wire592), .wire553(reg502), .wire555(reg496), .clk(clk), .wire554(reg498), .wire552(reg488));
  always
    @(posedge clk) begin
      reg594 <= (wire548[(2'h3):(1'h0)] ?
          (reg502 ?
              (7'h41) : $signed({(8'ha6)})) : $unsigned(reg488[(3'h4):(1'h0)]));
      reg595 <= (~^$unsigned((-(|(reg496 <= wire592)))));
      if (reg513)
        begin
          reg596 <= {$unsigned(wire481[(5'h11):(4'h9)])};
        end
      else
        begin
          if (reg595[(4'h9):(4'h9)])
            begin
              reg596 <= reg596;
              reg597 <= $signed((($signed((wire550 + reg491)) | (|(reg490 ?
                      reg494 : reg485))) ?
                  $unsigned({(reg496 | reg486),
                      $unsigned(reg498)}) : $signed(reg511)));
              reg598 <= ($unsigned(({reg512, reg487[(3'h7):(2'h2)]} ?
                      $unsigned($signed(reg492)) : $signed(reg494))) ?
                  ($unsigned((|reg498[(4'h9):(3'h7)])) ^~ reg489[(4'h9):(4'h9)]) : (reg596 != $signed(reg597[(1'h1):(1'h0)])));
            end
          else
            begin
              reg596 <= $signed(reg598);
              reg597 <= (+reg489[(3'h7):(1'h0)]);
              reg598 <= (^$signed(($unsigned(reg506) ^~ ({reg497, reg498} ?
                  (~&reg495) : (wire480 && reg488)))));
              reg599 <= ($unsigned(((~&((8'haa) ^~ reg512)) ?
                      reg510 : $unsigned(((8'hbc) ? (8'hbd) : reg500)))) ?
                  ($unsigned(((reg492 ? reg595 : reg510) ?
                          (^~reg488) : (reg594 - reg499))) ?
                      reg485 : $signed($unsigned((reg598 ?
                          reg508 : reg492)))) : $unsigned($unsigned(reg503[(1'h0):(1'h0)])));
              reg600 <= reg598[(4'hc):(4'h8)];
            end
          reg601 <= ($signed($signed((reg594 >>> (8'hae)))) ?
              (reg489 | $unsigned(($signed((8'hac)) + $unsigned(reg500)))) : ((~(&reg508[(3'h6):(2'h3)])) ?
                  (wire592 >> ($signed(reg509) << (8'ha9))) : (^(reg511 <= (reg499 | reg488)))));
          if ((~($unsigned({((8'hb6) != reg509), (reg507 << reg512)}) ?
              $signed($unsigned({reg508})) : (^~$signed($signed(wire548))))))
            begin
              reg602 <= (~&($unsigned({$unsigned(wire478),
                  {reg482, reg598}}) || ((^$unsigned(reg485)) ?
                  (~reg596) : {reg486[(3'h6):(3'h4)]})));
              reg603 <= (-(8'had));
              reg604 <= $signed((8'hb5));
              reg605 <= {$unsigned((~|$signed(reg505))),
                  {$signed($unsigned((wire550 ? reg499 : reg513)))}};
            end
          else
            begin
              reg602 <= (~&reg604);
              reg603 <= {reg603};
              reg604 <= reg506[(3'h4):(3'h4)];
              reg605 <= reg497[(5'h13):(1'h1)];
            end
          reg606 <= $unsigned((($signed(reg484[(2'h2):(1'h1)]) ?
              $signed({(8'ha0), reg602}) : reg602[(3'h4):(2'h3)]) << wire480));
          reg607 <= wire479;
        end
      if ({((|reg488) << reg504[(1'h0):(1'h0)]),
          $unsigned(($unsigned((-reg494)) ~^ ($unsigned(wire479) | (reg493 ?
              (8'h9c) : reg505))))})
        begin
          reg608 <= ((+$unsigned((~wire480[(2'h2):(1'h1)]))) ?
              (($unsigned(reg485[(2'h2):(2'h2)]) - $unsigned(reg498)) ?
                  ($signed((reg600 ~^ wire481)) ?
                      reg508 : reg503[(3'h7):(3'h7)]) : (8'h9d)) : {$unsigned((+(reg490 ?
                      reg508 : reg498))),
                  $signed(reg483[(1'h0):(1'h0)])});
          reg609 <= (($signed(($signed(reg505) >>> reg511)) ^ $signed({reg600[(3'h4):(2'h3)],
                  $signed(reg510)})) ?
              wire478[(3'h6):(1'h0)] : ($unsigned(($unsigned(reg598) ?
                  {reg596, reg512} : $signed(reg489))) | $signed(((~^reg605) ?
                  (+wire481) : (^reg594)))));
          reg610 <= (reg509[(4'ha):(2'h2)] ?
              {(8'ha2)} : wire481[(3'h7):(1'h0)]);
        end
      else
        begin
          reg608 <= (~|wire478[(2'h2):(1'h1)]);
          reg609 <= $signed((reg486[(1'h1):(1'h1)] ?
              reg512[(3'h7):(3'h7)] : ({(~&(8'ha9)),
                  (+reg511)} <<< (^~(~^reg595)))));
          if (($signed(($signed((reg491 ? (8'hb9) : reg502)) ?
              (8'hb8) : reg605)) >= $unsigned(((reg504[(1'h1):(1'h0)] ?
                  (^reg492) : {reg492, (7'h41)}) ?
              reg506[(3'h7):(3'h5)] : ({reg488} ?
                  (reg493 ? (8'haa) : reg595) : (|reg485))))))
            begin
              reg610 <= (reg493[(4'h9):(3'h5)] | (reg610 >> reg491[(3'h7):(3'h5)]));
              reg611 <= ((7'h43) ?
                  ((({wire478, reg484} ?
                          {reg490, (8'ha3)} : $signed(reg489)) | (&(reg496 ?
                          (8'h9f) : reg511))) ?
                      $signed(reg492) : $signed(((^~reg609) ?
                          {reg490,
                              reg513} : $signed(reg482)))) : $signed((~&reg604)));
              reg612 <= $signed(((8'hae) ?
                  (reg508[(4'h8):(2'h2)] && $unsigned(((8'hbe) | reg509))) : (-(~$signed(reg483)))));
            end
          else
            begin
              reg610 <= (|reg484[(2'h2):(2'h2)]);
              reg611 <= ($signed((wire481[(4'hf):(4'ha)] << reg603)) ?
                  (&(~^(&reg594[(1'h1):(1'h0)]))) : reg504);
              reg612 <= reg608[(3'h5):(1'h0)];
            end
          if ($unsigned(reg487[(4'ha):(3'h7)]))
            begin
              reg613 <= reg599[(2'h2):(2'h2)];
              reg614 <= (~$unsigned($unsigned(reg504[(3'h6):(3'h6)])));
              reg615 <= reg483;
              reg616 <= (-$unsigned(({reg505, $signed(wire480)} ?
                  ($signed(reg508) && reg596) : $signed((reg506 && reg509)))));
              reg617 <= $unsigned((($signed((reg508 >= reg486)) <= reg596) <<< (7'h43)));
            end
          else
            begin
              reg613 <= reg504;
              reg614 <= (!reg488);
              reg615 <= (reg494 ?
                  reg600 : ({reg492[(3'h5):(3'h4)]} ?
                      (!((8'h9c) ?
                          reg484 : $unsigned(reg490))) : ($unsigned({(7'h44),
                          wire481}) & {(^~(8'hac))})));
            end
        end
    end
  assign wire618 = {$signed(((~^$signed(reg501)) ?
                           ({wire548} ?
                               (reg487 ? reg489 : reg599) : ((8'ha3) ?
                                   reg506 : reg495)) : reg607)),
                       ($unsigned(reg493[(3'h5):(1'h1)]) ?
                           reg511[(3'h4):(3'h4)] : (reg596[(3'h5):(3'h4)] ~^ ((reg492 ?
                               wire478 : (8'hb5)) < $unsigned(reg606))))};
  assign wire619 = (((($signed(reg502) + (^(8'hbd))) > wire550[(3'h7):(2'h3)]) < $unsigned(reg604)) >= (~^$unsigned(($signed(wire480) ?
                       {reg613, wire548} : $signed(reg501)))));
  always
    @(posedge clk) begin
      reg620 <= ($unsigned(($unsigned((reg505 ?
          reg489 : (8'hac))) | ($signed(reg509) ?
          (reg614 ?
              wire618 : wire478) : (reg484 ^~ (8'hb6))))) != (reg485[(1'h1):(1'h1)] ?
          ({(reg614 == wire481), {reg614}} ?
              (&{wire619}) : ((reg594 ? reg614 : reg599) ?
                  $unsigned((8'hb5)) : $signed(wire550))) : $unsigned({(reg489 + reg494)})));
      reg621 <= (!$unsigned({$signed(reg482[(2'h2):(2'h2)]),
          $unsigned({(8'hba), reg497})}));
      reg622 <= reg498[(3'h4):(2'h3)];
      reg623 <= $unsigned(wire480);
      reg624 <= $unsigned(((~&(wire479[(4'hd):(4'ha)] ?
              reg612 : $signed(reg616))) ?
          {$unsigned((~^(8'ha8))),
              $signed($unsigned(reg494))} : $unsigned($signed($unsigned((7'h42))))));
    end
  assign wire625 = $unsigned((^~reg594));
  always
    @(posedge clk) begin
      reg626 <= (^~(^wire625[(1'h1):(1'h0)]));
      if ($unsigned(({$signed({(8'ha5), reg626}),
          ($signed((8'ha2)) >> reg611)} >= (~wire625[(3'h5):(3'h5)]))))
        begin
          reg627 <= reg511;
          reg628 <= (|wire548[(3'h5):(3'h5)]);
        end
      else
        begin
          if ((((~&(reg596[(4'hc):(1'h0)] ?
                      (reg492 < reg597) : (reg628 <= reg610))) ?
                  reg492[(1'h0):(1'h0)] : {(^~$unsigned(wire592))}) ?
              reg594 : $signed(reg594)))
            begin
              reg627 <= {reg509[(1'h1):(1'h1)],
                  {reg616,
                      (((reg513 ? reg495 : reg624) ?
                              $signed(reg626) : (-reg498)) ?
                          reg503 : reg611)}};
              reg628 <= (+(-((^$unsigned(reg606)) ?
                  reg623[(2'h3):(1'h0)] : reg598)));
            end
          else
            begin
              reg627 <= ($signed(reg606) & $unsigned($unsigned($unsigned((-reg602)))));
            end
          reg629 <= (^$unsigned((!{(wire618 ? reg622 : reg599), reg503})));
          if ($unsigned($unsigned(reg615[(4'ha):(1'h0)])))
            begin
              reg630 <= reg602;
              reg631 <= reg606;
            end
          else
            begin
              reg630 <= reg607[(1'h0):(1'h0)];
              reg631 <= $unsigned(reg615[(3'h5):(3'h5)]);
            end
          if ({reg617})
            begin
              reg632 <= reg601[(1'h1):(1'h1)];
              reg633 <= (-(((~^(reg491 <= reg628)) ?
                  ({reg612, reg510} ?
                      reg493 : (reg606 == reg482)) : (~reg631[(2'h2):(2'h2)])) > (((reg623 ?
                      wire479 : reg612) ?
                  (reg487 || reg508) : $signed(reg616)) <= reg609[(4'h9):(4'h9)])));
              reg634 <= (reg613 ?
                  (!({wire478[(1'h0):(1'h0)]} & reg633)) : {(reg633 > reg630[(4'hd):(3'h4)])});
              reg635 <= reg595;
              reg636 <= ($unsigned(($signed($signed(reg483)) ?
                      {(&reg511)} : reg628)) ?
                  (^{reg598[(4'h9):(3'h5)],
                      ($unsigned(reg600) ?
                          reg512[(1'h1):(1'h0)] : $signed(reg604))}) : reg603[(3'h4):(1'h1)]);
            end
          else
            begin
              reg632 <= wire618;
              reg633 <= reg617[(4'ha):(1'h1)];
              reg634 <= (~^(($signed((reg501 ? reg488 : reg495)) ?
                      reg634 : {(reg607 ? reg605 : (8'ha7)), $signed(reg598)}) ?
                  reg510 : (reg485 ?
                      $unsigned((-(8'ha0))) : $unsigned({reg486}))));
              reg635 <= $signed(((8'h9d) ^ $signed(reg624[(1'h0):(1'h0)])));
            end
          if ({(!$signed(((reg596 ?
                  reg622 : wire480) != reg489[(1'h0):(1'h0)]))),
              reg513})
            begin
              reg637 <= (((~&((reg504 ?
                  reg612 : reg483) == $unsigned(reg628))) ^ reg483[(4'ha):(1'h1)]) - ($signed({$signed(reg595)}) >> (wire619 ?
                  $unsigned(wire479[(3'h7):(1'h0)]) : (8'ha7))));
              reg638 <= (~|$signed((^$signed((wire619 ? (8'hb5) : reg491)))));
            end
          else
            begin
              reg637 <= $unsigned($signed((((reg507 ?
                      reg632 : reg492) ^~ (|reg600)) ?
                  $unsigned((reg614 + wire550)) : (~^wire592[(4'h9):(1'h1)]))));
              reg638 <= {reg485[(1'h0):(1'h0)]};
            end
        end
      reg639 <= (^($signed((~&$unsigned(reg600))) ?
          $signed(reg492) : $unsigned(($unsigned(wire478) ?
              (wire479 ? (8'hac) : (8'hba)) : (~^reg501)))));
      reg640 <= $unsigned((&((-(8'ha0)) ?
          (reg631[(3'h6):(3'h5)] < reg614[(3'h7):(3'h6)]) : (~^{reg594,
              reg631}))));
      if ((^reg484[(1'h1):(1'h0)]))
        begin
          reg641 <= $unsigned(wire625);
          if ($signed(reg482))
            begin
              reg642 <= reg603;
            end
          else
            begin
              reg642 <= {(reg482 ~^ $signed(reg597[(4'h8):(2'h3)])), reg615};
              reg643 <= ({$unsigned(($signed(reg497) ?
                      reg632 : reg640[(4'hd):(3'h6)])),
                  $unsigned({$unsigned(reg594)})} * ($unsigned(((8'hae) >>> (reg512 << reg629))) <<< reg630));
              reg644 <= (((reg613 + reg499[(1'h1):(1'h1)]) ~^ (|{reg620})) ~^ (reg500[(4'ha):(2'h2)] ?
                  (($signed(reg603) <= $unsigned((7'h42))) == (~&$signed(wire619))) : $unsigned(((~^(8'hbe)) ?
                      reg492 : wire618[(2'h3):(2'h2)]))));
              reg645 <= $unsigned((($unsigned(((8'hba) ?
                      (8'ha1) : reg603)) && ((8'hbb) ?
                      reg629 : $unsigned(reg620))) ?
                  $unsigned($unsigned($unsigned(reg486))) : reg631));
            end
          reg646 <= reg494;
          reg647 <= {$unsigned({$signed($unsigned(reg496))})};
          reg648 <= $unsigned(reg607[(2'h2):(1'h0)]);
        end
      else
        begin
          if (wire625[(2'h3):(2'h2)])
            begin
              reg641 <= (|((((reg633 ? reg631 : reg604) ?
                      {reg627} : reg489) > $signed($unsigned(reg594))) ?
                  $signed(((|reg604) ?
                      (reg613 > reg493) : reg492[(3'h7):(2'h3)])) : (7'h42)));
            end
          else
            begin
              reg641 <= $unsigned(($signed(((reg630 ? (8'hac) : reg616) ?
                      reg631[(4'hf):(2'h3)] : reg488)) ?
                  reg612 : (({reg611} ?
                          (reg498 ? reg630 : reg613) : $unsigned(reg634)) ?
                      reg608[(1'h0):(1'h0)] : ((reg637 >> reg601) + $unsigned(reg614)))));
              reg642 <= ((reg483[(4'h8):(2'h2)] ?
                      (($signed(reg635) ~^ (reg623 + reg492)) + {reg621[(1'h0):(1'h0)],
                          (reg489 ?
                              reg501 : reg645)}) : {($signed(reg614) - $signed((7'h43))),
                          (8'hbd)}) ?
                  (^~(&(-(reg648 ?
                      reg497 : reg611)))) : $signed(($signed($signed(reg627)) | reg630)));
              reg643 <= {((!$signed((&reg602))) & ((&$unsigned(reg508)) >>> (wire481 ?
                      (^(8'hb2)) : $unsigned(reg604)))),
                  reg648};
              reg644 <= reg601;
            end
          reg645 <= {{{$unsigned(((8'ha0) ? reg612 : reg646))}, reg512}};
        end
    end
  assign wire649 = (+wire480[(3'h5):(3'h5)]);
  module650 modinst684 (wire683, clk, reg488, reg634, reg505, reg509);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module650
#( parameter param681 = ((^~(-((~^(8'hb2)) ? {(8'ha3), (8'hb2)} : ((8'hb9) > (8'ha2))))) ? (((^((8'hb8) ? (8'hbb) : (8'hb0))) || (^~{(8'ha9)})) << (|({(8'hb8), (8'had)} ? ((8'ha4) <= (8'ha6)) : ((8'hac) || (7'h41))))) : ((~&((-(8'h9c)) ? ((8'haa) ? (8'h9f) : (8'hbd)) : (-(8'hb9)))) ? ((~&((8'hb9) ? (8'had) : (8'ha8))) ? (~^(~|(8'hb3))) : (^(~|(8'hb7)))) : {(((8'ha0) ? (8'hb6) : (8'ha1)) ? ((8'ha2) ? (8'haa) : (8'hb2)) : (8'hac)), (~((8'had) ? (8'hb8) : (8'hac)))}))
, parameter param682 = (((((param681 ? (8'haf) : param681) != (param681 >>> (8'hbc))) * param681) ? param681 : (((~|param681) ? (param681 + param681) : (param681 ? param681 : param681)) ? param681 : {param681})) >= ({(param681 ? (param681 ? param681 : param681) : (+param681))} - {(~^(~param681))})) )
(y, clk, wire654, wire653, wire652, wire651);
  output wire [(32'h130):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire654;
  input wire [(2'h3):(1'h0)] wire653;
  input wire signed [(4'ha):(1'h0)] wire652;
  input wire [(5'h14):(1'h0)] wire651;
  reg signed [(5'h11):(1'h0)] reg680 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg679 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg678 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg677 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg676 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg675 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg674 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg673 = (1'h0);
  reg [(4'hb):(1'h0)] reg672 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg671 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg670 = (1'h0);
  reg [(5'h13):(1'h0)] reg669 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg668 = (1'h0);
  reg [(3'h7):(1'h0)] reg667 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg666 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg664 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg663 = (1'h0);
  reg [(3'h5):(1'h0)] reg662 = (1'h0);
  reg [(4'hd):(1'h0)] reg661 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg660 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg659 = (1'h0);
  reg [(5'h13):(1'h0)] reg658 = (1'h0);
  wire [(2'h3):(1'h0)] wire657;
  wire signed [(5'h14):(1'h0)] wire656;
  wire signed [(3'h4):(1'h0)] wire655;
  assign y = {reg680,
                 reg679,
                 reg678,
                 reg677,
                 reg676,
                 reg675,
                 reg674,
                 reg673,
                 reg672,
                 reg671,
                 reg670,
                 reg669,
                 reg668,
                 reg667,
                 reg666,
                 reg665,
                 reg664,
                 reg663,
                 reg662,
                 reg661,
                 reg660,
                 reg659,
                 reg658,
                 wire657,
                 wire656,
                 wire655,
                 (1'h0)};
  assign wire655 = $unsigned(($unsigned((^~{wire654})) << {wire654}));
  assign wire656 = wire654;
  assign wire657 = $unsigned($signed($unsigned($unsigned({wire652}))));
  always
    @(posedge clk) begin
      if ((((-($unsigned(wire653) == (wire656 ~^ wire654))) >= {wire657,
          wire654[(3'h6):(2'h2)]}) + {(|(wire651 || {wire656, (8'hb6)}))}))
        begin
          reg658 <= $unsigned(($signed(({wire653, wire652} < wire651)) ?
              (!wire656[(4'he):(3'h7)]) : {wire653[(2'h2):(2'h2)],
                  (wire653 ^ (~&wire654))}));
        end
      else
        begin
          if ((wire653 == (~&(^~$signed(wire657[(2'h3):(1'h0)])))))
            begin
              reg658 <= $unsigned(wire656[(1'h1):(1'h1)]);
              reg659 <= (~wire651[(4'hb):(3'h5)]);
            end
          else
            begin
              reg658 <= (((wire656 ? $signed((wire655 - reg658)) : reg659) ?
                  (|(&$signed(wire653))) : reg659) <= wire653[(2'h2):(1'h0)]);
              reg659 <= ((8'ha9) ?
                  reg659[(4'h9):(3'h4)] : ($signed((8'hba)) ?
                      wire653 : wire653));
              reg660 <= (+$signed($signed((wire654[(3'h4):(1'h0)] >>> (-wire655)))));
              reg661 <= (wire656[(3'h4):(2'h2)] ?
                  wire652 : $signed($signed((^{(8'hbc)}))));
              reg662 <= wire653;
            end
          if ({(+(-wire652[(3'h5):(2'h2)]))})
            begin
              reg663 <= (reg658 ?
                  ((8'hae) <= (((wire653 ? (8'ha4) : wire651) ?
                      (reg661 <= reg658) : $signed(reg658)) ^~ wire657)) : $unsigned(($unsigned($unsigned(wire655)) ?
                      (^wire657[(1'h0):(1'h0)]) : wire656)));
              reg664 <= (reg659[(3'h4):(1'h1)] - {{$unsigned($signed(wire653)),
                      {{wire653}}}});
              reg665 <= reg663;
              reg666 <= $unsigned((^$signed($unsigned((|reg659)))));
            end
          else
            begin
              reg663 <= reg662;
              reg664 <= ({$unsigned(($signed(wire652) ?
                          {reg665, wire657} : $signed(wire656)))} ?
                  wire652 : {reg664[(1'h0):(1'h0)], wire651});
              reg665 <= (^~wire652);
              reg666 <= (&reg660);
            end
          reg667 <= {{$signed(reg659[(2'h3):(2'h2)]), wire655}};
        end
      if ((&(((&(wire651 < reg660)) ? $unsigned({reg667}) : reg662) ?
          {((reg661 ? reg660 : wire657) ?
                  (+reg658) : (wire654 ? wire657 : wire654))} : ((7'h44) ?
              ({reg662, wire652} ?
                  $unsigned(reg662) : $signed((8'hac))) : $signed((reg665 ^~ wire654))))))
        begin
          if ($unsigned((8'ha0)))
            begin
              reg668 <= (~$signed($signed((|reg660))));
            end
          else
            begin
              reg668 <= $signed($unsigned((8'hbb)));
              reg669 <= $unsigned(wire654);
            end
          if ((~reg664[(1'h0):(1'h0)]))
            begin
              reg670 <= wire654;
              reg671 <= wire653;
              reg672 <= wire657;
              reg673 <= (8'hbe);
              reg674 <= ((+reg670[(4'hd):(3'h6)]) ?
                  $unsigned(reg667) : {($signed(wire651[(4'he):(4'h9)]) ?
                          wire655[(1'h1):(1'h0)] : ((8'hb4) == ((8'hb5) - (8'ha6))))});
            end
          else
            begin
              reg670 <= (8'hbb);
              reg671 <= (reg659 != reg671);
              reg672 <= reg666;
              reg673 <= (8'hbc);
            end
          if ((8'hb8))
            begin
              reg675 <= wire652;
              reg676 <= ((reg673[(1'h1):(1'h0)] ?
                  (~reg663) : $unsigned((~^$unsigned(reg661)))) && $signed((~^$signed($unsigned(reg662)))));
              reg677 <= ($unsigned($signed((8'hb0))) == $signed({(~&reg667),
                  reg667}));
              reg678 <= (reg666 == {((~^(reg671 ?
                      reg667 : reg671)) | (+(reg676 ? reg672 : wire653)))});
            end
          else
            begin
              reg675 <= ((+(reg662 << (-(reg678 != (8'haf))))) ?
                  (wire654[(5'h12):(2'h2)] <= $signed(reg673[(2'h3):(2'h2)])) : (wire653 ?
                      {(~$unsigned(wire652)),
                          $unsigned(reg670[(3'h6):(3'h5)])} : (!(~&reg663[(1'h0):(1'h0)]))));
              reg676 <= reg668[(1'h1):(1'h1)];
              reg677 <= (wire653[(2'h2):(1'h0)] ?
                  (~|(wire657[(2'h3):(2'h3)] ~^ $unsigned((8'hb1)))) : (!(((reg678 ?
                      reg667 : wire652) == reg674) >> $signed(reg660[(1'h0):(1'h0)]))));
              reg678 <= (&(^~(($unsigned(reg659) ?
                      (wire656 ? reg670 : reg674) : (reg665 ?
                          (7'h41) : reg674)) ?
                  (reg677 ?
                      reg664 : $signed(reg661)) : reg673[(2'h3):(2'h3)])));
              reg679 <= ((-$signed($signed(reg664))) ?
                  $unsigned($signed((~^reg663))) : reg666[(4'h8):(3'h4)]);
            end
        end
      else
        begin
          reg668 <= reg675;
          reg669 <= ((~|((reg674[(4'h8):(3'h7)] ?
                  $signed(wire652) : (reg671 ? (8'hbd) : reg675)) ?
              {wire653, reg672} : ($unsigned(reg665) ?
                  (reg678 ? reg673 : reg668) : {reg676,
                      reg679}))) <<< ($signed($unsigned($unsigned(reg669))) ?
              reg669[(5'h13):(3'h7)] : $signed($signed((8'had)))));
          if (reg665)
            begin
              reg670 <= $signed($unsigned(reg677));
            end
          else
            begin
              reg670 <= $signed($unsigned(wire654));
              reg671 <= (($signed(wire651[(2'h2):(1'h1)]) ?
                  ((+$signed(wire651)) ?
                      reg659 : wire654[(4'h9):(2'h3)]) : ((~^reg671[(4'hc):(1'h0)]) <= reg678)) && wire654[(5'h14):(3'h6)]);
              reg672 <= (+$signed((^~wire656)));
              reg673 <= $unsigned(reg678[(1'h0):(1'h0)]);
            end
          reg674 <= ((^(8'hb1)) >> (-reg674));
        end
      reg680 <= reg672[(3'h4):(2'h2)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module551
#( parameter param590 = (~&((({(7'h44)} ? ((8'h9c) ? (8'hb3) : (8'hac)) : ((8'hba) >> (7'h42))) ? ((~^(8'ha6)) ? ((8'haa) ? (8'hbc) : (8'hb0)) : ((8'hba) ? (8'hba) : (8'hb5))) : (~^(~(8'hb7)))) << (!(((8'hb2) == (8'h9f)) ^ (!(8'h9c))))))
, parameter param591 = ({(~{(param590 + (8'h9c)), ((8'hb9) || param590)})} ? (&(8'hab)) : ({(((7'h44) ? param590 : param590) <= (param590 >= param590))} >> param590)) )
(y, clk, wire555, wire554, wire553, wire552);
  output wire [(32'h177):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire555;
  input wire signed [(3'h4):(1'h0)] wire554;
  input wire signed [(2'h2):(1'h0)] wire553;
  input wire [(2'h2):(1'h0)] wire552;
  wire [(5'h15):(1'h0)] wire589;
  wire signed [(5'h13):(1'h0)] wire588;
  wire signed [(4'h8):(1'h0)] wire587;
  wire signed [(3'h6):(1'h0)] wire586;
  wire signed [(4'ha):(1'h0)] wire585;
  wire [(4'hf):(1'h0)] wire584;
  wire signed [(4'hc):(1'h0)] wire583;
  wire signed [(2'h3):(1'h0)] wire582;
  wire [(3'h6):(1'h0)] wire581;
  wire [(5'h12):(1'h0)] wire580;
  reg [(5'h10):(1'h0)] reg579 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg578 = (1'h0);
  reg [(5'h15):(1'h0)] reg577 = (1'h0);
  reg [(4'hf):(1'h0)] reg576 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg575 = (1'h0);
  reg [(4'hf):(1'h0)] reg574 = (1'h0);
  reg [(2'h2):(1'h0)] reg573 = (1'h0);
  reg [(3'h5):(1'h0)] reg572 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg571 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg570 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg569 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg568 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg567 = (1'h0);
  reg [(5'h10):(1'h0)] reg566 = (1'h0);
  reg [(5'h13):(1'h0)] reg565 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg564 = (1'h0);
  reg [(3'h5):(1'h0)] reg563 = (1'h0);
  reg [(3'h7):(1'h0)] reg562 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg561 = (1'h0);
  reg [(3'h4):(1'h0)] reg560 = (1'h0);
  reg [(5'h10):(1'h0)] reg559 = (1'h0);
  reg [(3'h7):(1'h0)] reg558 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire557;
  wire [(5'h11):(1'h0)] wire556;
  assign y = {wire589,
                 wire588,
                 wire587,
                 wire586,
                 wire585,
                 wire584,
                 wire583,
                 wire582,
                 wire581,
                 wire580,
                 reg579,
                 reg578,
                 reg577,
                 reg576,
                 reg575,
                 reg574,
                 reg573,
                 reg572,
                 reg571,
                 reg570,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 reg565,
                 reg564,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 reg558,
                 wire557,
                 wire556,
                 (1'h0)};
  assign wire556 = $signed($signed({{(^wire554)},
                       $signed($unsigned(wire555))}));
  assign wire557 = {{wire555[(3'h7):(1'h1)], $unsigned((~&(!wire556)))},
                       $signed(wire553[(2'h2):(1'h0)])};
  always
    @(posedge clk) begin
      if (wire553)
        begin
          if (wire556[(3'h6):(2'h3)])
            begin
              reg558 <= {{(-$signed((8'hb2))), wire556[(4'h8):(3'h4)]}};
              reg559 <= $unsigned(wire556[(4'ha):(2'h2)]);
              reg560 <= wire555;
            end
          else
            begin
              reg558 <= (+{$unsigned($signed($unsigned((8'h9d))))});
            end
          reg561 <= (wire553[(2'h2):(1'h0)] ?
              ({$signed((reg559 != reg560)),
                      ((|wire557) ? (8'hac) : (-wire557))} ?
                  $signed(($signed(wire555) ^~ $unsigned(wire555))) : {reg560}) : $signed(wire552));
          if ($unsigned($unsigned(($unsigned((^~wire552)) ?
              ((reg559 ? wire556 : reg559) <<< $unsigned(wire554)) : {(wire554 ?
                      wire552 : (8'hba)),
                  {wire554}}))))
            begin
              reg562 <= (reg560 ?
                  ($signed(reg558[(1'h1):(1'h1)]) ?
                      ({(wire553 ? (8'hb5) : reg561),
                          (~wire554)} | {(^wire553)}) : reg560) : (^~({(wire555 && wire557),
                      wire553[(1'h0):(1'h0)]} ^~ wire555[(2'h3):(2'h2)])));
              reg563 <= (reg558[(3'h6):(3'h5)] > {$signed($unsigned(((8'hb9) >= reg561)))});
              reg564 <= ($signed((reg558 ?
                      $unsigned((wire555 != wire556)) : (~^(wire552 ?
                          wire554 : reg561)))) ?
                  (8'had) : $unsigned({reg559[(5'h10):(2'h2)]}));
              reg565 <= ((-wire554[(2'h2):(2'h2)]) >> $signed($signed(($unsigned(wire553) ?
                  $unsigned(wire552) : (reg562 == reg558)))));
            end
          else
            begin
              reg562 <= wire554[(1'h1):(1'h1)];
            end
          reg566 <= ({{({wire553} < $unsigned(reg565)),
                  $signed($signed(wire553))},
              {$signed(((8'hb2) >>> (8'ha6)))}} ^ (~^reg560));
        end
      else
        begin
          reg558 <= ((&((~|(~|reg565)) ?
                  $unsigned((&reg561)) : reg561[(3'h5):(3'h5)])) ?
              ((^~((reg566 ? reg566 : (8'ha0)) * (reg560 ? reg561 : reg559))) ?
                  (~({wire553} * (~&reg563))) : reg558) : (|$signed($unsigned((reg558 >= wire556)))));
          reg559 <= reg566;
          reg560 <= $signed($signed(wire557));
        end
      if ((reg559 <<< ((~$signed((!wire552))) ?
          $unsigned(wire552[(2'h2):(1'h1)]) : $unsigned(((wire554 ?
                  reg564 : reg565) ?
              $signed(reg558) : {reg561})))))
        begin
          if (reg566[(5'h10):(1'h0)])
            begin
              reg567 <= (|(($unsigned((-reg565)) != {(8'hb1)}) & $signed((~^reg564))));
              reg568 <= {reg567};
              reg569 <= ($signed($signed(reg560)) && $signed({($signed(wire553) ^~ $unsigned((7'h40))),
                  reg561}));
              reg570 <= $signed(wire555[(3'h5):(1'h1)]);
            end
          else
            begin
              reg567 <= $unsigned(((reg564[(2'h2):(1'h0)] >> (~^$unsigned((8'ha0)))) * (wire553[(1'h0):(1'h0)] ?
                  reg563 : (8'hb3))));
            end
          reg571 <= wire556;
          if (reg562)
            begin
              reg572 <= {($signed(reg566) ?
                      ($unsigned((~|reg569)) ?
                          ($unsigned(wire552) ?
                              (wire556 ?
                                  reg563 : (8'hb9)) : wire555[(2'h2):(1'h0)]) : reg558[(3'h5):(1'h1)]) : wire553),
                  reg560[(2'h3):(1'h0)]};
              reg573 <= wire557[(4'he):(3'h6)];
              reg574 <= (reg559[(3'h4):(2'h3)] ?
                  (~&(($signed(reg571) ?
                      $unsigned((8'h9d)) : $signed(reg565)) > $unsigned(reg558[(3'h7):(3'h5)]))) : {{$signed((~reg560))},
                      reg564[(2'h2):(1'h0)]});
              reg575 <= {(+wire552[(1'h1):(1'h0)])};
            end
          else
            begin
              reg572 <= reg560;
              reg573 <= $unsigned(reg568);
              reg574 <= (reg560 ?
                  reg568[(1'h0):(1'h0)] : wire556[(4'hc):(1'h1)]);
              reg575 <= {reg566[(4'hf):(4'he)]};
            end
          reg576 <= $signed($signed(reg572[(2'h2):(1'h1)]));
          if ($signed($signed(({reg569} ?
              reg571 : ($signed((8'ha1)) ? reg564 : $unsigned(reg568))))))
            begin
              reg577 <= ($unsigned($signed(($unsigned(reg559) >= (reg571 ^ reg570)))) ?
                  (8'hbe) : reg575[(1'h0):(1'h0)]);
            end
          else
            begin
              reg577 <= wire554;
              reg578 <= $signed((reg567 ?
                  ((7'h43) || ((reg559 ? reg564 : reg576) && {reg577,
                      reg567})) : (reg577[(5'h12):(4'hf)] ?
                      (reg562[(3'h7):(3'h5)] ?
                          {(8'hb4), wire552} : (reg567 ?
                              reg564 : wire553)) : (~|reg572))));
              reg579 <= $signed((wire553[(1'h0):(1'h0)] ? (8'ha3) : wire552));
            end
        end
      else
        begin
          reg567 <= $signed((((reg579 >>> $unsigned(reg571)) ~^ ($signed(reg578) ?
                  $signed(wire555) : wire556)) ?
              ($unsigned((!reg573)) ?
                  ((wire556 ? wire557 : reg558) ?
                      {reg578} : $unsigned(wire553)) : (&(^~reg560))) : (~reg565)));
          if (((8'hb0) ?
              (-(~&reg558[(2'h3):(1'h1)])) : $signed($signed(((^reg579) ?
                  (-reg567) : reg560[(1'h1):(1'h0)])))))
            begin
              reg568 <= reg569;
              reg569 <= (-$signed((^wire555)));
              reg570 <= $unsigned({$unsigned(reg559)});
            end
          else
            begin
              reg568 <= ((|{((reg565 != (8'hbd)) ~^ wire557[(3'h6):(3'h4)]),
                      reg566}) ?
                  reg568 : reg578);
              reg569 <= $unsigned($signed({$unsigned((reg576 ?
                      (7'h41) : reg560))}));
            end
        end
    end
  assign wire580 = (reg566[(4'hb):(2'h3)] ?
                       {reg568} : (~|($signed({reg562}) || reg572)));
  assign wire581 = ((~&(+$unsigned((-(7'h43))))) == (((&reg577) != (|reg558[(1'h1):(1'h0)])) >> $signed(reg558)));
  assign wire582 = reg565[(1'h0):(1'h0)];
  assign wire583 = reg566[(4'h9):(4'h9)];
  assign wire584 = (8'had);
  assign wire585 = (($signed(reg574[(3'h6):(3'h4)]) && $unsigned($unsigned((+wire583)))) ?
                       (^(((reg564 ?
                               (8'hb0) : reg561) >= reg561[(1'h1):(1'h1)]) ?
                           (reg565[(3'h4):(2'h3)] ?
                               reg569 : reg561[(3'h5):(2'h3)]) : (!(wire580 - wire583)))) : wire555);
  assign wire586 = $unsigned(reg568);
  assign wire587 = ((7'h42) ?
                       {reg579,
                           (!(((8'hbc) >>> wire584) | {wire582,
                               (8'hb4)}))} : {$signed(($unsigned(reg572) ?
                               reg562 : (^wire557))),
                           (reg561[(3'h4):(2'h3)] ?
                               (~(reg559 ?
                                   reg567 : (8'hb8))) : $unsigned((reg575 ?
                                   wire554 : (8'h9c))))});
  assign wire588 = wire552;
  assign wire589 = $signed((-(7'h42)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module514  (y, clk, wire518, wire517, wire516, wire515);
  output wire [(32'h16f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire518;
  input wire [(5'h11):(1'h0)] wire517;
  input wire signed [(4'hc):(1'h0)] wire516;
  input wire [(5'h13):(1'h0)] wire515;
  wire signed [(4'hc):(1'h0)] wire547;
  wire signed [(4'ha):(1'h0)] wire546;
  wire [(3'h5):(1'h0)] wire545;
  wire [(3'h7):(1'h0)] wire544;
  reg signed [(4'h9):(1'h0)] reg543 = (1'h0);
  reg [(5'h11):(1'h0)] reg542 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg541 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg540 = (1'h0);
  reg [(4'hb):(1'h0)] reg539 = (1'h0);
  reg [(4'ha):(1'h0)] reg538 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg537 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg536 = (1'h0);
  reg [(5'h10):(1'h0)] reg535 = (1'h0);
  reg [(4'he):(1'h0)] reg534 = (1'h0);
  reg [(4'h8):(1'h0)] reg533 = (1'h0);
  reg [(4'he):(1'h0)] reg532 = (1'h0);
  reg [(4'he):(1'h0)] reg531 = (1'h0);
  reg [(3'h7):(1'h0)] reg530 = (1'h0);
  reg [(5'h14):(1'h0)] reg529 = (1'h0);
  reg [(4'hd):(1'h0)] reg528 = (1'h0);
  reg [(3'h7):(1'h0)] reg527 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg526 = (1'h0);
  reg [(5'h11):(1'h0)] reg525 = (1'h0);
  wire [(4'he):(1'h0)] wire524;
  reg signed [(4'h8):(1'h0)] reg523 = (1'h0);
  reg [(4'he):(1'h0)] reg522 = (1'h0);
  reg [(5'h14):(1'h0)] reg521 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg520 = (1'h0);
  wire [(4'hd):(1'h0)] wire519;
  assign y = {wire547,
                 wire546,
                 wire545,
                 wire544,
                 reg543,
                 reg542,
                 reg541,
                 reg540,
                 reg539,
                 reg538,
                 reg537,
                 reg536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 wire524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 wire519,
                 (1'h0)};
  assign wire519 = $unsigned(wire517[(1'h1):(1'h0)]);
  always
    @(posedge clk) begin
      reg520 <= $unsigned({{$signed({wire517})},
          (wire516[(2'h3):(2'h3)] ?
              $unsigned($unsigned(wire516)) : wire517[(2'h2):(2'h2)])});
      reg521 <= wire519;
      if (((|reg521[(4'ha):(2'h3)]) || ((+$unsigned((wire516 <= wire519))) ?
          $unsigned($signed((wire519 ?
              wire515 : wire517))) : ((reg520[(3'h6):(3'h5)] <<< $unsigned(reg521)) | $unsigned($unsigned((8'h9d)))))))
        begin
          reg522 <= ({(~|$signed((8'ha2))),
                  $unsigned(((wire515 ? wire517 : wire519) && (+wire515)))} ?
              {(wire518 ?
                      ($signed(wire517) ?
                          (&wire518) : $unsigned(wire515)) : reg521[(5'h14):(2'h2)])} : ($signed($signed((wire516 ?
                      reg521 : (8'hb9)))) ?
                  {$signed({wire519, (8'hab)}),
                      (wire515[(4'h8):(1'h0)] == $unsigned(wire519))} : $unsigned(((~wire518) ~^ {reg520}))));
        end
      else
        begin
          reg522 <= wire516;
        end
      reg523 <= (reg522 ?
          wire516[(2'h3):(1'h1)] : {$signed((|{wire516, wire517})),
              $unsigned(((8'hae) ? (^wire515) : {reg521, wire517}))});
    end
  assign wire524 = $unsigned(wire516);
  always
    @(posedge clk) begin
      if ($unsigned(($unsigned((&$unsigned(reg520))) ?
          ((8'ha9) ?
              $signed(wire518) : ((+reg520) || $signed(wire519))) : wire519[(4'hd):(4'h9)])))
        begin
          reg525 <= {{(^~({(8'hbf)} - (wire516 >>> wire517))),
                  $unsigned(reg523[(4'h8):(2'h3)])},
              (wire516 ?
                  $unsigned((wire524[(1'h1):(1'h1)] * {reg521})) : ((^~reg520) ~^ wire524[(2'h2):(2'h2)]))};
          reg526 <= (($unsigned(reg520) ?
              ((^(-wire516)) <<< (wire524 - $unsigned((7'h40)))) : (((reg525 ^ reg523) ?
                  $signed(wire524) : $unsigned(reg522)) & {(reg522 ?
                      wire518 : reg523),
                  $signed((8'h9c))})) < wire515[(3'h7):(3'h6)]);
        end
      else
        begin
          if ($signed(($signed($unsigned($unsigned(wire515))) && ($unsigned(reg522) > ((reg523 ?
                  wire519 : wire515) ?
              $signed(wire516) : (&reg520))))))
            begin
              reg525 <= wire519;
              reg526 <= reg521;
              reg527 <= $unsigned({((&$unsigned(wire516)) ?
                      (!wire515[(4'hd):(2'h2)]) : (~|(reg522 >= wire524)))});
            end
          else
            begin
              reg525 <= (8'ha8);
            end
        end
      reg528 <= $unsigned({(((wire519 ? reg523 : (8'h9c)) ?
                  (8'hbc) : $signed(reg525)) ?
              ((wire519 * (8'hba)) - $signed((8'hb9))) : $signed((~reg520)))});
      reg529 <= reg526;
    end
  always
    @(posedge clk) begin
      if ($signed({(-wire516), (reg520 ? wire517[(5'h10):(3'h5)] : reg521)}))
        begin
          if (reg522)
            begin
              reg530 <= $unsigned({reg526[(4'hf):(4'hd)],
                  ((8'haa) ?
                      reg527[(3'h5):(2'h3)] : $signed((reg528 & reg520)))});
              reg531 <= $unsigned(reg521);
              reg532 <= {(7'h44)};
              reg533 <= reg529[(3'h5):(3'h4)];
            end
          else
            begin
              reg530 <= (wire516 - reg523[(4'h8):(1'h0)]);
            end
          if (($signed(((~^$signed(wire518)) ?
                  reg522 : ($unsigned(reg532) ?
                      {reg528, reg528} : reg527[(3'h7):(1'h0)]))) ?
              reg528[(4'hc):(4'ha)] : ((({reg521} ?
                          $unsigned(reg529) : $signed(wire517)) ?
                      reg522[(2'h3):(1'h1)] : $signed((~^reg523))) ?
                  {((wire518 != reg533) ? (^~(8'hb7)) : reg523[(1'h0):(1'h0)]),
                      ((7'h40) >>> (reg531 ?
                          wire515 : reg528))} : reg532[(4'hc):(3'h4)])))
            begin
              reg534 <= (!reg521[(5'h13):(4'hf)]);
              reg535 <= (reg523[(3'h4):(1'h1)] ?
                  wire515 : $signed(wire518[(4'hd):(2'h2)]));
              reg536 <= {({reg523, (+(8'haf))} ?
                      $signed($unsigned($signed((8'h9c)))) : (($unsigned((8'ha0)) <= {reg535}) || ((reg521 ?
                              reg534 : (8'hbe)) ?
                          $unsigned(wire518) : reg530[(3'h6):(3'h5)])))};
              reg537 <= (($signed(($unsigned((8'hbd)) == {reg527, reg527})) ?
                      reg534 : $unsigned({reg530})) ?
                  {(((wire519 != reg534) <= reg536[(3'h5):(1'h0)]) & ((~&reg527) >= wire519)),
                      (($signed(reg534) >= $signed(reg530)) ?
                          $signed((&wire515)) : $unsigned(reg534[(4'ha):(3'h4)]))} : ((({wire518} ?
                          (-reg534) : reg534) ?
                      (^~(7'h41)) : ((reg522 + wire518) >> {reg527})) & $unsigned(reg530[(3'h5):(2'h3)])));
              reg538 <= reg520;
            end
          else
            begin
              reg534 <= ($signed($signed(wire524)) & ((^(~^(reg528 ?
                      (8'hbb) : reg529))) ?
                  $signed($signed($unsigned(wire516))) : reg522));
              reg535 <= (+($signed($signed($signed(wire518))) ?
                  ($signed(((8'hab) ?
                      wire516 : wire518)) ~^ $signed($signed(reg523))) : $unsigned($signed(reg521[(1'h0):(1'h0)]))));
              reg536 <= ((($unsigned($signed(reg520)) || reg526[(5'h11):(3'h7)]) != $signed(reg526)) ~^ reg536);
              reg537 <= (~reg536[(4'hd):(4'hd)]);
              reg538 <= (($unsigned(($signed(reg529) ?
                      $signed(wire515) : {(8'hbc),
                          reg522})) >= {reg535[(3'h7):(3'h4)],
                      ((|reg520) ^ $unsigned(reg533))}) ?
                  (($unsigned({reg526, reg523}) ^~ wire519[(1'h1):(1'h0)]) ?
                      $unsigned(reg526[(3'h7):(3'h5)]) : reg528[(3'h6):(3'h5)]) : reg520);
            end
          reg539 <= (reg520 ~^ (reg538 + $unsigned($signed((reg521 ?
              reg520 : (8'h9e))))));
          reg540 <= ($signed((-((|reg530) ^ (reg528 ?
              wire519 : reg528)))) && (^~(($signed(reg521) ?
                  reg526[(1'h0):(1'h0)] : {(8'ha4)}) ?
              reg525 : $signed(reg529))));
          if (($unsigned($unsigned({(reg520 >>> wire518), reg532})) ?
              reg532[(4'h8):(3'h5)] : $signed(((^reg525[(3'h4):(2'h2)]) << $unsigned((reg529 ?
                  reg528 : reg530))))))
            begin
              reg541 <= (((reg531 && $signed($signed(wire516))) ?
                      $unsigned($signed(wire518)) : (wire516[(3'h4):(2'h2)] >= $signed($unsigned(reg535)))) ?
                  {(((reg520 ? reg537 : wire515) ?
                          reg525[(4'hb):(3'h4)] : ((8'hb6) < reg538)) != $signed(reg537[(3'h4):(2'h3)])),
                      $signed((^~{wire518}))} : $signed((~&(reg523 ?
                      $unsigned((8'hb5)) : $signed(wire517)))));
            end
          else
            begin
              reg541 <= reg541[(1'h1):(1'h0)];
              reg542 <= wire518;
              reg543 <= {(reg531 && reg535[(3'h7):(3'h7)]),
                  reg541[(3'h6):(3'h6)]};
            end
        end
      else
        begin
          if ($signed((8'ha5)))
            begin
              reg530 <= (~&{$signed(reg539), reg530});
              reg531 <= {(reg533 ?
                      (reg521[(5'h10):(4'h9)] ?
                          ($unsigned(wire524) | reg541) : ((+reg521) ?
                              reg523 : reg529[(4'h9):(3'h7)])) : $unsigned(reg527[(2'h2):(1'h1)])),
                  reg540};
              reg532 <= wire518[(4'he):(4'ha)];
              reg533 <= (reg521[(5'h11):(5'h10)] ?
                  (^$unsigned(reg537)) : (^{$unsigned((wire516 - reg522))}));
              reg534 <= (wire519[(4'hd):(4'h9)] ?
                  {reg526[(3'h4):(2'h3)]} : (reg529 ?
                      $unsigned(reg522) : reg542));
            end
          else
            begin
              reg530 <= (8'ha5);
              reg531 <= reg540;
              reg532 <= $signed(($unsigned(reg528) ?
                  reg537 : ($signed($unsigned(wire519)) ?
                      ((reg522 ? reg522 : wire524) ?
                          (reg520 * (8'ha8)) : $unsigned(reg529)) : ($unsigned(reg542) - (wire519 ?
                          reg536 : reg523)))));
            end
          reg535 <= reg531[(1'h0):(1'h0)];
          if (reg531[(4'hb):(1'h1)])
            begin
              reg536 <= reg522;
            end
          else
            begin
              reg536 <= (8'ha1);
              reg537 <= reg531[(4'he):(4'hd)];
            end
          reg538 <= {(^(8'ha5)), ((!{(reg538 < reg525)}) || reg537)};
          reg539 <= (|($signed($unsigned($signed(reg526))) ?
              $unsigned(($unsigned(reg537) ?
                  $unsigned(wire519) : $unsigned((8'hab)))) : $unsigned($unsigned($unsigned(reg523)))));
        end
    end
  assign wire544 = $signed(reg538);
  assign wire545 = ((^~reg539) ?
                       $unsigned($unsigned({(reg527 >> reg540),
                           (reg537 ?
                               reg522 : (8'hbd))})) : (~^reg534[(4'h9):(4'h9)]));
  assign wire546 = reg542;
  assign wire547 = $unsigned($unsigned((~&$unsigned($signed(reg530)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module733
#( parameter param1914 = (((|((-(8'ha8)) ? ((8'hb4) ? (8'hb2) : (7'h44)) : {(8'ha7)})) | ((((8'hba) << (8'h9e)) + (+(8'hae))) ? {(-(8'hba))} : (~|((8'hab) < (8'hb7))))) | ((((!(8'hb7)) == ((8'ha3) >> (7'h42))) ? (~|((8'hbe) || (8'hbf))) : (~&{(8'hb5)})) >>> ((^~{(8'hb1)}) ? ({(8'had), (8'hb8)} - ((8'haa) << (8'ha9))) : ((|(8'h9c)) ? ((8'ha8) >>> (8'ha9)) : (+(8'hbf)))))) )
(y, clk, wire734, wire735, wire736, wire737, wire738);
  output wire [(32'h139):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire734;
  input wire [(5'h15):(1'h0)] wire735;
  input wire signed [(5'h15):(1'h0)] wire736;
  input wire signed [(5'h15):(1'h0)] wire737;
  input wire [(5'h12):(1'h0)] wire738;
  wire signed [(4'hf):(1'h0)] wire1913;
  wire [(4'hd):(1'h0)] wire1912;
  wire signed [(5'h10):(1'h0)] wire1911;
  wire signed [(3'h6):(1'h0)] wire1910;
  wire signed [(4'h9):(1'h0)] wire1340;
  wire signed [(5'h14):(1'h0)] wire824;
  wire [(4'he):(1'h0)] wire823;
  reg [(5'h11):(1'h0)] reg739 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire740;
  wire signed [(4'hd):(1'h0)] wire821;
  wire signed [(2'h3):(1'h0)] wire1342;
  wire [(4'h8):(1'h0)] wire1343;
  wire [(4'h8):(1'h0)] wire1344;
  wire signed [(4'hb):(1'h0)] wire1417;
  wire signed [(4'hb):(1'h0)] wire1419;
  reg signed [(5'h15):(1'h0)] reg1420 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1421 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1422 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1423 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1424 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1425 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1426 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1427 = (1'h0);
  wire [(4'ha):(1'h0)] wire1908;
  assign y = {wire1913,
                 wire1912,
                 wire1911,
                 wire1910,
                 wire1340,
                 wire824,
                 wire823,
                 reg739,
                 wire740,
                 wire821,
                 wire1342,
                 wire1343,
                 wire1344,
                 wire1417,
                 wire1419,
                 reg1420,
                 reg1421,
                 reg1422,
                 reg1423,
                 reg1424,
                 reg1425,
                 reg1426,
                 reg1427,
                 wire1908,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg739 <= ((((wire736 >>> wire735[(4'hd):(1'h1)]) ?
                  wire738[(3'h5):(2'h2)] : wire738) ?
              wire738[(2'h3):(1'h1)] : {(wire737 << (wire735 == wire734)),
                  (((8'hb1) >>> wire734) + wire738)}) ?
          $signed((~^{$signed((8'ha1))})) : (^($unsigned((~^(8'hb3))) ?
              $signed($signed(wire738)) : wire737)));
    end
  assign wire740 = $unsigned($signed($signed((^~$unsigned(wire734)))));
  module741 modinst822 (.y(wire821), .wire746(reg739), .wire745(wire737), .wire744(wire738), .wire743(wire740), .wire742(wire736), .clk(clk));
  assign wire823 = wire740;
  assign wire824 = wire740[(5'h12):(1'h0)];
  module825 modinst1341 (wire1340, clk, reg739, wire738, wire735, wire736, wire740);
  assign wire1342 = wire735[(4'hb):(2'h3)];
  assign wire1343 = $unsigned($unsigned(wire738[(1'h0):(1'h0)]));
  assign wire1344 = (8'hae);
  module1345 modinst1418 (wire1417, clk, wire740, wire1343, wire735, wire738);
  assign wire1419 = ((({wire740, (wire1344 + wire735)} <= wire738) <= ((8'hbc) ?
                        ((wire738 << wire737) ^ $unsigned(wire737)) : $signed((wire823 != wire736)))) - {wire734});
  always
    @(posedge clk) begin
      reg1420 <= wire1344[(1'h0):(1'h0)];
      if ({(~$unsigned((|(|wire824)))), wire1343[(1'h1):(1'h0)]})
        begin
          reg1421 <= reg739;
          reg1422 <= (&($signed(wire740[(5'h13):(5'h12)]) ?
              wire1417 : $unsigned($signed((wire738 - wire1344)))));
          reg1423 <= wire735[(4'hd):(3'h5)];
          reg1424 <= ((&reg739[(5'h10):(4'he)]) + wire1340[(2'h2):(1'h1)]);
        end
      else
        begin
          if ($signed(reg1420))
            begin
              reg1421 <= ((wire736 != $signed((^~(wire1419 ?
                  reg1422 : wire1340)))) && reg1424);
              reg1422 <= (&(-reg1421));
              reg1423 <= $unsigned(reg1420[(5'h14):(5'h11)]);
              reg1424 <= wire1342[(2'h3):(1'h1)];
              reg1425 <= $unsigned(wire821);
            end
          else
            begin
              reg1421 <= (!$signed(reg1421[(4'h9):(4'h8)]));
            end
          reg1426 <= $unsigned($unsigned((($signed(wire1343) ?
              (reg1422 ?
                  wire823 : reg1422) : $unsigned((8'hbd))) <<< reg1425[(4'ha):(1'h1)])));
          reg1427 <= wire1340;
        end
    end
  module1428 modinst1909 (wire1908, clk, wire738, reg1427, reg1426, wire823, wire824);
  assign wire1910 = (~reg1421[(3'h6):(3'h4)]);
  assign wire1911 = $signed(($signed({(wire735 < reg1422),
                            (reg1427 ? (8'had) : wire734)}) ?
                        (((^~wire823) & (reg1424 ?
                            wire1343 : wire735)) < (wire1910 ?
                            (+reg1421) : {wire738, wire823})) : wire735));
  assign wire1912 = (|wire1910[(1'h0):(1'h0)]);
  assign wire1913 = (7'h42);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1428
#( parameter param1907 = (~(((((8'hbc) ? (8'ha8) : (7'h41)) ? (~&(7'h42)) : {(8'hb5), (8'h9f)}) >>> ((-(7'h43)) ? ((8'hb1) ^ (8'hbb)) : {(8'ha6)})) ? {{(+(8'ha5))}, (8'ha2)} : {{((8'hbe) >= (8'hb8))}, ((&(8'hb0)) ^~ ((8'h9d) < (8'h9d)))})) )
(y, clk, wire1429, wire1430, wire1431, wire1432, wire1433);
  output wire [(32'h12c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire1429;
  input wire signed [(5'h13):(1'h0)] wire1430;
  input wire [(4'hd):(1'h0)] wire1431;
  input wire [(4'he):(1'h0)] wire1432;
  input wire [(5'h14):(1'h0)] wire1433;
  wire signed [(2'h2):(1'h0)] wire1906;
  wire signed [(5'h13):(1'h0)] wire1905;
  wire signed [(3'h4):(1'h0)] wire1903;
  wire [(4'ha):(1'h0)] wire1883;
  wire signed [(4'ha):(1'h0)] wire1882;
  wire [(3'h7):(1'h0)] wire1881;
  wire [(4'hf):(1'h0)] wire1880;
  wire [(5'h14):(1'h0)] wire1757;
  wire signed [(4'hd):(1'h0)] wire1566;
  wire signed [(5'h10):(1'h0)] wire1565;
  wire signed [(5'h15):(1'h0)] wire1564;
  wire [(5'h10):(1'h0)] wire1563;
  wire [(5'h15):(1'h0)] wire1562;
  reg [(5'h11):(1'h0)] reg1561 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1560 = (1'h0);
  reg [(5'h13):(1'h0)] reg1559 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1558 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire1434;
  wire signed [(5'h15):(1'h0)] wire1556;
  wire signed [(5'h15):(1'h0)] wire1759;
  wire [(3'h7):(1'h0)] wire1878;
  assign y = {wire1906,
                 wire1905,
                 wire1903,
                 wire1883,
                 wire1882,
                 wire1881,
                 wire1880,
                 wire1757,
                 wire1566,
                 wire1565,
                 wire1564,
                 wire1563,
                 wire1562,
                 reg1561,
                 reg1560,
                 reg1559,
                 reg1558,
                 wire1434,
                 wire1556,
                 wire1759,
                 wire1878,
                 (1'h0)};
  assign wire1434 = $unsigned(((+$signed(wire1431)) ?
                        wire1431 : wire1431[(2'h3):(1'h0)]));
  module1435 modinst1557 (.wire1438(wire1433), .clk(clk), .y(wire1556), .wire1439(wire1434), .wire1437(wire1429), .wire1440(wire1430), .wire1436(wire1431));
  always
    @(posedge clk) begin
      reg1558 <= $unsigned($unsigned({wire1430[(4'he):(4'ha)]}));
      reg1559 <= ($unsigned(($signed($signed(wire1433)) <<< wire1429[(3'h5):(1'h1)])) ?
          wire1433[(4'hd):(3'h5)] : $unsigned(wire1556));
      reg1560 <= (({(wire1434[(5'h12):(3'h7)] <<< (wire1430 ?
                  reg1559 : wire1433))} | $unsigned(wire1432[(4'hc):(2'h3)])) ?
          wire1430 : $unsigned((~^($unsigned(wire1433) ?
              (wire1434 ? (8'had) : wire1430) : $signed(wire1432)))));
      reg1561 <= (+$signed((~^$signed((!(8'hb8))))));
    end
  assign wire1562 = (|$signed(((^$signed(wire1429)) ~^ $signed({(8'hba),
                        wire1432}))));
  assign wire1563 = $unsigned($signed(wire1434));
  assign wire1564 = $unsigned((8'ha6));
  assign wire1565 = $unsigned($unsigned(wire1563));
  assign wire1566 = wire1433;
  module1567 modinst1758 (.wire1570(wire1433), .y(wire1757), .wire1572(wire1556), .clk(clk), .wire1569(wire1431), .wire1568(wire1562), .wire1571(reg1561));
  assign wire1759 = $unsigned(wire1434);
  module1760 modinst1879 (wire1878, clk, reg1559, wire1563, wire1430, reg1558, wire1564);
  assign wire1880 = $signed(reg1558[(4'hd):(1'h1)]);
  assign wire1881 = {$signed($signed($signed((^~reg1560)))),
                        $signed(wire1759[(4'hc):(3'h6)])};
  assign wire1882 = (8'ha1);
  assign wire1883 = reg1561;
  module1884 modinst1904 (wire1903, clk, wire1757, wire1556, reg1559, wire1878);
  assign wire1905 = wire1564[(3'h5):(2'h2)];
  assign wire1906 = wire1759[(5'h13):(3'h7)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1345  (y, clk, wire1349, wire1348, wire1347, wire1346);
  output wire [(32'h1bf):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire1349;
  input wire [(4'h8):(1'h0)] wire1348;
  input wire [(4'h9):(1'h0)] wire1347;
  input wire [(3'h5):(1'h0)] wire1346;
  reg [(4'hc):(1'h0)] reg1416 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1415 = (1'h0);
  reg [(5'h14):(1'h0)] reg1414 = (1'h0);
  reg [(3'h4):(1'h0)] reg1413 = (1'h0);
  wire [(5'h15):(1'h0)] wire1412;
  wire [(4'ha):(1'h0)] wire1411;
  reg signed [(3'h5):(1'h0)] reg1410 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1409 = (1'h0);
  reg [(4'hb):(1'h0)] reg1408 = (1'h0);
  reg [(2'h3):(1'h0)] reg1407 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1406 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1405 = (1'h0);
  reg [(3'h7):(1'h0)] reg1404 = (1'h0);
  reg [(2'h2):(1'h0)] reg1403 = (1'h0);
  reg [(4'hf):(1'h0)] reg1402 = (1'h0);
  reg [(4'hf):(1'h0)] reg1401 = (1'h0);
  reg [(3'h5):(1'h0)] reg1400 = (1'h0);
  reg [(2'h3):(1'h0)] reg1399 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1398 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1397 = (1'h0);
  reg [(4'ha):(1'h0)] reg1396 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1395 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1394 = (1'h0);
  reg [(4'hd):(1'h0)] reg1393 = (1'h0);
  reg [(5'h14):(1'h0)] reg1392 = (1'h0);
  reg [(4'he):(1'h0)] reg1391 = (1'h0);
  wire [(5'h13):(1'h0)] wire1390;
  wire [(5'h15):(1'h0)] wire1389;
  wire [(4'hf):(1'h0)] wire1388;
  wire signed [(5'h11):(1'h0)] wire1387;
  wire signed [(3'h6):(1'h0)] wire1386;
  wire signed [(3'h4):(1'h0)] wire1384;
  wire [(5'h11):(1'h0)] wire1353;
  wire [(4'hc):(1'h0)] wire1352;
  wire [(4'hf):(1'h0)] wire1351;
  wire signed [(5'h15):(1'h0)] wire1350;
  assign y = {reg1416,
                 reg1415,
                 reg1414,
                 reg1413,
                 wire1412,
                 wire1411,
                 reg1410,
                 reg1409,
                 reg1408,
                 reg1407,
                 reg1406,
                 reg1405,
                 reg1404,
                 reg1403,
                 reg1402,
                 reg1401,
                 reg1400,
                 reg1399,
                 reg1398,
                 reg1397,
                 reg1396,
                 reg1395,
                 reg1394,
                 reg1393,
                 reg1392,
                 reg1391,
                 wire1390,
                 wire1389,
                 wire1388,
                 wire1387,
                 wire1386,
                 wire1384,
                 wire1353,
                 wire1352,
                 wire1351,
                 wire1350,
                 (1'h0)};
  assign wire1350 = (^(wire1348[(1'h1):(1'h0)] <<< ({$signed(wire1349),
                        {wire1349, wire1346}} != {(!wire1347)})));
  assign wire1351 = ($unsigned((wire1348[(2'h2):(1'h1)] ?
                        wire1350 : wire1348)) - $signed(wire1350));
  assign wire1352 = ($unsigned($unsigned(wire1347)) ^~ wire1351);
  assign wire1353 = $unsigned((-(((!wire1346) ?
                        (wire1346 ?
                            wire1348 : (8'hbe)) : (wire1348 & wire1351)) * wire1351[(3'h5):(2'h3)])));
  module1354 modinst1385 (.wire1356(wire1352), .clk(clk), .y(wire1384), .wire1357(wire1348), .wire1358(wire1349), .wire1355(wire1353));
  assign wire1386 = $unsigned(((wire1347 ?
                        {$unsigned(wire1350)} : wire1351) <= (!(((7'h42) ?
                        wire1348 : wire1348) + (wire1351 ?
                        wire1350 : wire1348)))));
  assign wire1387 = (wire1347 >>> $unsigned((wire1353[(3'h6):(3'h5)] > $signed($unsigned(wire1348)))));
  assign wire1388 = ((wire1352[(1'h1):(1'h1)] ?
                        wire1384 : (($signed((7'h44)) ?
                            wire1384[(1'h1):(1'h0)] : $unsigned(wire1351)) & (~^$unsigned(wire1352)))) == $unsigned($unsigned(($unsigned(wire1346) ?
                        {wire1350} : $unsigned(wire1387)))));
  assign wire1389 = (wire1388 ?
                        $signed(((!{wire1348}) ?
                            (8'ha7) : ((8'hab) <= $unsigned(wire1388)))) : $unsigned(wire1349[(4'hc):(3'h4)]));
  assign wire1390 = ($signed(wire1351) >>> {(~^(^wire1387[(2'h3):(2'h3)]))});
  always
    @(posedge clk) begin
      if (((wire1353[(5'h10):(4'hc)] ?
              $signed($signed((^~wire1346))) : ((8'hb3) ?
                  (8'h9c) : $unsigned({wire1353}))) ?
          (((wire1389 ? ((8'ha5) ? wire1390 : wire1386) : $unsigned(wire1388)) ?
              (~^(~^wire1352)) : wire1390[(4'hd):(4'h8)]) || {((wire1350 ?
                  wire1346 : wire1352) ^~ $signed(wire1389)),
              {(wire1388 ? (8'hbb) : wire1389),
                  wire1389[(2'h2):(1'h0)]}}) : (!(~$signed((wire1387 ?
              wire1388 : wire1347))))))
        begin
          reg1391 <= ((((~$signed(wire1350)) ?
                      $unsigned((wire1352 ?
                          wire1347 : wire1353)) : $unsigned($signed((7'h44)))) ?
                  wire1387 : (wire1389 ?
                      (wire1388 ?
                          {(8'hba)} : ((8'h9d) ?
                              wire1348 : wire1388)) : (~^{wire1386,
                          wire1349}))) ?
              $unsigned(((wire1387[(4'hd):(3'h4)] ?
                      $unsigned(wire1386) : $signed((7'h42))) ?
                  wire1347 : ((+wire1386) ?
                      wire1387[(4'h9):(2'h3)] : wire1386[(1'h0):(1'h0)]))) : wire1347);
          reg1392 <= $unsigned(($signed({{wire1384,
                  wire1352}}) && ($unsigned(wire1346[(2'h3):(1'h1)]) <<< $unsigned(wire1389[(3'h4):(3'h4)]))));
        end
      else
        begin
          if ((((8'hbe) | ($unsigned({wire1349,
                  wire1390}) || $signed(wire1386[(2'h2):(1'h1)]))) ?
              (wire1346 >> $signed($signed($unsigned(wire1386)))) : $signed(((((8'had) ?
                      wire1347 : wire1350) ?
                  $signed(wire1350) : (wire1386 * wire1352)) == (wire1388[(4'hd):(4'hc)] ?
                  (wire1388 ? (8'haa) : wire1348) : {wire1348})))))
            begin
              reg1391 <= $unsigned((wire1348 && $unsigned($unsigned($signed(wire1347)))));
              reg1392 <= $unsigned(wire1386[(3'h6):(3'h5)]);
            end
          else
            begin
              reg1391 <= wire1387[(2'h3):(2'h3)];
            end
        end
      if ($signed((wire1384[(2'h2):(2'h2)] > (7'h42))))
        begin
          reg1393 <= reg1392;
          reg1394 <= (($unsigned(((wire1353 & wire1352) ?
                  wire1349 : (reg1391 < wire1353))) ?
              (wire1387 & $signed(wire1346[(3'h5):(2'h2)])) : wire1346[(3'h4):(2'h2)]) >> $signed($unsigned({(wire1353 ?
                  wire1389 : (8'hb0))})));
          if ((wire1346 ? {(8'ha1), wire1349} : reg1393[(3'h4):(3'h4)]))
            begin
              reg1395 <= (!((wire1387[(3'h4):(1'h1)] * $unsigned(wire1388)) >= (~|wire1389)));
              reg1396 <= {($signed(reg1394) <<< (&wire1388[(3'h6):(3'h6)]))};
              reg1397 <= (reg1393[(3'h4):(3'h4)] <<< wire1349[(2'h3):(2'h2)]);
              reg1398 <= (~&wire1347);
            end
          else
            begin
              reg1395 <= $signed($signed($signed($unsigned($signed(wire1348)))));
              reg1396 <= (~|($signed(wire1347[(3'h4):(2'h3)]) + $signed($unsigned(wire1346))));
              reg1397 <= {{($unsigned(wire1349) ?
                          (~$signed((7'h41))) : $signed({reg1397, wire1353}))}};
              reg1398 <= (wire1387 * (+($unsigned(reg1392) >> $unsigned((wire1351 ?
                  reg1396 : wire1346)))));
            end
        end
      else
        begin
          reg1393 <= wire1351[(2'h3):(2'h2)];
        end
      reg1399 <= {(&$signed(((+wire1346) ?
              $unsigned(wire1384) : wire1388[(3'h7):(1'h1)])))};
      if (wire1348)
        begin
          reg1400 <= {$unsigned((~$unsigned(reg1398[(4'hb):(3'h5)]))),
              (wire1351[(1'h0):(1'h0)] == wire1353)};
          reg1401 <= wire1348[(3'h5):(2'h3)];
          if ($unsigned($signed((^wire1390[(2'h2):(1'h1)]))))
            begin
              reg1402 <= $unsigned(((reg1395 ?
                  (!(+wire1390)) : $unsigned(wire1386)) & ((^wire1389[(4'hf):(4'h9)]) < reg1393[(2'h2):(2'h2)])));
              reg1403 <= wire1352[(2'h2):(1'h0)];
              reg1404 <= ((wire1348 ?
                  $signed((reg1393 ?
                      $signed(wire1348) : $unsigned(wire1347))) : $signed(wire1347)) <= $unsigned(reg1391));
            end
          else
            begin
              reg1402 <= ((&reg1400) == wire1347[(3'h5):(2'h2)]);
              reg1403 <= (~^(&wire1351[(3'h5):(3'h5)]));
            end
        end
      else
        begin
          reg1400 <= reg1396[(4'h8):(2'h2)];
          if ((reg1404 ?
              $unsigned($signed((wire1388 >= (reg1394 >>> reg1399)))) : ($signed($unsigned({(8'ha6)})) < $unsigned(wire1346))))
            begin
              reg1401 <= ($unsigned({($unsigned(wire1349) <<< reg1396)}) ?
                  (~|{reg1398[(5'h12):(4'hc)]}) : (8'haf));
              reg1402 <= $signed(((((reg1398 * reg1394) & $unsigned((8'hb8))) && reg1404[(2'h3):(2'h2)]) ?
                  $signed($signed((wire1352 ?
                      reg1393 : (7'h42)))) : wire1346[(1'h1):(1'h1)]));
              reg1403 <= (!(^$signed((~&{wire1389, (8'hb7)}))));
              reg1404 <= wire1388[(4'hd):(1'h0)];
              reg1405 <= (reg1400[(3'h5):(3'h4)] ?
                  reg1392 : (~^(wire1347 ?
                      $unsigned($signed(reg1404)) : reg1395[(1'h1):(1'h0)])));
            end
          else
            begin
              reg1401 <= ($signed(reg1399[(2'h2):(2'h2)]) ?
                  (reg1395 ?
                      ($signed((reg1400 ? wire1351 : wire1386)) ?
                          ((reg1395 == reg1395) != $signed(reg1405)) : ({reg1399,
                                  reg1404} ?
                              {reg1392,
                                  wire1386} : $signed(reg1393))) : wire1346) : $unsigned(((~^(wire1353 - reg1402)) == ((~^(7'h43)) ?
                      $signed(reg1394) : {wire1384, wire1348}))));
              reg1402 <= {((^~$unsigned(reg1403)) - wire1388[(3'h7):(3'h6)])};
              reg1403 <= ($signed($signed((|reg1391[(1'h0):(1'h0)]))) >= $unsigned((wire1347[(2'h2):(1'h0)] || ({reg1399,
                  wire1388} && reg1405))));
            end
          if ($signed($signed((^~(!(~^wire1351))))))
            begin
              reg1406 <= ((wire1351[(3'h7):(2'h3)] > (((reg1393 ^~ reg1393) <= reg1400) ?
                      $signed((~&wire1384)) : wire1390)) ?
                  wire1386 : (~|(~^wire1390[(3'h5):(1'h1)])));
            end
          else
            begin
              reg1406 <= $unsigned((~&(($unsigned(reg1394) ?
                  $signed((8'hbd)) : (reg1392 ?
                      wire1351 : wire1386)) + reg1397)));
              reg1407 <= {((wire1349 ?
                          (reg1400[(2'h2):(1'h1)] <<< $signed(reg1393)) : ((reg1397 != reg1400) ?
                              reg1399 : wire1390[(5'h10):(4'hb)])) ?
                      (8'hbc) : ($unsigned($unsigned(reg1393)) && $unsigned($unsigned(wire1388))))};
              reg1408 <= {{reg1397[(3'h6):(3'h6)], wire1386[(3'h5):(2'h2)]},
                  (((+wire1390) ?
                          (!reg1400[(2'h3):(1'h0)]) : ((reg1398 ?
                              wire1387 : reg1403) * $signed(reg1400))) ?
                      $signed(reg1393[(4'hd):(4'hb)]) : reg1398)};
              reg1409 <= ($signed(wire1387[(1'h0):(1'h0)]) ?
                  $signed($signed($signed((wire1384 ?
                      wire1351 : (8'hb8))))) : wire1388[(3'h4):(2'h2)]);
              reg1410 <= (+(+$signed($signed((wire1384 ?
                  (7'h40) : wire1348)))));
            end
        end
    end
  assign wire1411 = ((-wire1346[(3'h4):(3'h4)]) ?
                        $unsigned($unsigned((reg1406 ?
                            $unsigned(reg1403) : {wire1389}))) : ((($unsigned(reg1401) ?
                                (wire1390 ?
                                    reg1402 : reg1410) : reg1398[(5'h12):(1'h1)]) << (reg1394 > {reg1396})) ?
                            $unsigned($signed((+wire1346))) : $unsigned(reg1409[(4'h8):(3'h5)])));
  assign wire1412 = {(reg1409 << wire1348)};
  always
    @(posedge clk) begin
      if (($signed($signed(reg1392[(5'h12):(3'h4)])) << (~&$signed(((wire1412 & wire1351) ?
          $unsigned(wire1352) : wire1352[(4'ha):(3'h4)])))))
        begin
          reg1413 <= (($unsigned((reg1408 ^ {reg1395})) * $signed(((reg1395 * reg1402) ?
                  $unsigned(reg1404) : $unsigned(reg1400)))) ?
              (((8'ha9) >= reg1397) ?
                  {(8'hb0)} : (((wire1349 <= reg1406) || wire1352) ?
                      ((reg1393 ?
                          reg1391 : reg1406) >>> reg1398[(3'h7):(3'h4)]) : $signed(((8'hba) ?
                          (8'hb6) : reg1401)))) : $signed($unsigned(wire1411)));
          reg1414 <= wire1351;
          reg1415 <= $signed(((~(wire1352[(4'hc):(1'h0)] ?
              reg1405[(1'h1):(1'h1)] : (reg1399 ~^ reg1403))) ~^ reg1396));
          reg1416 <= $signed($unsigned((&(reg1415[(1'h1):(1'h0)] || (+reg1394)))));
        end
      else
        begin
          reg1413 <= reg1393[(4'h8):(1'h1)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module825
#( parameter param1339 = (({((8'hbc) && {(8'hb6)}), {{(8'ha4), (8'hb3)}}} | (|(~^{(8'hbf), (8'hb0)}))) >> (^~{(8'haf), {((8'hac) <<< (8'h9e))}})) )
(y, clk, wire830, wire829, wire828, wire827, wire826);
  output wire [(32'hed):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire830;
  input wire signed [(4'hb):(1'h0)] wire829;
  input wire [(5'h15):(1'h0)] wire828;
  input wire [(5'h15):(1'h0)] wire827;
  input wire [(5'h13):(1'h0)] wire826;
  wire signed [(3'h6):(1'h0)] wire1046;
  wire [(4'h8):(1'h0)] wire1048;
  wire [(5'h11):(1'h0)] wire1049;
  wire [(5'h11):(1'h0)] wire1050;
  wire [(4'h8):(1'h0)] wire1051;
  wire signed [(4'ha):(1'h0)] wire1052;
  wire [(3'h4):(1'h0)] wire1196;
  wire signed [(3'h6):(1'h0)] wire1198;
  wire signed [(5'h10):(1'h0)] wire1199;
  reg signed [(4'h9):(1'h0)] reg1200 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1201 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1202 = (1'h0);
  reg [(4'hc):(1'h0)] reg1203 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1204 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1205 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1206 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1207 = (1'h0);
  reg [(5'h11):(1'h0)] reg1208 = (1'h0);
  wire [(4'hf):(1'h0)] wire1209;
  wire signed [(4'hb):(1'h0)] wire1337;
  assign y = {wire1046,
                 wire1048,
                 wire1049,
                 wire1050,
                 wire1051,
                 wire1052,
                 wire1196,
                 wire1198,
                 wire1199,
                 reg1200,
                 reg1201,
                 reg1202,
                 reg1203,
                 reg1204,
                 reg1205,
                 reg1206,
                 reg1207,
                 reg1208,
                 wire1209,
                 wire1337,
                 (1'h0)};
  module831 modinst1047 (.wire834(wire828), .y(wire1046), .wire832(wire827), .wire835(wire830), .clk(clk), .wire836(wire829), .wire833(wire826));
  assign wire1048 = ({(((8'hac) ? (^wire1046) : wire830[(5'h10):(2'h3)]) ?
                            wire829[(4'hb):(4'hb)] : $unsigned(wire827[(5'h15):(4'hf)])),
                        ({wire1046[(1'h0):(1'h0)], (wire830 || wire829)} ?
                            ((wire827 == wire826) ?
                                wire826 : (wire827 > wire826)) : wire827)} <= (+wire827[(1'h0):(1'h0)]));
  assign wire1049 = wire829;
  assign wire1050 = $unsigned((+wire826));
  assign wire1051 = ($signed((|$signed(wire827))) || ((&(8'h9d)) ?
                        (+((8'had) ^ $signed(wire826))) : $signed(wire1050[(3'h4):(2'h3)])));
  assign wire1052 = (($signed(((|wire1048) ?
                        $signed(wire826) : (wire829 ?
                            wire830 : wire829))) > $signed(($unsigned(wire1049) ?
                        (wire830 ?
                            wire828 : wire1051) : $signed(wire1048)))) || (8'had));
  module1053 modinst1197 (.wire1056(wire830), .wire1055(wire1050), .wire1054(wire1049), .y(wire1196), .wire1057(wire828), .clk(clk));
  assign wire1198 = {($unsigned({(wire1051 || (8'hab))}) >> (7'h41))};
  assign wire1199 = wire828[(4'h9):(4'h8)];
  always
    @(posedge clk) begin
      reg1200 <= $unsigned(((($unsigned(wire828) ?
          wire1196[(1'h1):(1'h1)] : $signed((8'hbf))) + ((wire828 > wire1049) ?
          $signed((8'h9e)) : wire830[(2'h3):(1'h0)])) ~^ (wire1199[(1'h0):(1'h0)] | $unsigned(wire827))));
      if ((wire1052[(2'h2):(1'h0)] - wire1046[(1'h1):(1'h0)]))
        begin
          if ($unsigned($unsigned((^~((&wire829) < (8'ha8))))))
            begin
              reg1201 <= wire827;
            end
          else
            begin
              reg1201 <= (wire1196[(2'h2):(1'h1)] ?
                  ($signed($unsigned(reg1200[(1'h0):(1'h0)])) <= (^~$signed({wire1048}))) : $signed((wire1196[(1'h0):(1'h0)] ?
                      $signed($unsigned(wire1198)) : (wire1051[(3'h6):(1'h0)] == $unsigned(wire828)))));
            end
          if (((($unsigned(reg1200[(3'h6):(3'h4)]) > $unsigned((wire1198 & wire829))) ?
                  wire1048 : ($unsigned((8'hb9)) ?
                      ((wire830 ?
                          wire1198 : (8'hbb)) << $unsigned(wire1052)) : wire828[(4'hd):(4'hc)])) ?
              $signed((~&(wire829 && {reg1200}))) : {((~(wire828 < wire1048)) ?
                      ((~wire829) ?
                          $signed((8'hab)) : $unsigned(reg1201)) : wire1196)}))
            begin
              reg1202 <= (({wire830[(3'h4):(1'h1)]} - (^~wire828[(5'h11):(4'hf)])) ?
                  wire826 : $unsigned($unsigned($unsigned(wire827))));
              reg1203 <= $unsigned($unsigned((-($unsigned(wire1051) ?
                  (&wire1049) : $unsigned(wire1049)))));
              reg1204 <= wire1051[(3'h5):(1'h0)];
              reg1205 <= ($unsigned((~(|(-reg1201)))) || $unsigned((-($unsigned(wire829) ?
                  wire1051 : wire830))));
              reg1206 <= $signed((~^wire1048));
            end
          else
            begin
              reg1202 <= ($signed(wire1049[(4'hd):(1'h1)]) ?
                  wire1196 : (|{($unsigned(wire1199) ?
                          $unsigned(wire828) : $unsigned(reg1204))}));
            end
          reg1207 <= ($signed($unsigned(({wire1046} ?
              $signed(reg1201) : ((8'ha5) ?
                  (8'ha3) : wire826)))) == (($unsigned($signed(wire1048)) > reg1202[(3'h7):(3'h6)]) > (((wire1052 <= wire1051) < (reg1201 ^ wire1048)) ?
              ((reg1206 <= wire826) ?
                  (wire1046 ?
                      (7'h44) : wire1196) : (&wire1049)) : {wire1198[(2'h3):(2'h3)]})));
        end
      else
        begin
          if ((!($signed(((reg1206 ? wire1196 : wire829) ?
                  (reg1200 > wire829) : {(8'haf)})) ?
              $unsigned({$unsigned(wire829)}) : $unsigned((8'h9e)))))
            begin
              reg1201 <= reg1207[(2'h3):(1'h1)];
              reg1202 <= (wire827 << {((((8'haa) >> reg1207) - wire1048) - wire1199),
                  wire829[(2'h3):(1'h1)]});
            end
          else
            begin
              reg1201 <= (~^wire829);
              reg1202 <= wire1046[(3'h5):(3'h4)];
            end
          reg1203 <= (reg1203[(1'h0):(1'h0)] ?
              reg1205 : $unsigned($signed($signed((reg1200 && wire828)))));
          if ((~(-$signed(((~^wire1052) ? (!(8'ha0)) : $signed((8'hb5)))))))
            begin
              reg1204 <= (reg1203 == reg1207[(4'h9):(2'h2)]);
              reg1205 <= ((!$unsigned(wire828[(2'h2):(1'h0)])) ?
                  (&(&$signed($unsigned(reg1203)))) : (|({wire1049[(4'he):(4'h9)]} || (+wire827))));
            end
          else
            begin
              reg1204 <= wire1198[(2'h2):(2'h2)];
              reg1205 <= $signed(((-((reg1207 || wire1049) ?
                      (-wire828) : reg1200)) ?
                  (-(~|$signed(wire1051))) : reg1205));
            end
        end
      reg1208 <= reg1205[(4'h9):(4'h8)];
    end
  assign wire1209 = $signed((wire827 > wire827[(4'h8):(4'h8)]));
  module1210 modinst1338 (.wire1212(reg1206), .wire1213(wire1199), .wire1215(wire1049), .y(wire1337), .wire1211(wire1050), .wire1214(reg1203), .clk(clk));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module741
#( parameter param820 = {(+(^(8'ha7))), (~|((((8'hbf) - (8'hb6)) ? ((8'ha4) ^~ (8'hbf)) : {(7'h41)}) ? (((8'had) || (8'hb8)) ? {(8'ha5), (8'haa)} : ((8'h9e) ? (8'ha8) : (7'h43))) : (8'haf)))} )
(y, clk, wire746, wire745, wire744, wire743, wire742);
  output wire [(32'h113):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire746;
  input wire signed [(5'h15):(1'h0)] wire745;
  input wire signed [(4'h8):(1'h0)] wire744;
  input wire signed [(4'ha):(1'h0)] wire743;
  input wire signed [(5'h12):(1'h0)] wire742;
  wire signed [(4'h9):(1'h0)] wire819;
  reg [(4'h9):(1'h0)] reg818 = (1'h0);
  reg [(4'h9):(1'h0)] reg817 = (1'h0);
  reg [(4'ha):(1'h0)] reg816 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg815 = (1'h0);
  reg [(4'hb):(1'h0)] reg814 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg813 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg812 = (1'h0);
  reg [(4'hf):(1'h0)] reg811 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg810 = (1'h0);
  reg [(5'h14):(1'h0)] reg809 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg808 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg807 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg806 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire805;
  wire signed [(5'h10):(1'h0)] wire804;
  wire [(4'hb):(1'h0)] wire802;
  wire [(3'h7):(1'h0)] wire753;
  wire signed [(5'h11):(1'h0)] wire752;
  wire [(4'hd):(1'h0)] wire751;
  wire signed [(5'h12):(1'h0)] wire750;
  wire signed [(4'hd):(1'h0)] wire749;
  wire signed [(2'h2):(1'h0)] wire748;
  wire [(5'h13):(1'h0)] wire747;
  assign y = {wire819,
                 reg818,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 reg812,
                 reg811,
                 reg810,
                 reg809,
                 reg808,
                 reg807,
                 reg806,
                 wire805,
                 wire804,
                 wire802,
                 wire753,
                 wire752,
                 wire751,
                 wire750,
                 wire749,
                 wire748,
                 wire747,
                 (1'h0)};
  assign wire747 = wire746[(3'h6):(2'h3)];
  assign wire748 = $unsigned(wire745[(2'h2):(1'h1)]);
  assign wire749 = ($signed(wire744) || wire743);
  assign wire750 = $signed((!(wire744 == wire746)));
  assign wire751 = wire744[(4'h8):(2'h2)];
  assign wire752 = ($signed((wire748 ?
                       ((8'ha3) ?
                           (wire744 != wire742) : $signed(wire742)) : (wire751 ?
                           wire749[(1'h1):(1'h0)] : $unsigned(wire743)))) + {(((wire743 - wire748) && wire748[(1'h1):(1'h1)]) << (|(+wire751)))});
  assign wire753 = ($unsigned(wire746[(2'h2):(1'h1)]) ?
                       ((wire746[(1'h1):(1'h0)] && ($signed(wire752) != (~&wire751))) | $unsigned((7'h44))) : ({wire744[(3'h6):(3'h6)],
                               $signed({wire747})} ?
                           $unsigned($unsigned($unsigned(wire747))) : (wire749[(2'h2):(1'h1)] ?
                               $signed((wire748 ?
                                   wire743 : wire747)) : ((wire745 <= wire752) ?
                                   (wire749 >= wire750) : $signed(wire746)))));
  module754 modinst803 (wire802, clk, wire752, wire743, wire749, wire745);
  assign wire804 = wire742[(1'h1):(1'h1)];
  assign wire805 = {$signed((wire742[(4'h8):(4'h8)] <= ((8'hb5) >> (-wire747))))};
  always
    @(posedge clk) begin
      if ($unsigned($unsigned({$unsigned($signed(wire752)),
          (~^$signed((8'haf)))})))
        begin
          if (((&(wire805 ?
                  {(+wire745)} : (wire753[(1'h1):(1'h1)] ?
                      wire802[(3'h4):(1'h0)] : wire748))) ?
              wire742 : (wire745 ? wire747 : {(^~$unsigned(wire748))})))
            begin
              reg806 <= {wire750};
            end
          else
            begin
              reg806 <= $unsigned((!((wire751 | $signed(wire743)) ^ $signed((~&reg806)))));
              reg807 <= ((+wire748[(1'h1):(1'h1)]) ?
                  $signed(wire749[(4'h9):(2'h2)]) : wire751[(4'ha):(2'h3)]);
              reg808 <= (((&((wire751 * wire802) && (wire749 ?
                  wire744 : wire752))) ^ $signed((8'h9c))) <= $signed($signed((wire749 ?
                  (wire747 ? (8'hac) : wire748) : (8'hac)))));
              reg809 <= $signed(wire748[(1'h0):(1'h0)]);
            end
          if ($unsigned($unsigned($signed($signed(((8'hac) <<< (8'hb1)))))))
            begin
              reg810 <= $unsigned(({wire743} ~^ ({(8'hb7),
                  wire805[(3'h5):(2'h2)]} > (wire805[(2'h3):(2'h3)] ?
                  $unsigned(wire750) : (reg809 < (8'h9e))))));
              reg811 <= $unsigned((^(+($signed(wire744) ?
                  $unsigned(reg809) : reg809[(4'hf):(3'h7)]))));
              reg812 <= wire749;
              reg813 <= ($unsigned(wire747[(5'h12):(1'h0)]) && $signed(wire745));
              reg814 <= ($unsigned({$unsigned(reg812),
                      $signed(((7'h41) ? wire742 : wire744))}) ?
                  (~|wire750) : reg811);
            end
          else
            begin
              reg810 <= wire742;
            end
          reg815 <= reg806;
          reg816 <= reg806;
          reg817 <= $signed($signed($unsigned(reg813)));
        end
      else
        begin
          reg806 <= (^$unsigned($signed(reg806[(2'h2):(1'h1)])));
          reg807 <= (^$unsigned(wire802[(3'h4):(1'h1)]));
          reg808 <= $unsigned(reg809[(4'h9):(4'h9)]);
          if (wire748)
            begin
              reg809 <= ((($unsigned((reg816 >= wire749)) ~^ ((reg808 ?
                              wire744 : wire743) ?
                          (!wire804) : (wire748 != (8'ha1)))) ?
                      (($unsigned(reg814) ? (reg812 <= wire745) : wire745) ?
                          $unsigned((reg816 * (8'hbc))) : wire749[(3'h7):(3'h5)]) : $signed(((reg815 ?
                          (8'hbd) : wire753) < (|reg814)))) ?
                  (wire753 ?
                      {(8'hb0),
                          {$unsigned(wire744)}} : wire749) : ((((wire746 >>> reg806) ?
                          $signed(wire744) : $signed(reg816)) ?
                      $signed(((8'ha0) | reg809)) : reg814[(1'h0):(1'h0)]) < $signed(((reg814 ?
                          reg812 : reg813) ?
                      $unsigned(reg807) : (reg816 & reg806)))));
              reg810 <= $signed({wire748, reg817});
              reg811 <= wire750;
              reg812 <= (~|($signed($unsigned(reg806[(1'h1):(1'h0)])) | (((^~wire805) <= (8'hbd)) + wire748[(1'h1):(1'h1)])));
              reg813 <= (|reg807[(1'h0):(1'h0)]);
            end
          else
            begin
              reg809 <= (^~({$unsigned((~&wire744)),
                  (-reg811)} << ($signed($unsigned((8'ha4))) + reg808[(3'h7):(3'h4)])));
              reg810 <= ((~|(~&$unsigned((wire750 ? wire752 : reg807)))) ?
                  $unsigned((|$signed((reg813 ?
                      wire748 : wire749)))) : $unsigned($unsigned(wire745[(5'h11):(4'hb)])));
              reg811 <= $signed((^~wire746[(2'h3):(2'h3)]));
              reg812 <= ($signed($signed(wire743)) & reg808);
            end
          if ($signed($unsigned((~&$unsigned({wire747})))))
            begin
              reg814 <= (~|(|wire749));
              reg815 <= reg816[(2'h2):(1'h1)];
              reg816 <= wire805;
              reg817 <= ($unsigned(($unsigned(wire804) || reg806)) ?
                  wire749[(3'h4):(2'h3)] : (~^$unsigned(((wire744 ?
                          (8'haf) : wire747) ?
                      {wire742} : $signed(wire804)))));
              reg818 <= reg813[(4'ha):(1'h0)];
            end
          else
            begin
              reg814 <= {$unsigned({($signed(wire751) + reg814),
                      ($signed(wire742) ?
                          $signed(reg817) : (reg812 && wire804))}),
                  $unsigned((wire805 ?
                      wire743[(3'h6):(3'h6)] : (~$unsigned(wire742))))};
              reg815 <= {reg817};
              reg816 <= reg808;
              reg817 <= (8'hb6);
            end
        end
    end
  assign wire819 = (((wire804 >> (!(-(8'hae)))) ?
                           ((^wire747[(5'h10):(5'h10)]) ?
                               {(wire743 <= wire750)} : $unsigned(reg813)) : reg808) ?
                       $signed($unsigned((~^reg810[(4'h9):(2'h3)]))) : $signed((|(-$signed(reg812)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module754  (y, clk, wire758, wire757, wire756, wire755);
  output wire [(32'hb6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire758;
  input wire signed [(4'h8):(1'h0)] wire757;
  input wire [(4'hd):(1'h0)] wire756;
  input wire signed [(4'he):(1'h0)] wire755;
  wire signed [(4'h8):(1'h0)] wire801;
  wire signed [(5'h12):(1'h0)] wire800;
  wire [(5'h14):(1'h0)] wire799;
  reg signed [(5'h12):(1'h0)] reg798 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg797 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg796 = (1'h0);
  reg [(5'h13):(1'h0)] reg795 = (1'h0);
  reg [(3'h6):(1'h0)] reg794 = (1'h0);
  reg [(4'hf):(1'h0)] reg793 = (1'h0);
  reg [(5'h11):(1'h0)] reg792 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire791;
  wire signed [(3'h7):(1'h0)] wire790;
  wire signed [(2'h3):(1'h0)] wire788;
  assign y = {wire801,
                 wire800,
                 wire799,
                 reg798,
                 reg797,
                 reg796,
                 reg795,
                 reg794,
                 reg793,
                 reg792,
                 wire791,
                 wire790,
                 wire788,
                 (1'h0)};
  module759 modinst789 (.y(wire788), .wire763(wire756), .wire761(wire757), .wire760((8'hbc)), .clk(clk), .wire764(wire758), .wire762(wire755));
  assign wire790 = (wire757[(2'h2):(1'h0)] ?
                       $unsigned($signed((wire755 ?
                           wire756[(2'h3):(1'h1)] : wire755))) : $signed($unsigned(wire756)));
  assign wire791 = $unsigned($unsigned(($unsigned(((8'hb3) ?
                       wire758 : wire790)) || {wire790})));
  always
    @(posedge clk) begin
      reg792 <= wire790;
      if (((8'hae) ? $unsigned(wire790) : $unsigned(wire790)))
        begin
          if ((~(~(&reg792[(4'hb):(3'h4)]))))
            begin
              reg793 <= (wire755 << ($unsigned((wire757 <= (wire756 ?
                      wire758 : reg792))) ?
                  ($unsigned(wire756) ?
                      (-wire791[(1'h0):(1'h0)]) : $signed(wire791)) : {(wire756[(3'h6):(2'h2)] ?
                          $unsigned(wire790) : $signed((8'haf)))}));
              reg794 <= ($unsigned($unsigned((wire788[(1'h0):(1'h0)] | (-(8'h9d))))) | wire790);
            end
          else
            begin
              reg793 <= reg793;
              reg794 <= $unsigned(wire755);
              reg795 <= wire755[(3'h7):(2'h2)];
              reg796 <= ((wire791 << $unsigned($signed((reg794 ?
                  (8'hb7) : wire756)))) & reg792);
            end
        end
      else
        begin
          if (wire788[(1'h1):(1'h0)])
            begin
              reg793 <= (~|$unsigned(reg792[(3'h5):(1'h0)]));
              reg794 <= (reg794 * {(+$signed((wire755 ? reg796 : wire791)))});
            end
          else
            begin
              reg793 <= $signed((wire788[(2'h2):(1'h0)] ?
                  $unsigned($unsigned(reg796[(4'he):(4'h8)])) : {$unsigned((wire788 == reg796)),
                      $unsigned((reg796 ? wire755 : reg792))}));
              reg794 <= reg794[(1'h1):(1'h1)];
              reg795 <= reg792;
              reg796 <= $unsigned($signed(($signed(wire755) ?
                  {(wire756 ? wire791 : wire788),
                      reg793[(3'h6):(1'h0)]} : {wire756, reg795})));
              reg797 <= ((wire756[(3'h7):(2'h3)] ?
                  (~|(8'hbb)) : {(8'ha7)}) != $unsigned(wire755[(2'h3):(1'h0)]));
            end
        end
      reg798 <= (wire790[(2'h2):(2'h2)] ?
          reg796 : ((wire755 <<< {{(8'hb4)}}) != (reg794[(3'h4):(2'h3)] != wire756[(1'h1):(1'h1)])));
    end
  assign wire799 = $signed(wire756);
  assign wire800 = (wire788 ?
                       {$signed(wire756[(2'h2):(1'h0)])} : (~($unsigned(((8'hbd) ?
                               wire790 : wire791)) ?
                           ($unsigned((8'hb3)) ?
                               wire790 : (wire755 >>> (8'haa))) : ((&reg792) ?
                               {(8'hbe), (8'hba)} : {wire755}))));
  assign wire801 = (^~$signed((|$signed($unsigned(reg797)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module759
#( parameter param786 = (((((^(8'hbe)) < {(8'hb1)}) ~^ (&(8'h9e))) || ((!((8'ha4) * (8'hbf))) ? (((8'ha5) ? (7'h41) : (8'hbb)) >>> (^~(8'hbb))) : (((8'hb6) <<< (7'h42)) | ((8'ha0) ~^ (8'hb1))))) ? (({(&(8'hb9)), (|(8'hab))} != (~^{(7'h42), (8'had)})) ? {(7'h40)} : (&(((8'hb3) < (8'hb3)) ? ((8'had) < (8'ha7)) : (~|(8'ha9))))) : (|(((~|(8'hb9)) > ((8'hbd) ? (8'h9f) : (8'hba))) ? (((8'ha0) ? (8'hba) : (8'haa)) ? {(8'hab)} : ((8'ha7) > (8'hb0))) : (~((7'h44) ? (8'hb1) : (8'hb6))))))
, parameter param787 = (&((8'hb3) << (((param786 * param786) ? (|param786) : (param786 ? param786 : param786)) ~^ {(param786 ^ param786), (|param786)}))) )
(y, clk, wire764, wire763, wire762, wire761, wire760);
  output wire [(32'hf1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire764;
  input wire [(4'hb):(1'h0)] wire763;
  input wire signed [(4'he):(1'h0)] wire762;
  input wire signed [(4'h8):(1'h0)] wire761;
  input wire signed [(2'h2):(1'h0)] wire760;
  wire [(4'h9):(1'h0)] wire785;
  wire signed [(4'hd):(1'h0)] wire784;
  wire signed [(2'h2):(1'h0)] wire783;
  reg [(3'h7):(1'h0)] reg782 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg781 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg780 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire779;
  wire [(3'h6):(1'h0)] wire778;
  wire [(5'h13):(1'h0)] wire777;
  wire signed [(5'h14):(1'h0)] wire776;
  wire signed [(5'h12):(1'h0)] wire775;
  reg signed [(3'h6):(1'h0)] reg774 = (1'h0);
  reg [(3'h7):(1'h0)] reg773 = (1'h0);
  reg [(4'ha):(1'h0)] reg772 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg771 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg770 = (1'h0);
  reg [(4'hd):(1'h0)] reg769 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg768 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg767 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg766 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire765;
  assign y = {wire785,
                 wire784,
                 wire783,
                 reg782,
                 reg781,
                 reg780,
                 wire779,
                 wire778,
                 wire777,
                 wire776,
                 wire775,
                 reg774,
                 reg773,
                 reg772,
                 reg771,
                 reg770,
                 reg769,
                 reg768,
                 reg767,
                 reg766,
                 wire765,
                 (1'h0)};
  assign wire765 = (((-$signed($unsigned(wire763))) < {(8'h9f),
                       $unsigned($unsigned((8'hbd)))}) << (+(~^(((8'ha9) ?
                       wire763 : wire763) << (wire761 ? wire764 : wire760)))));
  always
    @(posedge clk) begin
      if ((wire762 != (($unsigned($unsigned(wire762)) ?
          (~^$signed(wire761)) : $unsigned((~|(8'haf)))) - (-({wire761,
          wire761} < wire763)))))
        begin
          if (wire762)
            begin
              reg766 <= $signed({($signed((wire762 ^~ wire762)) ?
                      (~^{(8'hb6)}) : wire763[(4'hb):(3'h5)])});
              reg767 <= $unsigned($signed(wire761));
              reg768 <= $signed((~^wire763[(4'hb):(1'h0)]));
              reg769 <= (($unsigned(reg766[(3'h7):(3'h4)]) ?
                      $unsigned(((wire765 ? (8'had) : wire764) ?
                          (^~wire764) : (wire762 || reg768))) : reg768) ?
                  ((-$unsigned((wire765 ? wire763 : wire760))) ?
                      ((wire765 ? reg767[(5'h14):(5'h14)] : (~&reg767)) ?
                          {(wire764 ? reg766 : wire762)} : $signed(((8'ha1) ?
                              wire763 : reg766))) : $signed(reg768)) : $unsigned((({(8'hab),
                      wire762} < $unsigned(wire762)) == ({wire762,
                      (8'hae)} && (-wire764)))));
            end
          else
            begin
              reg766 <= (reg766[(3'h6):(2'h3)] < reg769);
              reg767 <= {$unsigned((($unsigned(wire761) ^~ $unsigned(reg766)) | {reg769,
                      (~|(8'hbc))})),
                  $unsigned({$unsigned($unsigned(wire765))})};
            end
          reg770 <= wire762[(2'h2):(1'h1)];
        end
      else
        begin
          reg766 <= (($unsigned((~^$unsigned(wire763))) ?
                  ((wire764[(5'h10):(4'h9)] ?
                      {(8'ha4)} : wire764) <<< (~^reg767[(4'hf):(4'h8)])) : reg769) ?
              ($unsigned(wire764) && $signed(wire761[(3'h7):(1'h1)])) : ($unsigned((wire761 ?
                      (reg768 ? wire763 : wire762) : ((8'had) ?
                          wire761 : (8'hb1)))) ?
                  $signed($signed((-(8'hab)))) : wire763));
          reg767 <= reg767[(1'h0):(1'h0)];
          reg768 <= wire765;
        end
      reg771 <= (wire763[(2'h2):(1'h0)] ? wire763[(3'h6):(3'h4)] : wire763);
      reg772 <= reg770;
      reg773 <= reg769;
      reg774 <= reg767;
    end
  assign wire775 = $unsigned({(reg773 <<< wire765)});
  assign wire776 = reg767[(4'ha):(2'h2)];
  assign wire777 = $unsigned((wire764[(3'h7):(2'h3)] ?
                       (^wire776) : $signed($signed($unsigned(reg768)))));
  assign wire778 = $unsigned((8'hbc));
  assign wire779 = (^$signed($unsigned((reg771 || ((8'had) >>> reg773)))));
  always
    @(posedge clk) begin
      reg780 <= $signed({(~|((-reg766) > {wire763, wire765}))});
      reg781 <= reg773[(1'h1):(1'h0)];
      reg782 <= (~|$unsigned(((!(^~wire765)) ?
          $signed(reg774) : (((8'hb2) && reg772) ?
              ((8'hbc) ~^ wire777) : (^~wire765)))));
    end
  assign wire783 = reg769[(3'h4):(2'h3)];
  assign wire784 = reg769;
  assign wire785 = reg782[(3'h6):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1210  (y, clk, wire1215, wire1214, wire1213, wire1212, wire1211);
  output wire [(32'h116):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire1215;
  input wire signed [(4'hc):(1'h0)] wire1214;
  input wire [(5'h10):(1'h0)] wire1213;
  input wire signed [(4'hf):(1'h0)] wire1212;
  input wire signed [(4'ha):(1'h0)] wire1211;
  wire [(3'h6):(1'h0)] wire1336;
  reg [(2'h3):(1'h0)] reg1335 = (1'h0);
  reg [(5'h15):(1'h0)] reg1334 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1333 = (1'h0);
  wire [(3'h5):(1'h0)] wire1332;
  wire [(5'h13):(1'h0)] wire1331;
  wire signed [(3'h5):(1'h0)] wire1330;
  wire signed [(5'h12):(1'h0)] wire1329;
  wire [(5'h13):(1'h0)] wire1328;
  wire signed [(4'h9):(1'h0)] wire1327;
  wire signed [(2'h2):(1'h0)] wire1326;
  wire signed [(5'h10):(1'h0)] wire1293;
  wire [(5'h11):(1'h0)] wire1221;
  wire signed [(3'h4):(1'h0)] wire1220;
  wire [(4'ha):(1'h0)] wire1219;
  wire [(2'h2):(1'h0)] wire1218;
  wire signed [(5'h13):(1'h0)] wire1217;
  wire [(5'h15):(1'h0)] wire1216;
  wire signed [(5'h11):(1'h0)] wire1295;
  wire [(4'hc):(1'h0)] wire1296;
  wire [(4'hd):(1'h0)] wire1297;
  wire signed [(5'h15):(1'h0)] wire1298;
  wire [(4'h8):(1'h0)] wire1324;
  assign y = {wire1336,
                 reg1335,
                 reg1334,
                 reg1333,
                 wire1332,
                 wire1331,
                 wire1330,
                 wire1329,
                 wire1328,
                 wire1327,
                 wire1326,
                 wire1293,
                 wire1221,
                 wire1220,
                 wire1219,
                 wire1218,
                 wire1217,
                 wire1216,
                 wire1295,
                 wire1296,
                 wire1297,
                 wire1298,
                 wire1324,
                 (1'h0)};
  assign wire1216 = $unsigned($unsigned($signed($unsigned(wire1211[(1'h1):(1'h1)]))));
  assign wire1217 = {$signed($unsigned($unsigned($unsigned((8'ha2)))))};
  assign wire1218 = $signed(wire1213);
  assign wire1219 = {(^~wire1212), $unsigned((~^(8'ha1)))};
  assign wire1220 = (-wire1216);
  assign wire1221 = wire1220[(1'h1):(1'h0)];
  module1222 modinst1294 (.clk(clk), .wire1225(wire1211), .wire1224(wire1219), .wire1227(wire1216), .y(wire1293), .wire1223(wire1217), .wire1226(wire1215));
  assign wire1295 = ((|({(~|wire1221)} >>> ((wire1219 ? wire1219 : (8'ha8)) ?
                        (~&wire1213) : (wire1218 + wire1214)))) >>> (((~|(wire1219 ?
                            (8'hb4) : wire1211)) ?
                        $signed(wire1214[(4'hb):(3'h7)]) : wire1219[(1'h0):(1'h0)]) <<< (^~((wire1220 ?
                            wire1216 : wire1219) ?
                        wire1214[(4'h8):(1'h0)] : (wire1221 * wire1216)))));
  assign wire1296 = (~^$signed((~|$unsigned($signed(wire1221)))));
  assign wire1297 = $unsigned(wire1217);
  assign wire1298 = $unsigned(wire1217);
  module1299 modinst1325 (.wire1303(wire1298), .y(wire1324), .wire1304(wire1221), .wire1300(wire1212), .wire1302(wire1216), .wire1301(wire1217), .clk(clk));
  assign wire1326 = $signed((8'hb2));
  assign wire1327 = wire1216[(4'ha):(3'h6)];
  assign wire1328 = wire1211;
  assign wire1329 = wire1293[(5'h10):(2'h2)];
  assign wire1330 = ((($signed({wire1329}) + $signed($signed(wire1328))) ^ {($unsigned(wire1295) - wire1213[(3'h7):(3'h5)]),
                            {(~^wire1221)}}) ?
                        ($unsigned(wire1211[(4'ha):(1'h0)]) && (wire1215[(3'h4):(1'h0)] ?
                            (^~(wire1220 >>> wire1296)) : (~^(8'ha5)))) : (wire1326 ?
                            ((&(wire1219 == wire1296)) ?
                                (wire1328 ?
                                    (wire1297 >>> wire1326) : {wire1324,
                                        wire1324}) : (8'had)) : $unsigned(wire1328)));
  assign wire1331 = ((&$signed($unsigned($unsigned(wire1211)))) <<< (wire1329[(4'hd):(3'h5)] ?
                        {wire1216,
                            $unsigned((8'hac))} : (&{$unsigned(wire1297)})));
  assign wire1332 = ((-wire1328) ?
                        {wire1293,
                            $unsigned(wire1329)} : wire1326[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg1333 <= (8'hac);
      reg1334 <= wire1220[(1'h0):(1'h0)];
      reg1335 <= (wire1324 ? (~|wire1293[(4'hb):(3'h6)]) : wire1221);
    end
  assign wire1336 = (-wire1329[(5'h12):(4'hf)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1053
#(parameter param1195 = (8'had))
(y, clk, wire1054, wire1055, wire1056, wire1057);
  output wire [(32'h22d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire1054;
  input wire [(5'h11):(1'h0)] wire1055;
  input wire signed [(4'h8):(1'h0)] wire1056;
  input wire signed [(4'hb):(1'h0)] wire1057;
  wire [(5'h15):(1'h0)] wire1194;
  wire signed [(4'he):(1'h0)] wire1193;
  wire signed [(4'hf):(1'h0)] wire1192;
  wire [(5'h15):(1'h0)] wire1191;
  wire signed [(5'h14):(1'h0)] wire1190;
  wire [(4'hb):(1'h0)] wire1189;
  wire signed [(4'he):(1'h0)] wire1188;
  wire [(3'h7):(1'h0)] wire1187;
  wire [(4'ha):(1'h0)] wire1058;
  wire signed [(3'h7):(1'h0)] wire1059;
  wire signed [(5'h12):(1'h0)] wire1060;
  wire signed [(4'h9):(1'h0)] wire1061;
  reg [(5'h13):(1'h0)] reg1062 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1063 = (1'h0);
  reg [(4'hf):(1'h0)] reg1064 = (1'h0);
  reg [(4'h8):(1'h0)] reg1065 = (1'h0);
  reg [(3'h7):(1'h0)] reg1066 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1067 = (1'h0);
  reg [(5'h15):(1'h0)] reg1068 = (1'h0);
  reg [(3'h6):(1'h0)] reg1069 = (1'h0);
  reg [(4'hf):(1'h0)] reg1070 = (1'h0);
  reg [(3'h4):(1'h0)] reg1071 = (1'h0);
  wire [(4'hf):(1'h0)] wire1072;
  wire [(2'h3):(1'h0)] wire1073;
  reg signed [(3'h6):(1'h0)] reg1074 = (1'h0);
  reg [(4'hb):(1'h0)] reg1075 = (1'h0);
  reg [(5'h14):(1'h0)] reg1076 = (1'h0);
  reg [(4'he):(1'h0)] reg1077 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1078 = (1'h0);
  reg [(5'h11):(1'h0)] reg1079 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1080 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1081 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1082 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1083 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1084 = (1'h0);
  reg [(5'h11):(1'h0)] reg1085 = (1'h0);
  reg [(5'h13):(1'h0)] reg1086 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1087 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1088 = (1'h0);
  reg [(3'h5):(1'h0)] reg1089 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire1090;
  wire signed [(5'h10):(1'h0)] wire1185;
  assign y = {wire1194,
                 wire1193,
                 wire1192,
                 wire1191,
                 wire1190,
                 wire1189,
                 wire1188,
                 wire1187,
                 wire1058,
                 wire1059,
                 wire1060,
                 wire1061,
                 reg1062,
                 reg1063,
                 reg1064,
                 reg1065,
                 reg1066,
                 reg1067,
                 reg1068,
                 reg1069,
                 reg1070,
                 reg1071,
                 wire1072,
                 wire1073,
                 reg1074,
                 reg1075,
                 reg1076,
                 reg1077,
                 reg1078,
                 reg1079,
                 reg1080,
                 reg1081,
                 reg1082,
                 reg1083,
                 reg1084,
                 reg1085,
                 reg1086,
                 reg1087,
                 reg1088,
                 reg1089,
                 wire1090,
                 wire1185,
                 (1'h0)};
  assign wire1058 = ({$unsigned(wire1055)} + (($signed((wire1054 ?
                        wire1055 : (8'hb6))) != ({wire1055, (8'hab)} ?
                        $unsigned((8'ha4)) : ((8'haf) ?
                            (8'ha6) : wire1057))) > {wire1056, wire1056}));
  assign wire1059 = $unsigned(($unsigned((((8'ha6) <<< wire1057) > wire1056)) ?
                        wire1057 : $unsigned((~|wire1054))));
  assign wire1060 = ((+$signed(wire1058[(4'ha):(1'h1)])) && wire1059[(2'h3):(1'h0)]);
  assign wire1061 = ((|(8'h9e)) + $signed(wire1054));
  always
    @(posedge clk) begin
      reg1062 <= ({wire1055} && wire1060);
      reg1063 <= $unsigned(wire1057);
      reg1064 <= (((^~((wire1054 ? wire1055 : wire1054) && {reg1063})) ?
          wire1059[(3'h7):(1'h1)] : $unsigned((^$unsigned((8'hae))))) || {$unsigned(wire1056[(2'h2):(1'h1)])});
      if (wire1057[(2'h2):(1'h0)])
        begin
          reg1065 <= (~&(^~(8'h9d)));
          reg1066 <= ($unsigned(($signed((~wire1056)) ?
                  (|(7'h42)) : $signed((reg1062 ? wire1060 : wire1058)))) ?
              reg1063[(4'h9):(2'h2)] : wire1055[(4'h8):(2'h2)]);
          reg1067 <= (~^(~|$unsigned((wire1056[(3'h6):(1'h0)] >> wire1055[(5'h10):(2'h3)]))));
        end
      else
        begin
          if (((((+reg1066) <<< wire1061) >>> wire1061[(3'h7):(1'h1)]) ?
              $unsigned(reg1066) : $signed((((~^wire1060) ?
                      ((8'hb0) ? wire1060 : wire1054) : ((8'hb8) <<< (7'h44))) ?
                  $unsigned($signed((8'hb4))) : wire1058))))
            begin
              reg1065 <= (8'haa);
              reg1066 <= reg1063[(1'h1):(1'h1)];
              reg1067 <= $signed(wire1058);
              reg1068 <= $signed($signed(reg1067));
            end
          else
            begin
              reg1065 <= ($unsigned(reg1063) - wire1060);
              reg1066 <= ($signed((8'hbe)) ?
                  wire1055 : (|reg1062[(2'h2):(1'h1)]));
              reg1067 <= (wire1060 ?
                  reg1064[(4'ha):(4'h8)] : (wire1061[(2'h2):(1'h1)] < (((8'hab) - reg1068) ?
                      {(~&wire1058)} : $signed(wire1055))));
              reg1068 <= (({(wire1059 ?
                              (reg1066 < reg1065) : reg1068[(2'h2):(1'h1)]),
                          $signed(((8'hb7) ? wire1054 : wire1061))} ?
                      wire1059[(3'h7):(3'h4)] : wire1058) ?
                  $signed($unsigned((8'ha7))) : (+reg1066[(3'h7):(2'h3)]));
            end
          reg1069 <= $signed($unsigned($unsigned($signed($signed(wire1054)))));
          reg1070 <= {wire1056, reg1069[(3'h4):(2'h2)]};
          reg1071 <= {((+wire1058) >> $signed(($unsigned(reg1065) > (reg1065 ?
                  reg1065 : (8'had))))),
              $signed($signed($unsigned((~|reg1070))))};
        end
    end
  assign wire1072 = wire1060[(4'hc):(3'h4)];
  assign wire1073 = {($signed(wire1058) >>> (&{wire1056}))};
  always
    @(posedge clk) begin
      reg1074 <= $unsigned(reg1066);
      reg1075 <= reg1068[(4'hb):(2'h3)];
      if (wire1060[(2'h2):(1'h0)])
        begin
          if ((wire1061 ?
              {(!((8'hbb) ? reg1075 : (reg1070 ? wire1073 : wire1057))),
                  reg1074[(3'h4):(2'h2)]} : (($signed($signed(wire1058)) <= ((reg1063 && (8'hb8)) + ((8'ha5) ~^ wire1058))) ?
                  (8'hb8) : reg1066)))
            begin
              reg1076 <= ((((&(reg1067 == reg1067)) > (|(8'hb8))) ?
                  (((wire1072 <<< wire1058) > $signed(wire1072)) ?
                      (~|reg1068) : $signed((reg1065 ^ reg1075))) : ((reg1065 + $unsigned((8'hb7))) >= $unsigned({reg1071,
                      wire1073}))) & (({reg1067[(1'h0):(1'h0)]} ?
                  {(reg1069 ? reg1071 : wire1056),
                      reg1068[(4'h8):(3'h5)]} : ({wire1054} ?
                      $unsigned(wire1055) : $unsigned(reg1064))) | (8'hb8)));
              reg1077 <= ($signed(((~wire1058) >= reg1063)) <= ({{$unsigned((7'h42))},
                      reg1066[(3'h7):(1'h1)]} ?
                  reg1064 : (reg1063 >> ($signed(wire1073) >> (8'ha8)))));
              reg1078 <= reg1066[(2'h3):(1'h1)];
              reg1079 <= $signed(reg1069[(2'h2):(1'h1)]);
              reg1080 <= $unsigned(((reg1078 ?
                  ((reg1065 && reg1075) ?
                      $signed(wire1056) : reg1063) : $unsigned(((7'h43) ?
                      (8'hab) : wire1057))) & {reg1078,
                  $unsigned($signed(reg1067))}));
            end
          else
            begin
              reg1076 <= (+reg1068);
              reg1077 <= $unsigned($signed(reg1062[(4'h8):(3'h6)]));
              reg1078 <= reg1062[(4'hd):(4'hc)];
            end
          if (reg1069)
            begin
              reg1081 <= (~|(-(|(!$signed(reg1077)))));
              reg1082 <= ((^reg1066) ?
                  $signed((-wire1060[(3'h5):(3'h4)])) : reg1069);
              reg1083 <= (&(~reg1077[(4'hb):(3'h4)]));
              reg1084 <= $unsigned($signed(((reg1080[(1'h1):(1'h0)] <= (wire1054 ?
                      reg1077 : reg1064)) ?
                  reg1076 : (reg1081 ?
                      reg1079[(2'h3):(1'h1)] : (wire1073 ?
                          (8'hab) : wire1058)))));
              reg1085 <= reg1062;
            end
          else
            begin
              reg1081 <= (7'h43);
              reg1082 <= $unsigned(reg1076[(1'h1):(1'h1)]);
              reg1083 <= (~&wire1072);
              reg1084 <= (~^$signed((($signed(reg1075) - $signed(wire1054)) ?
                  wire1056[(3'h7):(3'h5)] : ({(8'hb1), reg1069} < (8'ha7)))));
              reg1085 <= $unsigned((-$signed(wire1058)));
            end
          reg1086 <= $signed(reg1069);
          reg1087 <= $signed(reg1063);
          reg1088 <= wire1054[(4'hd):(1'h0)];
        end
      else
        begin
          if (wire1056)
            begin
              reg1076 <= reg1062;
              reg1077 <= ((((reg1076[(5'h10):(4'hd)] * (reg1088 ?
                  reg1074 : wire1057)) <= ((wire1056 ? (8'hba) : (8'hb6)) ?
                  (reg1079 ? wire1058 : wire1058) : (reg1087 ?
                      reg1084 : reg1075))) << $signed((reg1081[(5'h11):(3'h5)] & ((8'hbd) ?
                  reg1066 : reg1086)))) & ($unsigned((reg1069 ?
                      (-reg1083) : (wire1061 != reg1082))) ?
                  (+$unsigned({(8'hb9)})) : reg1071[(2'h2):(2'h2)]));
              reg1078 <= $unsigned((($unsigned($signed(wire1060)) ?
                  (8'ha8) : (~|reg1085)) > $unsigned((&reg1079[(1'h0):(1'h0)]))));
              reg1079 <= $unsigned((~&(wire1055[(3'h6):(3'h5)] ?
                  $signed(reg1065) : (-(!(8'ha5))))));
              reg1080 <= ((&$signed(wire1058)) ?
                  $unsigned((^~$signed($signed(reg1087)))) : reg1069[(2'h3):(2'h3)]);
            end
          else
            begin
              reg1076 <= reg1064;
              reg1077 <= reg1079;
              reg1078 <= ((~((8'haa) << (^{wire1057,
                  wire1073}))) <= {wire1060[(4'hf):(2'h3)], reg1070});
              reg1079 <= (((+(~&reg1066[(3'h4):(3'h4)])) ?
                  (+(^~(~^reg1071))) : wire1055[(2'h2):(1'h0)]) + $signed(wire1073));
            end
          reg1081 <= (^~reg1070[(3'h5):(3'h5)]);
          if (reg1086)
            begin
              reg1082 <= (8'hb5);
              reg1083 <= $unsigned(reg1065[(1'h0):(1'h0)]);
              reg1084 <= ({(~&(~reg1069))} ?
                  ((reg1068[(5'h10):(3'h4)] < $unsigned((reg1077 > reg1082))) <= $signed(reg1083[(2'h3):(2'h2)])) : (reg1070 + reg1069[(1'h0):(1'h0)]));
            end
          else
            begin
              reg1082 <= $unsigned({reg1084,
                  ({reg1077} <<< $signed($unsigned(wire1061)))});
              reg1083 <= (^reg1088);
            end
          if ($unsigned($unsigned(wire1059)))
            begin
              reg1085 <= (reg1074[(1'h1):(1'h1)] ?
                  $unsigned((-({reg1085} & (reg1067 ^~ reg1080)))) : ((~&(wire1056 ?
                          reg1081[(5'h13):(2'h3)] : (reg1079 | reg1064))) ?
                      (+{((8'hbc) != (8'hbf))}) : {(wire1060[(4'hc):(3'h5)] == reg1062[(5'h13):(3'h6)]),
                          $signed($unsigned(reg1076))}));
              reg1086 <= $unsigned($unsigned((((reg1067 ? (8'ha8) : (8'hbe)) ?
                      (|reg1087) : $signed(wire1058)) ?
                  (~&{wire1057}) : $unsigned(wire1054[(2'h3):(1'h1)]))));
              reg1087 <= ($signed(reg1087) ?
                  (~&{reg1068[(3'h5):(1'h0)]}) : $signed({($signed(reg1063) || ((7'h42) ?
                          reg1088 : wire1056))}));
              reg1088 <= (((($signed(reg1079) ?
                  (~&reg1076) : (~wire1055)) && reg1083[(2'h2):(1'h0)]) == {wire1061,
                  (reg1087[(3'h7):(3'h5)] ~^ reg1070[(4'h9):(2'h2)])}) ^~ $signed((~|$unsigned(wire1060))));
            end
          else
            begin
              reg1085 <= reg1079[(3'h5):(1'h1)];
              reg1086 <= (reg1070[(3'h4):(3'h4)] * (|reg1078[(4'hc):(1'h0)]));
              reg1087 <= ({{$signed(((8'h9e) < reg1066)),
                      wire1059[(3'h5):(1'h1)]}} || $unsigned($unsigned((~^(+reg1069)))));
              reg1088 <= ($signed((~(reg1083 ?
                  $signed(reg1083) : (~&reg1078)))) << reg1071);
            end
          reg1089 <= $unsigned((~^$signed($signed((wire1061 ?
              reg1066 : (7'h43))))));
        end
    end
  assign wire1090 = $signed($signed($signed(((~&reg1087) ?
                        (reg1084 && wire1055) : wire1061))));
  module1091 modinst1186 (wire1185, clk, reg1062, reg1077, reg1088, reg1068, reg1067);
  assign wire1187 = {reg1089[(3'h5):(1'h1)]};
  assign wire1188 = wire1056;
  assign wire1189 = (wire1185[(2'h3):(1'h0)] ?
                        (8'hb1) : reg1086[(4'he):(1'h1)]);
  assign wire1190 = ((~&(wire1185 <= ((8'hac) >> $unsigned(wire1185)))) ?
                        (reg1081[(4'hb):(2'h2)] ?
                            (!$unsigned((reg1070 ?
                                reg1067 : wire1073))) : $signed(((wire1061 <= wire1061) ?
                                (wire1061 ?
                                    wire1188 : reg1069) : (~reg1070)))) : (($signed(wire1054[(4'hf):(4'ha)]) ?
                                (8'hb4) : $signed((-wire1055))) ?
                            $signed($signed((reg1079 ?
                                reg1074 : reg1078))) : wire1054));
  assign wire1191 = ({(-wire1090[(4'hf):(4'h9)])} > (-$unsigned(((reg1078 | wire1189) & reg1071[(2'h3):(1'h0)]))));
  assign wire1192 = $unsigned((^$unsigned(reg1069[(1'h0):(1'h0)])));
  assign wire1193 = $signed($unsigned($unsigned(reg1084[(2'h3):(2'h2)])));
  assign wire1194 = (!(reg1067[(4'hc):(1'h0)] > (wire1061 | ((reg1077 ?
                        reg1064 : reg1085) ^~ $unsigned((8'hb0))))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module831  (y, clk, wire832, wire833, wire834, wire835, wire836);
  output wire [(32'hdb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire832;
  input wire signed [(5'h11):(1'h0)] wire833;
  input wire signed [(5'h10):(1'h0)] wire834;
  input wire signed [(5'h10):(1'h0)] wire835;
  input wire signed [(4'hb):(1'h0)] wire836;
  reg [(4'hc):(1'h0)] reg1045 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1044 = (1'h0);
  reg [(4'hd):(1'h0)] reg1043 = (1'h0);
  reg [(5'h10):(1'h0)] reg1042 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1041 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1040 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1039 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1038 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1037 = (1'h0);
  reg [(2'h2):(1'h0)] reg1036 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1035 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire1034;
  wire [(4'hb):(1'h0)] wire1033;
  reg signed [(4'hb):(1'h0)] reg1032 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1031 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1030 = (1'h0);
  reg [(2'h3):(1'h0)] reg1029 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1028 = (1'h0);
  reg [(2'h2):(1'h0)] reg1027 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire1026;
  wire signed [(4'hd):(1'h0)] wire1025;
  wire signed [(5'h11):(1'h0)] wire948;
  wire [(4'h9):(1'h0)] wire1023;
  assign y = {reg1045,
                 reg1044,
                 reg1043,
                 reg1042,
                 reg1041,
                 reg1040,
                 reg1039,
                 reg1038,
                 reg1037,
                 reg1036,
                 reg1035,
                 wire1034,
                 wire1033,
                 reg1032,
                 reg1031,
                 reg1030,
                 reg1029,
                 reg1028,
                 reg1027,
                 wire1026,
                 wire1025,
                 wire948,
                 wire1023,
                 (1'h0)};
  module837 modinst949 (wire948, clk, wire835, wire834, wire836, wire833);
  module950 modinst1024 (wire1023, clk, wire832, wire836, wire833, wire948, wire835);
  assign wire1025 = (~|$unsigned($unsigned((wire948 ?
                        (wire833 <<< wire834) : wire836[(4'h8):(2'h2)]))));
  assign wire1026 = wire1025;
  always
    @(posedge clk) begin
      if ((-wire1023[(2'h2):(1'h0)]))
        begin
          if (wire1023[(3'h6):(3'h5)])
            begin
              reg1027 <= (^~((~|($unsigned(wire948) ?
                  wire833 : (wire1026 ? wire948 : (8'hbc)))) == (((wire834 ?
                      wire833 : wire948) ?
                  $unsigned(wire834) : $unsigned(wire836)) && ((wire834 <<< wire832) ?
                  wire833[(4'hb):(4'ha)] : ((8'ha4) ? wire1025 : wire1023)))));
              reg1028 <= (+wire834[(1'h0):(1'h0)]);
              reg1029 <= $signed((((~&reg1028) << (wire832[(3'h7):(3'h7)] || (~|wire835))) < {wire836[(4'h8):(1'h1)],
                  $unsigned($unsigned(wire1026))}));
            end
          else
            begin
              reg1027 <= $unsigned(wire832[(5'h12):(4'h8)]);
              reg1028 <= ((~|((reg1027 & (wire832 && (7'h40))) ?
                  $signed($signed((8'ha4))) : wire835)) <<< ((wire833 >> {{(8'hb0)}}) ?
                  (($signed(wire836) > $signed(wire1023)) | (~(reg1029 - wire835))) : reg1029));
              reg1029 <= wire1023[(1'h0):(1'h0)];
            end
          reg1030 <= {((!reg1028[(4'h9):(3'h7)]) > (7'h40))};
          reg1031 <= (~^wire1023);
          reg1032 <= wire832;
        end
      else
        begin
          reg1027 <= (wire1023 != reg1029[(2'h3):(1'h1)]);
          reg1028 <= wire948[(3'h7):(3'h4)];
          reg1029 <= reg1027;
        end
    end
  assign wire1033 = ((~|reg1029) ?
                        ({wire832,
                            $signed((~&wire1025))} ~^ wire1026[(3'h4):(1'h1)]) : (~(^((wire836 ?
                                (8'hb2) : reg1031) ?
                            $signed(wire836) : $unsigned(reg1029)))));
  assign wire1034 = wire832[(3'h6):(1'h1)];
  always
    @(posedge clk) begin
      if (($unsigned((&(!reg1029[(1'h1):(1'h0)]))) ^ $signed($unsigned((wire1026 ?
          reg1030 : (wire948 ? wire1033 : (7'h41)))))))
        begin
          reg1035 <= $unsigned($unsigned((($signed(wire832) <<< $signed(reg1027)) >= (wire948 ?
              $unsigned(wire836) : (reg1028 ? wire1034 : (7'h42))))));
          reg1036 <= (&$unsigned(wire1034[(1'h0):(1'h0)]));
          reg1037 <= $signed($signed((wire1033 >= (|(|wire833)))));
        end
      else
        begin
          reg1035 <= wire836[(4'h8):(4'h8)];
          if ((^{(reg1031[(4'h8):(3'h7)] >>> ($signed(wire1026) << (reg1031 * reg1032)))}))
            begin
              reg1036 <= (8'h9f);
            end
          else
            begin
              reg1036 <= (-($signed((reg1036[(1'h0):(1'h0)] + (reg1032 < reg1035))) ?
                  {(~wire1034[(2'h2):(2'h2)]),
                      $signed($unsigned(reg1028))} : wire835));
              reg1037 <= $signed(reg1031[(4'h9):(3'h7)]);
              reg1038 <= ($unsigned({reg1027[(2'h2):(1'h1)], (8'hb3)}) ?
                  reg1028[(4'h9):(3'h6)] : $unsigned(reg1035));
            end
          if (wire1026[(2'h3):(1'h0)])
            begin
              reg1039 <= (wire1034 - (~$signed(reg1035[(1'h0):(1'h0)])));
            end
          else
            begin
              reg1039 <= wire836[(3'h7):(1'h0)];
              reg1040 <= {({$signed((wire1023 ? reg1029 : wire948)),
                      reg1029[(2'h3):(1'h1)]} != ($unsigned((^reg1036)) ^~ wire834[(4'h8):(2'h2)]))};
              reg1041 <= {(~^$unsigned((reg1040[(1'h0):(1'h0)] ?
                      (reg1032 ? (8'ha6) : wire832) : reg1029[(1'h0):(1'h0)]))),
                  $signed((^((reg1032 >> (8'hae)) > $signed(wire836))))};
              reg1042 <= {($unsigned(($signed(wire836) ?
                      $unsigned(wire836) : (+wire834))) < $unsigned(reg1038))};
              reg1043 <= ($unsigned((^~(~|$signed(reg1030)))) ?
                  (^~((8'ha5) ?
                      (^(reg1029 != reg1029)) : $unsigned((wire1025 ?
                          reg1027 : (8'hbc))))) : (($signed($signed(wire948)) ?
                          $unsigned((~|reg1027)) : reg1035) ?
                      reg1040[(1'h1):(1'h0)] : $unsigned(wire1023)));
            end
        end
      reg1044 <= $unsigned(wire1023[(2'h3):(1'h1)]);
      reg1045 <= (+(((~&wire836) ?
              reg1040[(2'h3):(2'h3)] : $signed($signed(wire1026))) ?
          reg1043 : $unsigned((^~$signed(wire1034)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module950
#(parameter param1022 = (^{{(+(7'h41)), ((~|(8'ha1)) - {(8'h9f)})}}))
(y, clk, wire955, wire954, wire953, wire952, wire951);
  output wire [(32'h310):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire955;
  input wire signed [(4'hb):(1'h0)] wire954;
  input wire signed [(2'h2):(1'h0)] wire953;
  input wire signed [(5'h11):(1'h0)] wire952;
  input wire [(5'h10):(1'h0)] wire951;
  wire signed [(5'h15):(1'h0)] wire1021;
  reg [(4'hc):(1'h0)] reg1020 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1019 = (1'h0);
  reg [(4'h8):(1'h0)] reg1018 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1017 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1016 = (1'h0);
  reg [(5'h10):(1'h0)] reg1015 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1014 = (1'h0);
  reg [(2'h3):(1'h0)] reg1013 = (1'h0);
  reg [(4'h9):(1'h0)] reg1012 = (1'h0);
  reg [(5'h13):(1'h0)] reg1011 = (1'h0);
  reg [(4'hc):(1'h0)] reg1010 = (1'h0);
  reg [(5'h10):(1'h0)] reg1009 = (1'h0);
  reg [(2'h2):(1'h0)] reg1008 = (1'h0);
  reg [(4'h9):(1'h0)] reg1007 = (1'h0);
  reg [(4'hd):(1'h0)] reg1006 = (1'h0);
  reg [(4'hd):(1'h0)] reg1005 = (1'h0);
  reg [(4'hf):(1'h0)] reg1004 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1003 = (1'h0);
  reg [(3'h5):(1'h0)] reg1002 = (1'h0);
  reg [(5'h12):(1'h0)] reg1001 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1000 = (1'h0);
  reg [(3'h6):(1'h0)] reg999 = (1'h0);
  reg [(5'h11):(1'h0)] reg998 = (1'h0);
  reg [(5'h14):(1'h0)] reg997 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg996 = (1'h0);
  reg [(4'hb):(1'h0)] reg995 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg994 = (1'h0);
  reg [(5'h14):(1'h0)] reg993 = (1'h0);
  reg signed [(4'he):(1'h0)] reg992 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg991 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg990 = (1'h0);
  reg [(5'h14):(1'h0)] reg989 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg988 = (1'h0);
  reg [(4'ha):(1'h0)] reg987 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg986 = (1'h0);
  reg [(4'h8):(1'h0)] reg985 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg984 = (1'h0);
  reg [(4'h8):(1'h0)] reg983 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg982 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg981 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg980 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg979 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire978;
  wire [(2'h3):(1'h0)] wire977;
  wire signed [(5'h12):(1'h0)] wire976;
  wire signed [(2'h3):(1'h0)] wire975;
  reg [(5'h10):(1'h0)] reg974 = (1'h0);
  reg [(3'h4):(1'h0)] reg973 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg972 = (1'h0);
  reg [(5'h11):(1'h0)] reg971 = (1'h0);
  reg signed [(4'he):(1'h0)] reg970 = (1'h0);
  reg [(3'h7):(1'h0)] reg969 = (1'h0);
  reg [(5'h15):(1'h0)] reg968 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg967 = (1'h0);
  reg [(3'h5):(1'h0)] reg966 = (1'h0);
  reg [(3'h7):(1'h0)] reg965 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg964 = (1'h0);
  reg [(5'h14):(1'h0)] reg963 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg962 = (1'h0);
  reg [(4'h8):(1'h0)] reg961 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg960 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg959 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg958 = (1'h0);
  reg [(5'h13):(1'h0)] reg957 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg956 = (1'h0);
  assign y = {wire1021,
                 reg1020,
                 reg1019,
                 reg1018,
                 reg1017,
                 reg1016,
                 reg1015,
                 reg1014,
                 reg1013,
                 reg1012,
                 reg1011,
                 reg1010,
                 reg1009,
                 reg1008,
                 reg1007,
                 reg1006,
                 reg1005,
                 reg1004,
                 reg1003,
                 reg1002,
                 reg1001,
                 reg1000,
                 reg999,
                 reg998,
                 reg997,
                 reg996,
                 reg995,
                 reg994,
                 reg993,
                 reg992,
                 reg991,
                 reg990,
                 reg989,
                 reg988,
                 reg987,
                 reg986,
                 reg985,
                 reg984,
                 reg983,
                 reg982,
                 reg981,
                 reg980,
                 reg979,
                 wire978,
                 wire977,
                 wire976,
                 wire975,
                 reg974,
                 reg973,
                 reg972,
                 reg971,
                 reg970,
                 reg969,
                 reg968,
                 reg967,
                 reg966,
                 reg965,
                 reg964,
                 reg963,
                 reg962,
                 reg961,
                 reg960,
                 reg959,
                 reg958,
                 reg957,
                 reg956,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((wire951 + wire955[(2'h3):(1'h1)]))
        begin
          if (wire952[(5'h10):(3'h7)])
            begin
              reg956 <= (|wire952[(3'h6):(3'h4)]);
              reg957 <= wire954[(1'h0):(1'h0)];
            end
          else
            begin
              reg956 <= reg956;
              reg957 <= $unsigned($signed($signed(((wire953 > reg956) ?
                  $unsigned(reg957) : {wire952}))));
            end
          reg958 <= ({(wire953 != $unsigned(wire951[(1'h0):(1'h0)]))} ?
              wire953[(2'h2):(1'h0)] : wire951);
          reg959 <= $signed(((|(^~reg956)) * $unsigned((((8'hba) ?
              wire951 : wire951) && {wire953, wire953}))));
        end
      else
        begin
          reg956 <= wire955[(1'h0):(1'h0)];
          if ({({($signed(reg958) ~^ (wire955 + wire951)), (~(~|reg958))} ?
                  reg956[(2'h2):(1'h0)] : wire951[(3'h6):(3'h5)])})
            begin
              reg957 <= wire955[(2'h3):(1'h0)];
            end
          else
            begin
              reg957 <= wire952[(5'h10):(1'h1)];
              reg958 <= $unsigned((^$signed((|(wire953 ? (8'hbe) : wire954)))));
              reg959 <= (wire953 ^~ (wire953[(1'h0):(1'h0)] ?
                  $signed($unsigned({wire953,
                      reg959})) : wire953[(1'h1):(1'h1)]));
              reg960 <= {$signed($unsigned($unsigned($unsigned(reg956))))};
            end
          if ($signed(({$unsigned({wire955,
                  reg960})} >= $signed({(~^reg958)}))))
            begin
              reg961 <= $signed($unsigned(reg958[(5'h10):(4'hf)]));
              reg962 <= ((~|reg959[(2'h3):(2'h2)]) ?
                  ((8'hb5) >> ((~{(8'hbb)}) ?
                      (~|wire954) : (reg958[(4'hb):(2'h3)] || wire952[(4'ha):(4'ha)]))) : (wire952 < wire955));
              reg963 <= reg956[(3'h6):(3'h4)];
              reg964 <= $signed(((&(~$unsigned(wire954))) ?
                  wire955 : $unsigned($unsigned($unsigned(reg958)))));
            end
          else
            begin
              reg961 <= (wire954 ?
                  reg956 : (+($signed((wire954 < wire952)) != (|$unsigned(reg963)))));
              reg962 <= (reg962 ?
                  (wire955[(4'hc):(3'h7)] ?
                      $unsigned($unsigned(reg961)) : $unsigned((!reg958[(1'h1):(1'h0)]))) : ((($unsigned(reg961) ?
                              (-wire952) : (~^reg963)) ?
                          (-(^reg957)) : $unsigned({reg960})) ?
                      (-($unsigned(reg961) ?
                          (reg962 ?
                              reg962 : reg960) : $signed(reg956))) : wire955));
            end
          if (reg964)
            begin
              reg965 <= reg957[(2'h2):(2'h2)];
              reg966 <= $signed(wire952);
              reg967 <= (^~(reg962 ? (~&wire951[(1'h1):(1'h0)]) : reg960));
              reg968 <= (($signed((|((8'hb3) - reg967))) ?
                  (~^(^~(reg959 ?
                      reg963 : reg962))) : ($unsigned((reg961 | (8'hba))) & reg967[(5'h10):(3'h5)])) ^ (~|$signed($signed(reg967))));
            end
          else
            begin
              reg965 <= reg956;
              reg966 <= (+reg966);
              reg967 <= $unsigned(wire955[(1'h1):(1'h0)]);
              reg968 <= $unsigned(reg968);
              reg969 <= $unsigned((($unsigned({(8'haa),
                      reg956}) && (~&reg962)) ?
                  ((((8'haf) ? (8'ha0) : reg962) ?
                      $unsigned(reg965) : reg963) < reg964[(5'h11):(4'hc)]) : reg961));
            end
          reg970 <= $unsigned(wire954);
        end
      reg971 <= $unsigned({(-($signed(wire951) ? reg967 : reg970)),
          reg963[(1'h0):(1'h0)]});
      if ((((7'h42) >> $signed((+wire952))) ?
          $unsigned((8'ha1)) : $signed((8'hb0))))
        begin
          reg972 <= $unsigned((^$unsigned(reg970)));
          reg973 <= (^((reg962 * $unsigned($signed((8'ha8)))) ?
              ($signed((reg960 ? reg963 : (7'h43))) ?
                  ($signed((8'ha8)) ?
                      (reg966 ?
                          reg959 : reg962) : $signed(wire954)) : reg966) : (reg972[(3'h5):(1'h0)] ?
                  $unsigned((8'hb7)) : (reg958[(4'h8):(2'h3)] ^ (^~reg968)))));
          reg974 <= $signed((|$signed($signed(reg961))));
        end
      else
        begin
          reg972 <= $signed(((reg968[(3'h6):(2'h3)] ?
                  $signed((reg968 != (8'ha9))) : ((&reg958) ?
                      $signed(reg974) : $unsigned((8'ha6)))) ?
              $signed(($signed((8'hba)) >> (reg968 ~^ reg965))) : (8'ha5)));
          reg973 <= reg963;
          reg974 <= $unsigned($unsigned($signed($unsigned((~|(8'h9f))))));
        end
    end
  assign wire975 = reg965;
  assign wire976 = (|wire952);
  assign wire977 = wire955;
  assign wire978 = (^~({{wire955[(4'he):(1'h0)], $signed(reg959)},
                           ((reg957 ? reg962 : wire955) < reg958)} ?
                       reg964 : $unsigned($signed($unsigned((8'h9e))))));
  always
    @(posedge clk) begin
      if (wire951[(5'h10):(4'h9)])
        begin
          reg979 <= $signed({reg966, (&reg969)});
          reg980 <= ((wire976 ?
              (~|$unsigned(wire952)) : {$signed((reg956 ~^ reg973))}) != reg956);
          reg981 <= (reg974[(4'hd):(4'hc)] ?
              (wire952[(4'hf):(4'h8)] ?
                  reg965 : $unsigned($unsigned($signed(reg973)))) : {{$signed($signed((8'ha5)))}});
          if ({reg966[(2'h2):(1'h0)],
              (((~&$signed(reg957)) & ((^reg966) << reg980[(2'h2):(2'h2)])) ?
                  (reg967 ?
                      ((reg980 ? reg956 : reg966) ?
                          ((8'ha6) ?
                              reg959 : reg974) : (wire976 ~^ reg965)) : ((|wire951) ?
                          reg956 : $signed((8'hab)))) : $unsigned(((wire952 ~^ wire954) ?
                      $unsigned((8'ha1)) : {reg974, reg967})))})
            begin
              reg982 <= $unsigned((reg957[(2'h3):(1'h0)] ?
                  ((~&reg967[(1'h1):(1'h0)]) ~^ wire977) : $unsigned(($unsigned(wire975) > $unsigned(reg980)))));
              reg983 <= $signed(((reg971 ^~ $signed(((8'ha1) ?
                  wire951 : reg959))) >> (^~{$signed((8'hbd)),
                  reg959[(3'h5):(1'h1)]})));
            end
          else
            begin
              reg982 <= $signed((($unsigned(reg958[(2'h3):(2'h3)]) ?
                  wire953[(2'h2):(1'h0)] : ((-reg983) >>> wire953[(1'h0):(1'h0)])) || wire953));
              reg983 <= $unsigned({$signed(($signed((8'ha4)) - reg961)),
                  reg968});
              reg984 <= (8'haf);
              reg985 <= $unsigned(wire951);
            end
        end
      else
        begin
          if (wire951[(4'hd):(3'h5)])
            begin
              reg979 <= (~^wire951);
              reg980 <= (wire951 >> ((~&$signed((~|reg958))) ?
                  (((reg971 ? (8'ha8) : reg962) > reg969[(2'h2):(1'h1)]) ?
                      ((wire976 * reg984) + $unsigned(wire955)) : ($unsigned(reg980) ?
                          (reg956 >= reg962) : wire955)) : {wire978[(4'ha):(3'h5)]}));
            end
          else
            begin
              reg979 <= {($signed($unsigned(wire975[(1'h0):(1'h0)])) ?
                      reg963[(4'he):(3'h7)] : reg956[(1'h1):(1'h1)])};
              reg980 <= $signed(reg972);
            end
        end
      if ((((-$signed(wire977[(1'h0):(1'h0)])) ?
              (8'hac) : reg964[(4'hd):(4'hd)]) ?
          ((((reg966 <= wire975) ?
              {reg980} : (8'h9d)) ~^ (+$unsigned(reg971))) < {($unsigned(reg961) ?
                  (8'hbb) : (^reg980))}) : {reg956[(1'h1):(1'h1)],
              reg961[(3'h6):(2'h3)]}))
        begin
          reg986 <= ($unsigned((|(reg970 ?
              reg970[(4'ha):(3'h6)] : wire954))) ^~ reg967);
        end
      else
        begin
          reg986 <= $signed(reg968);
          reg987 <= reg964;
          reg988 <= reg979[(1'h1):(1'h0)];
          if ($signed((~^($unsigned(reg986) && reg963))))
            begin
              reg989 <= ($signed(((8'ha8) | $unsigned((reg968 ?
                  reg982 : reg988)))) | $unsigned((~|$unsigned(((8'ha2) != (8'hb4))))));
              reg990 <= {((wire978 ?
                      $unsigned((|wire953)) : $unsigned((wire955 ?
                          wire954 : wire952))) < reg972),
                  reg980};
              reg991 <= ((($unsigned($signed(reg982)) ^~ ((8'hae) ?
                      (reg989 | (8'h9f)) : reg969)) ?
                  reg985[(3'h6):(3'h5)] : ((^reg957) & (wire954 - reg981))) >= wire955);
            end
          else
            begin
              reg989 <= ($signed((wire954[(1'h0):(1'h0)] * $signed(reg963[(4'he):(3'h6)]))) & reg979[(1'h1):(1'h1)]);
            end
        end
      if (((reg981 ? (~$signed($unsigned(reg983))) : $unsigned(reg970)) ?
          ($signed(({reg967} ~^ {reg962})) ?
              reg991 : (reg985 ?
                  $unsigned($signed(reg979)) : wire975[(1'h0):(1'h0)])) : ((reg971[(4'hd):(3'h4)] && ((reg981 ?
              (8'hb0) : reg957) <= {(8'hbe),
              reg960})) ^ $signed($unsigned((~&reg964))))))
        begin
          if (($unsigned(($unsigned($unsigned((8'hbb))) ~^ ($signed(reg964) ~^ wire954))) ?
              (^~{(wire954[(4'hb):(1'h1)] <<< wire951[(3'h6):(1'h0)]),
                  (-wire952)}) : $unsigned(($signed((reg967 ?
                      reg990 : reg968)) ?
                  {(!reg973), $signed(reg960)} : $signed(reg988)))))
            begin
              reg992 <= reg957[(1'h0):(1'h0)];
            end
          else
            begin
              reg992 <= ($unsigned(($signed(reg968) != reg987[(2'h3):(2'h2)])) >= reg967);
              reg993 <= reg991;
              reg994 <= reg969;
            end
          if ((($signed(wire978[(4'h9):(2'h3)]) ?
                  $unsigned({$signed(wire976)}) : reg984[(3'h5):(2'h2)]) ?
              ((!$unsigned(reg960)) && wire953[(1'h0):(1'h0)]) : ($unsigned((~|reg987)) ?
                  ($signed($signed(reg967)) ^ ($unsigned(wire975) <= ((8'hb6) >= reg972))) : {((reg965 ?
                              reg981 : reg972) ?
                          $signed(reg972) : (+reg979)),
                      wire955})))
            begin
              reg995 <= (!{($signed(reg962[(1'h1):(1'h0)]) ?
                      wire975[(1'h0):(1'h0)] : $unsigned((reg973 ?
                          (8'haa) : (8'ha6))))});
              reg996 <= {(((8'ha4) ?
                          (~|{wire953}) : $unsigned(reg994[(1'h1):(1'h0)])) ?
                      $signed({$unsigned((7'h40)),
                          (~wire975)}) : $unsigned(reg972[(5'h11):(3'h5)]))};
            end
          else
            begin
              reg995 <= reg988[(1'h1):(1'h1)];
              reg996 <= {$signed((~&wire953))};
              reg997 <= ($unsigned(reg964) + $signed($signed({reg996,
                  (~|wire953)})));
              reg998 <= $signed(reg963[(4'hc):(3'h7)]);
              reg999 <= (^reg998[(4'hf):(4'hc)]);
            end
        end
      else
        begin
          reg992 <= reg960;
          reg993 <= (reg994[(3'h6):(3'h4)] ?
              $unsigned(reg993[(5'h11):(4'he)]) : wire951);
          if (($signed({reg973[(2'h3):(2'h3)], (~$signed(reg990))}) ?
              $signed(((reg988[(5'h11):(1'h1)] ?
                  reg968 : reg972) >> reg993[(4'hb):(1'h1)])) : ({($signed(reg979) ?
                      $signed((8'hae)) : (reg993 ?
                          reg988 : reg999))} - (&$signed(((8'haf) ?
                  (8'hb1) : reg958))))))
            begin
              reg994 <= $signed({$unsigned(($unsigned(reg988) ?
                      $unsigned(wire975) : (reg962 >= reg979))),
                  reg966[(1'h0):(1'h0)]});
              reg995 <= (^~$unsigned((reg967 << (8'hac))));
            end
          else
            begin
              reg994 <= reg956[(1'h0):(1'h0)];
              reg995 <= (|($unsigned(reg970) ?
                  $unsigned((wire951 ?
                      $signed(reg997) : (reg985 | (8'had)))) : $signed((-$signed(reg959)))));
              reg996 <= $unsigned((($signed((reg963 ?
                      reg990 : reg964)) <= (reg966 > $signed(reg999))) ?
                  ($unsigned((^~reg988)) ?
                      (reg974[(3'h4):(3'h4)] ?
                          $unsigned(reg987) : wire975[(1'h0):(1'h0)]) : reg995) : $unsigned((reg994 ?
                      {reg992} : (!wire975)))));
              reg997 <= $signed(($signed(((~&reg967) > wire977[(2'h3):(1'h1)])) || $signed((~&reg995[(4'h8):(3'h7)]))));
            end
        end
      reg1000 <= $unsigned((reg969[(3'h4):(1'h1)] ?
          $unsigned($signed(reg991[(2'h3):(2'h2)])) : (~^($unsigned(reg984) == reg980))));
    end
  always
    @(posedge clk) begin
      reg1001 <= $signed((^$unsigned($unsigned($unsigned(reg967)))));
      if ({(((~|$unsigned((8'ha8))) == reg982[(2'h3):(2'h3)]) ?
              {(~$signed(reg984))} : reg1001[(4'ha):(3'h7)])})
        begin
          if (($signed(($unsigned((8'hb6)) | (~|reg996))) >= reg989))
            begin
              reg1002 <= ((^~reg995[(4'ha):(3'h6)]) && (^~(({reg957} >> (reg987 ?
                      reg964 : reg972)) ?
                  reg979 : (reg964 >= reg967[(2'h3):(2'h3)]))));
              reg1003 <= reg992;
              reg1004 <= reg983[(3'h4):(1'h1)];
            end
          else
            begin
              reg1002 <= ($signed((~reg958[(4'he):(4'h9)])) + (^reg967));
              reg1003 <= reg979;
            end
          reg1005 <= {(!(wire977 >>> $signed((reg994 ? wire977 : reg989)))),
              (+(8'h9f))};
        end
      else
        begin
          reg1002 <= ($signed($unsigned($signed(((8'hb6) ?
                  wire951 : reg990)))) ?
              reg993[(2'h2):(1'h0)] : wire952);
          if (((reg986 ? $unsigned(reg969[(2'h3):(1'h1)]) : (~&reg968)) ?
              $signed((8'hae)) : $signed(reg998[(3'h5):(2'h2)])))
            begin
              reg1003 <= (($signed(wire953) ?
                      (reg957 ?
                          $unsigned(reg1002[(3'h4):(1'h1)]) : ($signed(reg961) <<< wire952)) : reg967[(3'h4):(1'h0)]) ?
                  wire954[(4'h9):(1'h1)] : reg968[(5'h13):(4'hd)]);
              reg1004 <= (!wire954[(2'h3):(2'h3)]);
              reg1005 <= $unsigned($unsigned(reg993));
              reg1006 <= (+(~reg972[(3'h5):(1'h1)]));
            end
          else
            begin
              reg1003 <= ((8'hbd) ? (~(^(8'ha3))) : reg988);
              reg1004 <= reg979;
              reg1005 <= $signed(reg992);
              reg1006 <= (reg964 ?
                  reg956 : (!$unsigned((reg1004 ?
                      (reg1003 * wire978) : reg995))));
              reg1007 <= $unsigned(({(~&reg991[(2'h3):(1'h1)])} != $unsigned({$unsigned((8'had)),
                  (wire955 - reg988)})));
            end
          reg1008 <= (($signed(($unsigned(reg979) <= ((8'ha4) > wire976))) ?
              reg990 : (reg1001 <<< $unsigned($unsigned(wire953)))) + ($unsigned($unsigned(reg981)) ?
              $unsigned(reg959) : reg959));
          if (($signed({wire953[(1'h1):(1'h1)],
                  ({reg965} - reg990[(1'h1):(1'h1)])}) ?
              wire952[(3'h4):(2'h2)] : reg1008[(1'h1):(1'h0)]))
            begin
              reg1009 <= (|$unsigned($signed(reg992)));
              reg1010 <= $signed(((+((reg997 ^ reg987) || $unsigned(reg969))) | ($unsigned((reg960 >>> reg956)) == (((8'hbc) ?
                      reg1005 : reg1007) ?
                  $signed((8'h9d)) : reg956[(3'h4):(3'h4)]))));
              reg1011 <= (reg1005 ?
                  (&((reg1004 ?
                      $unsigned(reg959) : $unsigned(reg963)) ~^ (!reg982[(1'h1):(1'h0)]))) : ((reg994 ?
                      (((8'haf) ? reg969 : reg987) ?
                          {reg971,
                              reg987} : reg974) : reg980[(4'h8):(3'h5)]) >> $signed($signed((~&reg970)))));
            end
          else
            begin
              reg1009 <= $unsigned(wire976[(3'h5):(1'h1)]);
              reg1010 <= {((8'hbe) < (((reg971 ?
                      reg1005 : reg963) ^~ reg994[(2'h3):(1'h1)]) << (((8'ha8) ?
                      reg985 : reg1000) >>> reg997)))};
              reg1011 <= $unsigned(((reg984[(2'h3):(1'h0)] ?
                  wire977 : ((reg982 < (8'hbb)) <<< $signed(reg979))) ^ $unsigned(((reg999 ?
                      wire952 : (8'ha1)) ?
                  (reg994 ? (8'hb9) : reg1008) : reg995[(3'h5):(3'h5)]))));
              reg1012 <= (7'h42);
              reg1013 <= $signed($signed((+reg979[(1'h0):(1'h0)])));
            end
          reg1014 <= $unsigned($unsigned((8'had)));
        end
      if (((!{reg959[(1'h0):(1'h0)]}) && reg958[(4'ha):(2'h2)]))
        begin
          reg1015 <= (($unsigned($unsigned({reg987,
              reg1003})) & reg1001) < ($signed(($unsigned(reg964) ^~ $unsigned(wire977))) ^ reg982[(1'h0):(1'h0)]));
          reg1016 <= {reg959, wire952[(4'hc):(2'h2)]};
          reg1017 <= reg983[(1'h1):(1'h0)];
          reg1018 <= {$unsigned(reg1005[(3'h7):(2'h2)])};
        end
      else
        begin
          if (($signed((!{$signed(reg1016)})) - (reg972[(5'h15):(5'h12)] ?
              $signed(($unsigned(reg962) ?
                  (reg1002 ?
                      wire975 : reg967) : reg971[(4'h8):(2'h2)])) : {((^~reg964) - (reg1013 ?
                      reg965 : (8'hac)))})))
            begin
              reg1015 <= ((+((^reg1018[(2'h2):(1'h0)]) <= $unsigned(reg969))) ?
                  (reg995[(2'h3):(2'h2)] > (|((reg995 <<< reg972) <= (8'ha8)))) : (({reg993[(3'h4):(1'h1)]} >> $signed(((8'h9e) ?
                      reg958 : reg988))) == $signed($unsigned($unsigned((8'hb3))))));
              reg1016 <= (reg1008[(2'h2):(2'h2)] ?
                  (reg995[(4'hb):(3'h7)] <= $unsigned($signed((reg992 ?
                      reg994 : reg957)))) : $signed((reg970 < (~&$signed(reg991)))));
              reg1017 <= (($signed(((~reg1007) ? (-reg966) : {reg971})) ?
                  (8'ha5) : (reg988[(4'h8):(1'h1)] ?
                      reg1008[(1'h1):(1'h0)] : ((~|reg994) > (reg983 ?
                          wire978 : wire952)))) ^ (reg972 ?
                  $signed({(reg1000 ?
                          (8'hb6) : (7'h43))}) : $unsigned((8'hbc))));
              reg1018 <= ($signed($unsigned($signed($unsigned(reg984)))) | (reg964 ?
                  {(8'hbd), $signed($signed(reg1016))} : {(((8'ha0) ?
                          reg986 : reg968) != $signed(reg1015)),
                      reg992[(4'ha):(2'h3)]}));
            end
          else
            begin
              reg1015 <= {(({$unsigned(reg983),
                      reg969[(3'h6):(3'h6)]} >> ($unsigned(reg981) ?
                      reg1005 : (7'h40))) >= reg959),
                  ($unsigned(($unsigned(reg970) ?
                          reg985[(4'h8):(3'h6)] : $signed(wire955))) ?
                      reg984 : (reg961[(2'h3):(1'h0)] && $unsigned((reg983 ?
                          reg974 : wire953))))};
              reg1016 <= $unsigned(reg973[(2'h3):(2'h2)]);
              reg1017 <= $signed((($signed($unsigned(reg1013)) << $unsigned($unsigned(reg990))) ?
                  reg980[(4'h8):(1'h1)] : $unsigned({$unsigned((8'hb1)),
                      (reg990 >> reg983)})));
              reg1018 <= $signed((~(~|reg1018)));
              reg1019 <= (!{$unsigned($signed($signed(reg1012))), (^reg1008)});
            end
        end
      reg1020 <= $unsigned((8'hab));
    end
  assign wire1021 = $unsigned({$signed($signed((&reg957)))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module837  (y, clk, wire841, wire840, wire839, wire838);
  output wire [(32'h4b0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire841;
  input wire [(5'h10):(1'h0)] wire840;
  input wire [(2'h2):(1'h0)] wire839;
  input wire [(5'h11):(1'h0)] wire838;
  wire signed [(4'ha):(1'h0)] wire947;
  wire signed [(5'h13):(1'h0)] wire946;
  reg signed [(5'h10):(1'h0)] reg945 = (1'h0);
  reg [(4'ha):(1'h0)] reg944 = (1'h0);
  reg [(4'hf):(1'h0)] reg943 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg942 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg941 = (1'h0);
  reg [(4'hf):(1'h0)] reg940 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg939 = (1'h0);
  reg [(5'h14):(1'h0)] reg938 = (1'h0);
  reg [(5'h10):(1'h0)] reg937 = (1'h0);
  reg [(5'h11):(1'h0)] reg936 = (1'h0);
  reg [(5'h12):(1'h0)] reg935 = (1'h0);
  reg [(4'h8):(1'h0)] reg934 = (1'h0);
  reg signed [(4'he):(1'h0)] reg933 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg932 = (1'h0);
  reg [(4'hb):(1'h0)] reg931 = (1'h0);
  reg [(4'he):(1'h0)] reg930 = (1'h0);
  reg [(4'h8):(1'h0)] reg929 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg928 = (1'h0);
  reg [(4'h8):(1'h0)] reg927 = (1'h0);
  reg [(3'h5):(1'h0)] reg926 = (1'h0);
  reg [(3'h5):(1'h0)] reg925 = (1'h0);
  reg [(4'h8):(1'h0)] reg924 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg923 = (1'h0);
  reg [(4'hf):(1'h0)] reg922 = (1'h0);
  reg [(4'h9):(1'h0)] reg921 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg920 = (1'h0);
  reg [(4'h8):(1'h0)] reg919 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg918 = (1'h0);
  reg [(2'h3):(1'h0)] reg917 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg916 = (1'h0);
  reg [(5'h13):(1'h0)] reg915 = (1'h0);
  reg [(3'h5):(1'h0)] reg914 = (1'h0);
  reg [(4'h8):(1'h0)] reg913 = (1'h0);
  reg [(3'h4):(1'h0)] reg912 = (1'h0);
  reg [(4'h8):(1'h0)] reg911 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg910 = (1'h0);
  reg [(5'h13):(1'h0)] reg909 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg908 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg907 = (1'h0);
  reg [(5'h14):(1'h0)] reg906 = (1'h0);
  reg [(3'h4):(1'h0)] reg905 = (1'h0);
  reg [(2'h2):(1'h0)] reg904 = (1'h0);
  reg [(5'h15):(1'h0)] reg903 = (1'h0);
  reg [(4'h8):(1'h0)] reg902 = (1'h0);
  reg [(5'h11):(1'h0)] reg901 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg899 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg898 = (1'h0);
  reg [(4'hc):(1'h0)] reg897 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg896 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg895 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg894 = (1'h0);
  reg [(4'hb):(1'h0)] reg893 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg892 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg891 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg890 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg889 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg888 = (1'h0);
  reg [(4'hc):(1'h0)] reg887 = (1'h0);
  reg [(4'he):(1'h0)] reg886 = (1'h0);
  wire [(4'hf):(1'h0)] wire885;
  wire [(5'h10):(1'h0)] wire884;
  wire signed [(3'h6):(1'h0)] wire883;
  wire [(4'h8):(1'h0)] wire882;
  reg signed [(4'h8):(1'h0)] reg881 = (1'h0);
  reg [(4'ha):(1'h0)] reg880 = (1'h0);
  reg [(3'h6):(1'h0)] reg879 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg878 = (1'h0);
  reg [(2'h2):(1'h0)] reg877 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg876 = (1'h0);
  reg [(4'hd):(1'h0)] reg875 = (1'h0);
  reg [(2'h2):(1'h0)] reg874 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg873 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg872 = (1'h0);
  reg [(3'h5):(1'h0)] reg871 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg870 = (1'h0);
  reg [(3'h4):(1'h0)] reg869 = (1'h0);
  reg [(3'h4):(1'h0)] reg868 = (1'h0);
  reg [(5'h11):(1'h0)] reg867 = (1'h0);
  reg [(4'he):(1'h0)] reg866 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg865 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg864 = (1'h0);
  reg [(3'h7):(1'h0)] reg863 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg862 = (1'h0);
  reg [(4'h8):(1'h0)] reg861 = (1'h0);
  wire signed [(4'he):(1'h0)] wire860;
  wire signed [(3'h6):(1'h0)] wire859;
  reg signed [(4'h9):(1'h0)] reg858 = (1'h0);
  reg [(4'hb):(1'h0)] reg857 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg856 = (1'h0);
  reg [(5'h15):(1'h0)] reg855 = (1'h0);
  reg [(2'h2):(1'h0)] reg854 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg853 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire852;
  reg signed [(4'hb):(1'h0)] reg851 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg850 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg849 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg848 = (1'h0);
  reg [(5'h12):(1'h0)] reg847 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg846 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg845 = (1'h0);
  reg [(4'h8):(1'h0)] reg844 = (1'h0);
  reg [(3'h4):(1'h0)] reg843 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire842;
  assign y = {wire947,
                 wire946,
                 reg945,
                 reg944,
                 reg943,
                 reg942,
                 reg941,
                 reg940,
                 reg939,
                 reg938,
                 reg937,
                 reg936,
                 reg935,
                 reg934,
                 reg933,
                 reg932,
                 reg931,
                 reg930,
                 reg929,
                 reg928,
                 reg927,
                 reg926,
                 reg925,
                 reg924,
                 reg923,
                 reg922,
                 reg921,
                 reg920,
                 reg919,
                 reg918,
                 reg917,
                 reg916,
                 reg915,
                 reg914,
                 reg913,
                 reg912,
                 reg911,
                 reg910,
                 reg909,
                 reg908,
                 reg907,
                 reg906,
                 reg905,
                 reg904,
                 reg903,
                 reg902,
                 reg901,
                 reg900,
                 reg899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 reg893,
                 reg892,
                 reg891,
                 reg890,
                 reg889,
                 reg888,
                 reg887,
                 reg886,
                 wire885,
                 wire884,
                 wire883,
                 wire882,
                 reg881,
                 reg880,
                 reg879,
                 reg878,
                 reg877,
                 reg876,
                 reg875,
                 reg874,
                 reg873,
                 reg872,
                 reg871,
                 reg870,
                 reg869,
                 reg868,
                 reg867,
                 reg866,
                 reg865,
                 reg864,
                 reg863,
                 reg862,
                 reg861,
                 wire860,
                 wire859,
                 reg858,
                 reg857,
                 reg856,
                 reg855,
                 reg854,
                 reg853,
                 wire852,
                 reg851,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 reg846,
                 reg845,
                 reg844,
                 reg843,
                 wire842,
                 (1'h0)};
  assign wire842 = $unsigned(($unsigned(wire841) ?
                       ((wire840[(4'h8):(3'h5)] & $signed(wire839)) ?
                           $unsigned(wire841[(4'hb):(3'h6)]) : ($signed((8'h9f)) ?
                               $signed((8'hbd)) : (wire839 ?
                                   (8'hb3) : wire841))) : ((wire840[(4'hd):(4'ha)] ?
                               $signed(wire841) : wire839) ?
                           ($unsigned(wire839) ?
                               $signed(wire838) : (^wire841)) : wire839)));
  always
    @(posedge clk) begin
      reg843 <= $unsigned((wire839 ?
          (7'h43) : $signed(($signed((8'ha3)) ?
              wire842[(4'hf):(3'h5)] : wire839))));
      reg844 <= {(wire842 ?
              (^$signed({wire838})) : $unsigned($signed((wire840 ?
                  (8'hbc) : wire842)))),
          $signed(wire838[(5'h11):(1'h1)])};
      if ({((+(wire841 ?
                  (wire842 ? wire841 : reg843) : (wire842 ?
                      wire839 : wire842))) ?
              $signed(($unsigned(reg844) << wire841)) : $signed(wire842))})
        begin
          reg845 <= (!wire839);
        end
      else
        begin
          reg845 <= $signed(((($signed(wire839) > {wire842, reg844}) ?
                  (^wire839[(1'h1):(1'h0)]) : $unsigned(wire842)) ?
              ($unsigned($unsigned(wire840)) != ((-wire839) ?
                  ((8'h9f) ~^ wire841) : wire842)) : $unsigned((wire839[(1'h0):(1'h0)] + (&wire839)))));
          if ($signed(reg845))
            begin
              reg846 <= (!(((reg845 ^ (8'ha1)) >> wire842) ?
                  (!({reg843, (8'h9e)} | (~|wire841))) : wire841));
              reg847 <= wire842;
              reg848 <= $signed({{(8'hbc), reg847}});
            end
          else
            begin
              reg846 <= reg845[(3'h7):(2'h2)];
              reg847 <= reg844[(1'h0):(1'h0)];
              reg848 <= $unsigned((8'ha7));
            end
          reg849 <= $unsigned((-wire841));
          reg850 <= $unsigned(wire839);
        end
      reg851 <= {((reg846[(1'h1):(1'h1)] ? {$unsigned(reg849)} : reg845) ?
              wire842[(4'h8):(2'h2)] : (~(wire839[(1'h0):(1'h0)] ?
                  $signed(wire840) : $signed(reg847)))),
          ($unsigned(wire841) != $signed({$signed(reg844)}))};
    end
  assign wire852 = $signed($signed(((wire840[(4'hc):(1'h0)] ?
                       {reg848} : (reg851 ?
                           reg844 : wire839)) & ($unsigned(reg844) || $unsigned(reg848)))));
  always
    @(posedge clk) begin
      if (wire838[(4'hc):(3'h6)])
        begin
          reg853 <= (+$signed({(&$signed(reg851))}));
          reg854 <= $unsigned({reg847});
        end
      else
        begin
          reg853 <= $signed(reg854);
          if (reg848[(1'h1):(1'h1)])
            begin
              reg854 <= reg854[(2'h2):(1'h1)];
              reg855 <= reg853[(3'h6):(2'h2)];
              reg856 <= ($unsigned(reg851) ?
                  $signed($unsigned(((~(8'hb7)) ?
                      {wire840,
                          wire840} : $unsigned(reg851)))) : $signed($unsigned(($unsigned(wire841) ?
                      (reg853 + wire838) : (!(7'h41))))));
            end
          else
            begin
              reg854 <= (~&(~($signed(reg845[(3'h5):(2'h2)]) ?
                  wire839[(1'h1):(1'h0)] : {(reg849 ? reg849 : reg848),
                      (8'hbe)})));
            end
        end
      reg857 <= $signed((!({$signed(reg855), {reg849, reg844}} ?
          (reg845 <<< (^reg856)) : (8'hb1))));
      reg858 <= reg847;
    end
  assign wire859 = (((^reg856[(4'hb):(3'h7)]) ?
                       wire840 : (reg854[(1'h0):(1'h0)] | $unsigned((~|wire852)))) | $unsigned(($unsigned(wire838) & ($unsigned(wire841) ?
                       (wire852 | reg858) : reg845[(3'h4):(1'h1)]))));
  assign wire860 = wire859;
  always
    @(posedge clk) begin
      if ($signed($unsigned(wire839[(1'h1):(1'h0)])))
        begin
          reg861 <= (^reg853[(1'h1):(1'h0)]);
          reg862 <= $unsigned($unsigned((($unsigned(reg849) <= wire852[(3'h5):(3'h4)]) ~^ reg846)));
          if ($signed((reg854[(1'h1):(1'h1)] * reg851)))
            begin
              reg863 <= (reg849 != (reg850 ? reg847 : reg844));
              reg864 <= ($signed($signed((|$unsigned(wire840)))) != (wire839 == $signed($signed((~^reg862)))));
              reg865 <= (({($signed((8'h9d)) >= $unsigned(wire859)),
                      reg854[(1'h0):(1'h0)]} ?
                  (^((reg854 <<< wire842) ?
                      wire838[(4'he):(4'ha)] : wire852)) : (((reg854 - reg853) ?
                      reg849 : (^~wire842)) > reg856[(5'h10):(4'ha)])) >>> ($signed(reg858[(1'h1):(1'h0)]) ?
                  wire840 : reg856[(2'h2):(1'h1)]));
            end
          else
            begin
              reg863 <= {$signed($signed(reg851)),
                  (reg847[(2'h3):(1'h1)] ?
                      $unsigned(reg857[(1'h0):(1'h0)]) : (8'ha2))};
              reg864 <= reg855;
              reg865 <= $unsigned($unsigned((~&{(~&reg846), wire859})));
              reg866 <= reg854[(1'h0):(1'h0)];
              reg867 <= ($signed(((reg850[(3'h6):(1'h0)] <= reg850[(3'h4):(1'h1)]) && reg861)) >= (8'h9f));
            end
        end
      else
        begin
          reg861 <= $unsigned(reg863);
          if (reg853)
            begin
              reg862 <= wire842;
            end
          else
            begin
              reg862 <= reg845;
              reg863 <= (+(8'had));
              reg864 <= (($signed(reg867) && wire840) >= (|$signed(($unsigned(reg856) >>> reg843))));
              reg865 <= {reg844,
                  {$signed(((reg849 ? reg850 : reg853) ?
                          (reg847 | reg853) : $unsigned(reg850)))}};
            end
          reg866 <= (+$signed($unsigned(reg855)));
          reg867 <= reg866;
          if ($unsigned($signed((8'ha9))))
            begin
              reg868 <= reg857;
              reg869 <= (^~wire860);
              reg870 <= reg868[(1'h0):(1'h0)];
              reg871 <= $unsigned({(reg862 > (^reg846[(4'hf):(4'hc)])),
                  $unsigned($unsigned($unsigned(wire840)))});
              reg872 <= {(reg865 ^ (~&reg847[(5'h10):(4'hc)])), reg855};
            end
          else
            begin
              reg868 <= reg865;
              reg869 <= (|wire841);
              reg870 <= $signed($unsigned((-reg872)));
            end
        end
      reg873 <= $unsigned(reg847[(4'hd):(3'h6)]);
      reg874 <= reg848;
    end
  always
    @(posedge clk) begin
      if ((&wire838[(4'ha):(2'h2)]))
        begin
          reg875 <= ($unsigned($unsigned((reg874[(2'h2):(1'h1)] || reg874))) ~^ wire860);
          reg876 <= reg871;
          reg877 <= $signed((reg876 ?
              $signed(reg858) : $signed(((~&wire839) ?
                  $signed(reg876) : (+reg875)))));
          reg878 <= ((7'h44) & (&wire841[(2'h3):(1'h0)]));
          if ($signed((8'ha8)))
            begin
              reg879 <= reg858[(3'h5):(3'h4)];
              reg880 <= ($signed((~&$signed($unsigned(reg875)))) ?
                  (reg863[(3'h4):(2'h3)] >= $unsigned(reg862)) : $signed(($signed(reg865) ^~ $signed($signed(reg863)))));
              reg881 <= ({(8'ha1)} ? reg875[(1'h1):(1'h1)] : wire840);
            end
          else
            begin
              reg879 <= $unsigned($unsigned(($signed((8'hb2)) ^~ reg844[(3'h4):(1'h1)])));
              reg880 <= $unsigned(reg857[(1'h1):(1'h0)]);
              reg881 <= {$signed($signed((&(reg869 ? (8'hba) : (8'hb7)))))};
            end
        end
      else
        begin
          reg875 <= $signed(($signed(reg870[(1'h0):(1'h0)]) ?
              $unsigned(($unsigned(reg874) ~^ reg862[(4'hb):(1'h0)])) : reg855));
          if ($unsigned($unsigned($signed(reg845))))
            begin
              reg876 <= (^~(((~(wire841 >= (8'hac))) ?
                      (reg863 && reg871) : $signed({(8'hbf)})) ?
                  (reg851 ? $signed((|reg864)) : $signed(reg865)) : reg866));
              reg877 <= reg872;
              reg878 <= (reg879 ?
                  reg862[(1'h0):(1'h0)] : (reg877[(2'h2):(2'h2)] - ({$unsigned(reg870),
                      $unsigned(reg854)} << reg866[(4'ha):(3'h5)])));
              reg879 <= {reg847, reg881};
            end
          else
            begin
              reg876 <= {$signed($unsigned($signed(wire838)))};
              reg877 <= reg854[(2'h2):(1'h0)];
            end
          reg880 <= ($signed((-($signed((8'h9c)) ?
                  (8'ha2) : reg856[(5'h13):(3'h4)]))) ?
              ($unsigned(($signed((8'ha1)) ^~ (reg881 ?
                  reg856 : reg844))) != (8'ha5)) : {(-$signed({reg849}))});
        end
    end
  assign wire882 = (((+((wire840 ? wire852 : reg862) ?
                           reg869[(2'h3):(1'h0)] : reg875)) ?
                       (((&reg878) ?
                               $signed(wire852) : (wire839 ? reg876 : reg864)) ?
                           (~{reg862,
                               reg877}) : (~&reg850)) : reg874[(2'h2):(2'h2)]) ~^ reg871);
  assign wire883 = wire882;
  assign wire884 = $unsigned(reg857[(4'h8):(4'h8)]);
  assign wire885 = wire839[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      if ($signed({wire839}))
        begin
          reg886 <= reg879;
          reg887 <= $signed((+{reg857[(3'h6):(1'h1)]}));
          reg888 <= $signed($signed({($unsigned((8'hba)) ?
                  (^(8'ha7)) : reg876[(2'h2):(2'h2)])}));
          if ((!$unsigned(({reg869, $unsigned(wire885)} ?
              (^reg876) : reg858[(2'h3):(2'h3)]))))
            begin
              reg889 <= reg866;
              reg890 <= $signed({reg843, (8'hae)});
              reg891 <= (!$unsigned({((reg855 ?
                      reg866 : reg887) | (&reg846))}));
              reg892 <= ((^(reg866 & $signed((~reg871)))) ?
                  (8'hb4) : ($signed(wire838[(1'h1):(1'h1)]) >= (^$unsigned((~&(8'hbf))))));
              reg893 <= $signed((~($signed(reg891[(1'h0):(1'h0)]) ?
                  (~$signed((8'hab))) : {{reg880, (7'h40)}})));
            end
          else
            begin
              reg889 <= (~&reg870[(1'h0):(1'h0)]);
              reg890 <= {(8'hb1), (-$unsigned({reg868}))};
            end
        end
      else
        begin
          if (((($unsigned((reg867 ? (8'hb5) : reg868)) ?
                  reg851[(2'h3):(1'h1)] : (~&(reg865 - (8'ha1)))) ?
              ($signed(((8'hbf) <<< reg876)) ?
                  ((|reg862) + reg872[(1'h1):(1'h1)]) : reg857) : reg857) - ((reg880 ?
                  ({reg880, wire852} ?
                      (reg844 ?
                          wire860 : reg854) : $signed((8'haf))) : reg855) ?
              {($unsigned(reg844) * reg889[(1'h1):(1'h0)]),
                  reg865} : (|(-(reg850 ? reg854 : reg864))))))
            begin
              reg886 <= $signed($signed({$signed({reg858})}));
              reg887 <= $signed(wire841);
              reg888 <= (8'ha4);
            end
          else
            begin
              reg886 <= {$unsigned(reg891[(1'h1):(1'h0)]),
                  $unsigned((~|$signed((-(8'haa)))))};
              reg887 <= {{(^$signed(wire838)), $signed(reg845)},
                  ((($unsigned(reg877) && $unsigned((8'ha7))) ?
                          ($signed(reg856) ?
                              wire884 : (reg846 << reg881)) : $signed($signed((8'ha9)))) ?
                      wire852[(2'h3):(2'h2)] : wire882[(3'h5):(3'h4)])};
              reg888 <= ($signed((wire842[(4'ha):(3'h6)] + $signed(reg893))) ?
                  $signed({$unsigned((~reg863)),
                      (wire841[(4'hb):(1'h0)] <= (~&reg847))}) : reg849);
              reg889 <= reg863[(2'h3):(1'h0)];
            end
          reg890 <= reg865;
          if ($unsigned($unsigned(reg892[(3'h6):(1'h0)])))
            begin
              reg891 <= ((((7'h41) & (((8'h9c) ? reg868 : reg849) ?
                      $unsigned(reg874) : $unsigned(reg873))) >>> ($unsigned((reg845 ?
                      reg853 : (8'hb0))) + reg892[(1'h1):(1'h0)])) ?
                  $signed((((reg878 ? reg849 : wire842) + (+(7'h40))) ?
                      (~^reg861[(2'h2):(1'h0)]) : ({reg861} ?
                          (reg868 >> reg871) : reg856[(5'h11):(3'h7)]))) : (reg857[(3'h5):(1'h0)] ?
                      reg890[(2'h2):(1'h0)] : $signed((|(reg889 ?
                          (8'had) : reg868)))));
              reg892 <= (($signed({$signed(reg857)}) ?
                  reg843[(2'h3):(2'h3)] : ($unsigned((reg877 ?
                          reg850 : reg858)) ?
                      (wire838[(2'h3):(2'h2)] ?
                          reg872[(1'h1):(1'h1)] : wire842) : reg886[(4'he):(4'h9)])) << wire842[(3'h4):(2'h2)]);
              reg893 <= wire882[(1'h1):(1'h0)];
            end
          else
            begin
              reg891 <= ((8'hbb) ?
                  (~|$unsigned((reg851[(4'h9):(3'h7)] > $unsigned(reg854)))) : (reg855[(5'h11):(1'h0)] & wire841));
              reg892 <= reg880[(3'h6):(3'h5)];
              reg893 <= ($signed($unsigned($unsigned(reg874))) || reg861[(1'h1):(1'h1)]);
            end
          reg894 <= (reg857[(3'h4):(1'h0)] ?
              reg863[(1'h0):(1'h0)] : ({{$unsigned(reg874)}} == ($unsigned(reg886) ?
                  reg889 : ($signed(reg889) >= $unsigned(wire838)))));
        end
      if (reg876[(4'hb):(2'h3)])
        begin
          reg895 <= (reg874 >= {reg891[(1'h0):(1'h0)], $signed(reg854)});
          reg896 <= $signed({(wire841[(4'hd):(4'h8)] ?
                  ({wire852,
                      reg875} == wire839[(1'h1):(1'h1)]) : $unsigned({(8'hbf),
                      reg894}))});
          if (($unsigned(reg881[(3'h7):(2'h2)]) ?
              (reg862 * (&(wire883[(1'h0):(1'h0)] && (reg846 ?
                  reg887 : reg846)))) : ((($unsigned(reg875) <= ((8'ha2) == reg880)) ?
                  {(reg847 ? wire838 : reg888), $signed((7'h41))} : ((wire859 ?
                      reg896 : reg865) + $signed(wire883))) ^~ ({$signed(reg863),
                  reg858} >> reg864[(2'h2):(1'h1)]))))
            begin
              reg897 <= (reg869[(1'h0):(1'h0)] ?
                  ((reg847 + $unsigned(reg871[(2'h3):(1'h0)])) || (reg844 > $signed($unsigned(reg864)))) : wire860[(4'hc):(3'h5)]);
              reg898 <= (reg889[(2'h3):(2'h2)] != ($signed($signed((reg845 && (7'h43)))) ?
                  (((7'h42) >= (|reg856)) ?
                      (reg849 ?
                          (reg892 ?
                              reg873 : reg851) : $signed((8'hb3))) : (8'haa)) : (&($unsigned((8'haf)) ?
                      $unsigned(reg869) : $signed((8'hae))))));
              reg899 <= (-$signed((~((reg887 ?
                  reg867 : wire859) >> $signed(wire839)))));
              reg900 <= (~^(-$unsigned($signed(reg887))));
              reg901 <= (|$unsigned(($signed($unsigned(reg866)) < reg890[(3'h5):(1'h0)])));
            end
          else
            begin
              reg897 <= $unsigned((reg895 + $signed((~&(wire839 || wire885)))));
              reg898 <= (~&{({$unsigned(wire842), reg900[(2'h3):(2'h3)]} ?
                      wire840[(4'hb):(1'h0)] : $signed((reg895 ?
                          reg847 : reg893))),
                  (~^(^~{reg871}))});
              reg899 <= wire885[(4'hf):(4'hb)];
            end
          reg902 <= reg863[(2'h2):(2'h2)];
          reg903 <= reg898[(5'h10):(4'hf)];
        end
      else
        begin
          if ($unsigned($signed($signed({((8'had) - reg890)}))))
            begin
              reg895 <= ((~|$unsigned({$unsigned(wire842)})) ?
                  ($unsigned(reg866) ?
                      ((-$unsigned(reg880)) ?
                          $unsigned((reg875 >> reg869)) : ({reg903, (8'hac)} ?
                              ((7'h42) ? wire839 : reg892) : (wire860 ?
                                  reg855 : reg896))) : (-(8'haf))) : (~^(reg903 ?
                      reg872[(1'h1):(1'h1)] : {wire838})));
              reg896 <= reg856[(5'h12):(5'h11)];
              reg897 <= ($unsigned(wire839) ? reg901 : reg849[(4'hf):(4'hf)]);
              reg898 <= $signed(wire883[(2'h2):(1'h1)]);
            end
          else
            begin
              reg895 <= $unsigned(reg880[(4'h8):(3'h7)]);
              reg896 <= (reg861 ^ (~^reg857[(4'ha):(2'h2)]));
              reg897 <= ($unsigned(reg900[(3'h5):(3'h5)]) * ($unsigned(wire840[(3'h4):(2'h2)]) >= $signed((wire859[(3'h5):(1'h1)] ?
                  {reg902, reg850} : reg898[(4'hf):(3'h6)]))));
              reg898 <= (&$unsigned($signed({(^wire859),
                  reg847[(4'hb):(4'ha)]})));
            end
          reg899 <= ((reg898 != $unsigned({(reg881 ? reg858 : reg886),
              $unsigned(reg850)})) ~^ reg872);
          if ((^~(reg853 ?
              wire859[(3'h5):(2'h3)] : ($signed((^(8'hb0))) ^~ ($unsigned(reg850) & $signed(reg889))))))
            begin
              reg900 <= {(((reg897 ? $unsigned(reg868) : (reg866 * wire852)) ?
                          $unsigned({(8'ha9),
                              reg894}) : reg871[(3'h5):(3'h4)]) ?
                      {((wire884 >>> (8'hbd)) >>> wire859),
                          (wire841 ?
                              (~|wire852) : (reg847 ?
                                  reg878 : reg879))} : $unsigned((8'hb6)))};
              reg901 <= {({{{wire839, reg878}, (reg871 < reg890)}} ?
                      $unsigned($signed((&reg843))) : $signed(wire859[(1'h0):(1'h0)]))};
              reg902 <= $unsigned((reg873 ?
                  ({reg890[(2'h3):(2'h3)], (^reg900)} * ($unsigned(reg862) ?
                      reg880[(1'h0):(1'h0)] : ((7'h40) ?
                          wire839 : reg894))) : $unsigned($signed((reg903 ?
                      reg862 : reg850)))));
            end
          else
            begin
              reg900 <= ((wire839 >>> {($unsigned(reg875) - reg868),
                  ($signed(reg858) >> reg855)}) >> (~((reg843[(2'h3):(1'h1)] > (wire859 ?
                  reg853 : reg862)) >>> (reg895 ?
                  (!reg858) : reg890[(3'h4):(3'h4)]))));
              reg901 <= reg887[(4'h9):(2'h2)];
              reg902 <= (reg869 ~^ (~|(reg881 ?
                  ($unsigned((8'hab)) <= (reg855 ~^ reg900)) : ($signed(wire842) << {reg898}))));
              reg903 <= ($unsigned((($signed(reg847) ?
                      (~|reg902) : $signed(wire860)) <= (&$signed(reg853)))) ?
                  ($unsigned((8'hb1)) ?
                      (reg865[(4'hf):(4'he)] <<< ($unsigned(wire842) > (wire883 ?
                          reg897 : reg894))) : reg899) : (!reg880));
              reg904 <= reg871;
            end
          reg905 <= (-(reg900[(3'h7):(3'h7)] ~^ (reg864[(1'h0):(1'h0)] >= $signed((-reg899)))));
          if (wire839[(1'h0):(1'h0)])
            begin
              reg906 <= $signed($unsigned($signed($signed((reg897 != reg851)))));
            end
          else
            begin
              reg906 <= reg895[(3'h6):(2'h3)];
              reg907 <= $unsigned($signed(wire883));
              reg908 <= {wire841};
            end
        end
      reg909 <= reg849[(4'hc):(1'h1)];
    end
  always
    @(posedge clk) begin
      if (reg905)
        begin
          if ($unsigned(reg851))
            begin
              reg910 <= $unsigned((+(wire842 && {{wire884}, (~|reg892)})));
            end
          else
            begin
              reg910 <= {$unsigned($signed(($unsigned(reg910) ?
                      (reg900 ~^ wire842) : (reg857 >= (8'ha6))))),
                  $signed(((7'h40) != wire838))};
              reg911 <= $unsigned(wire883[(1'h0):(1'h0)]);
            end
          reg912 <= ($unsigned($unsigned($signed(reg894[(3'h6):(2'h3)]))) ?
              $signed($unsigned($unsigned($unsigned((8'ha3))))) : (8'hb6));
          reg913 <= $unsigned(($signed(((reg888 ^ (8'hb9)) ?
                  $signed(reg877) : $unsigned(reg854))) ?
              $signed((!reg861)) : {$unsigned((~&reg889)),
                  (reg899[(4'hb):(3'h4)] ^ reg894)}));
          reg914 <= $unsigned((^~{($unsigned(reg863) ?
                  (reg894 ? reg909 : reg905) : {reg854})}));
        end
      else
        begin
          if ($unsigned(($unsigned($unsigned((~^wire882))) + (($unsigned(reg857) * reg843[(3'h4):(3'h4)]) <<< (~|reg857)))))
            begin
              reg910 <= reg878[(4'hb):(1'h1)];
              reg911 <= $unsigned($unsigned({$unsigned((8'hb8)),
                  {$signed(reg875)}}));
              reg912 <= reg868;
              reg913 <= wire859[(2'h3):(2'h2)];
            end
          else
            begin
              reg910 <= (+((reg851 ?
                  (((8'h9c) ^ reg880) ?
                      reg893[(2'h2):(1'h1)] : (~&(8'hb6))) : $signed((+reg867))) >>> {$signed((reg897 ?
                      reg844 : reg893)),
                  $signed(reg866)}));
              reg911 <= $signed((8'ha0));
              reg912 <= reg874;
              reg913 <= $unsigned($unsigned(reg903));
              reg914 <= ({reg857[(2'h3):(1'h1)]} >= reg894[(2'h3):(2'h2)]);
            end
          reg915 <= (^(8'ha4));
          reg916 <= (+(8'hae));
          if (reg907)
            begin
              reg917 <= reg846[(4'h8):(3'h7)];
              reg918 <= (8'h9f);
            end
          else
            begin
              reg917 <= reg858;
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg867[(3'h7):(3'h4)])
        begin
          reg919 <= (&(reg851 ?
              reg867[(3'h7):(2'h2)] : $signed(($signed(wire884) | $unsigned(reg905)))));
          reg920 <= (~$unsigned({reg903}));
          reg921 <= ($unsigned((&$signed(reg917))) ?
              $unsigned(reg871) : $unsigned({(&(reg844 && reg847)),
                  reg890[(3'h7):(1'h0)]}));
          reg922 <= ((((8'ha4) - reg893[(3'h4):(3'h4)]) * $unsigned(wire884)) ?
              {reg845[(2'h2):(1'h0)]} : (+reg919));
          reg923 <= ($unsigned({(!(^~wire842))}) ?
              wire860 : (reg894 ^~ reg892[(2'h2):(1'h0)]));
        end
      else
        begin
          reg919 <= (reg919 == $unsigned($unsigned((~^(reg917 == wire883)))));
          reg920 <= $signed({(-$signed($signed(reg911)))});
          reg921 <= wire883[(1'h0):(1'h0)];
          reg922 <= ((^(8'hb3)) ?
              reg903 : $signed($unsigned((reg875 != (wire859 ?
                  reg892 : reg891)))));
          reg923 <= reg858[(4'h9):(1'h1)];
        end
      if ($unsigned(reg891))
        begin
          reg924 <= ((&(((reg892 << reg873) ? (reg913 >= reg846) : (8'ha1)) ?
              $signed($unsigned((8'h9c))) : (&{reg865,
                  reg910}))) >> $unsigned(reg844[(2'h2):(1'h0)]));
        end
      else
        begin
          if ((!(((reg912 ?
                  $unsigned((8'ha5)) : (reg917 & reg863)) + $unsigned({reg856})) ?
              (~^reg914[(1'h0):(1'h0)]) : (((reg878 <<< reg858) ?
                      $unsigned(reg871) : $signed(reg894)) ?
                  $signed($unsigned(reg861)) : reg903[(1'h0):(1'h0)]))))
            begin
              reg924 <= reg890[(5'h13):(4'h9)];
              reg925 <= ((reg917 <<< (reg900 >= reg848)) ^ $signed((reg866[(4'ha):(3'h4)] ?
                  $signed((~reg862)) : {reg850[(3'h5):(2'h2)]})));
              reg926 <= ((-(~&{$unsigned(reg866)})) ?
                  reg902 : ($unsigned({(^reg900),
                      reg905}) ^~ ($unsigned($unsigned(reg901)) * $signed(reg907[(3'h5):(1'h0)]))));
            end
          else
            begin
              reg924 <= (reg906 ^~ (8'hb7));
              reg925 <= reg891;
              reg926 <= wire882[(2'h3):(1'h1)];
            end
          reg927 <= (({(^~((8'ha7) ? (8'hbb) : reg893)),
                      {reg912[(1'h0):(1'h0)], reg904[(1'h1):(1'h0)]}} ?
                  ($signed((-reg880)) + reg913[(2'h3):(1'h1)]) : reg886[(2'h2):(2'h2)]) ?
              wire852 : (^(~^$unsigned(wire840[(4'h9):(2'h3)]))));
        end
      if (reg923[(4'hb):(2'h2)])
        begin
          if (($signed(($unsigned((wire882 ? wire883 : reg900)) ?
                  $unsigned((&(8'hb8))) : reg900)) ?
              reg857[(4'ha):(2'h3)] : $unsigned((8'hb5))))
            begin
              reg928 <= wire859;
              reg929 <= wire885;
              reg930 <= $unsigned($unsigned(reg925));
              reg931 <= {(((reg865 ?
                      {reg902,
                          reg929} : (!(8'ha4))) < reg917[(2'h2):(1'h0)]) > (!((reg928 ?
                      reg910 : reg898) < (reg911 ? reg927 : wire885))))};
            end
          else
            begin
              reg928 <= $unsigned(reg916);
              reg929 <= reg900;
              reg930 <= $signed(reg879[(3'h6):(3'h4)]);
              reg931 <= $unsigned((reg867 ^~ $unsigned(wire839)));
              reg932 <= reg843[(2'h3):(2'h2)];
            end
        end
      else
        begin
          if ((8'hb9))
            begin
              reg928 <= (|((reg870[(2'h2):(2'h2)] ?
                      reg919 : reg922[(2'h3):(2'h2)]) ?
                  reg909 : wire841));
              reg929 <= (($signed((&(reg856 ? reg897 : reg901))) ?
                  reg870[(1'h1):(1'h0)] : $signed((&reg857[(3'h5):(1'h0)]))) | (reg910[(3'h7):(2'h2)] ?
                  reg861 : $unsigned(reg915[(5'h10):(4'ha)])));
              reg930 <= reg903[(5'h13):(2'h2)];
            end
          else
            begin
              reg928 <= reg855[(2'h2):(1'h0)];
              reg929 <= $signed(($signed(reg846) >= (reg899[(3'h5):(1'h1)] ?
                  (wire840 ? (~|reg930) : (&reg868)) : ((reg906 ~^ reg870) ?
                      reg920[(1'h1):(1'h1)] : $unsigned(reg867)))));
              reg930 <= {(-{($signed(reg846) ^~ (reg928 ? (8'hb2) : (8'h9c))),
                      reg903})};
              reg931 <= (7'h44);
              reg932 <= reg849;
            end
        end
      reg933 <= reg858[(3'h4):(1'h1)];
      if ((reg918 * (($signed($unsigned(reg933)) > (+$unsigned(reg915))) ?
          $signed(((reg894 - reg851) == (reg915 >= reg897))) : (~(reg877 ?
              (|reg919) : (^reg906))))))
        begin
          reg934 <= reg901;
          reg935 <= reg926[(3'h4):(2'h2)];
          reg936 <= reg914[(2'h3):(1'h1)];
        end
      else
        begin
          if ((-$unsigned(reg918)))
            begin
              reg934 <= reg872[(3'h7):(3'h6)];
              reg935 <= (({((!reg865) ?
                          (reg916 < reg909) : {reg869, wire839})} ^ reg844) ?
                  (reg855 << (+((reg923 ? reg843 : reg914) ?
                      (wire840 && reg891) : $unsigned(reg868)))) : (reg935[(5'h12):(4'he)] ?
                      ($unsigned((reg845 ?
                          reg896 : reg899)) ~^ {(reg867 >> reg908)}) : reg897[(4'h9):(2'h2)]));
              reg936 <= $unsigned($unsigned(wire884[(5'h10):(4'h8)]));
            end
          else
            begin
              reg934 <= {$signed((~^($signed(reg862) <<< {reg892})))};
              reg935 <= (-(~&(($unsigned(reg894) ?
                  (reg932 ? reg902 : reg900) : ((8'had) ?
                      reg919 : reg931)) ^ reg878)));
              reg936 <= ($unsigned($unsigned($signed($signed((8'ha9))))) ~^ reg866[(4'hd):(4'hb)]);
              reg937 <= $unsigned((reg936 << $unsigned({$unsigned(reg927),
                  (reg928 ? reg911 : wire885)})));
            end
          if (reg898[(3'h6):(3'h4)])
            begin
              reg938 <= reg907[(3'h4):(1'h0)];
            end
          else
            begin
              reg938 <= reg873;
              reg939 <= reg923;
            end
          reg940 <= (reg923 ?
              reg871 : ((~reg922) >> $signed((^~reg893[(3'h5):(3'h5)]))));
          reg941 <= $unsigned((((^$signed(reg938)) <<< ({reg881,
                  reg889} & $signed(reg857))) ?
              $unsigned(reg894[(3'h4):(3'h4)]) : $signed(($signed(reg851) ?
                  reg856 : ((8'haa) > wire838)))));
          if (reg857)
            begin
              reg942 <= ({{($unsigned(reg922) ?
                              $signed((8'haa)) : (reg925 - reg919)),
                          reg915},
                      $unsigned(reg931)} ?
                  (((!$unsigned(reg866)) ~^ (~$signed(reg899))) ?
                      $unsigned($unsigned(reg935)) : $signed($unsigned($unsigned(reg871)))) : $signed({$signed($signed(reg875))}));
            end
          else
            begin
              reg942 <= ((~|($signed((~^reg927)) ?
                  reg850 : (|(reg920 >= reg899)))) && (7'h40));
              reg943 <= (reg893 ?
                  (~^reg874[(2'h2):(1'h0)]) : reg866[(3'h5):(2'h3)]);
              reg944 <= reg935[(3'h5):(1'h0)];
              reg945 <= reg867[(5'h10):(4'ha)];
            end
        end
    end
  assign wire946 = reg918[(4'he):(4'ha)];
  assign wire947 = (({reg942} >> $unsigned(reg876[(3'h6):(3'h6)])) ?
                       $signed((($signed(reg924) > $unsigned((8'ha5))) ^~ (8'hb2))) : (&(((wire882 ?
                           reg877 : reg888) - $unsigned(reg916)) <= {reg876})));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1091  (y, clk, wire1096, wire1095, wire1094, wire1093, wire1092);
  output wire [(32'h3e5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire1096;
  input wire signed [(4'he):(1'h0)] wire1095;
  input wire signed [(3'h4):(1'h0)] wire1094;
  input wire signed [(5'h15):(1'h0)] wire1093;
  input wire signed [(4'hf):(1'h0)] wire1092;
  wire [(4'he):(1'h0)] wire1184;
  wire [(5'h10):(1'h0)] wire1183;
  reg [(4'ha):(1'h0)] reg1182 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1181 = (1'h0);
  reg [(3'h4):(1'h0)] reg1180 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1179 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1178 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1177 = (1'h0);
  reg [(4'he):(1'h0)] reg1176 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1175 = (1'h0);
  reg [(2'h3):(1'h0)] reg1174 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1173 = (1'h0);
  reg [(5'h10):(1'h0)] reg1172 = (1'h0);
  reg [(5'h11):(1'h0)] reg1171 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1170 = (1'h0);
  reg [(3'h5):(1'h0)] reg1169 = (1'h0);
  reg [(5'h15):(1'h0)] reg1168 = (1'h0);
  reg [(4'hf):(1'h0)] reg1167 = (1'h0);
  reg [(3'h4):(1'h0)] reg1166 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1165 = (1'h0);
  reg [(5'h15):(1'h0)] reg1164 = (1'h0);
  reg [(4'h9):(1'h0)] reg1163 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1162 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1161 = (1'h0);
  reg [(4'ha):(1'h0)] reg1160 = (1'h0);
  reg [(4'h8):(1'h0)] reg1159 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1158 = (1'h0);
  reg [(2'h2):(1'h0)] reg1157 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1156 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1155 = (1'h0);
  reg [(4'he):(1'h0)] reg1154 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1153 = (1'h0);
  reg [(4'h8):(1'h0)] reg1152 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1151 = (1'h0);
  reg [(5'h13):(1'h0)] reg1150 = (1'h0);
  reg [(2'h2):(1'h0)] reg1149 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1148 = (1'h0);
  reg [(4'hd):(1'h0)] reg1147 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1146 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1145 = (1'h0);
  reg [(5'h12):(1'h0)] reg1144 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1143 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1142 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1141 = (1'h0);
  reg [(4'hd):(1'h0)] reg1140 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1139 = (1'h0);
  wire [(4'ha):(1'h0)] wire1138;
  wire [(5'h13):(1'h0)] wire1137;
  wire signed [(3'h4):(1'h0)] wire1136;
  reg signed [(5'h10):(1'h0)] reg1135 = (1'h0);
  reg [(5'h13):(1'h0)] reg1134 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1133 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1132 = (1'h0);
  reg [(5'h14):(1'h0)] reg1131 = (1'h0);
  reg [(4'hf):(1'h0)] reg1130 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1129 = (1'h0);
  reg [(4'h8):(1'h0)] reg1128 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1127 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1126 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1125 = (1'h0);
  reg [(3'h5):(1'h0)] reg1124 = (1'h0);
  reg [(4'hb):(1'h0)] reg1123 = (1'h0);
  reg [(4'h8):(1'h0)] reg1122 = (1'h0);
  reg [(5'h11):(1'h0)] reg1121 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1120 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1119 = (1'h0);
  reg [(5'h13):(1'h0)] reg1118 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire1117;
  wire [(5'h11):(1'h0)] wire1116;
  wire [(2'h2):(1'h0)] wire1115;
  wire signed [(3'h4):(1'h0)] wire1114;
  reg [(4'hb):(1'h0)] reg1113 = (1'h0);
  reg [(5'h13):(1'h0)] reg1112 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1111 = (1'h0);
  reg [(5'h12):(1'h0)] reg1110 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1109 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1108 = (1'h0);
  reg [(5'h13):(1'h0)] reg1107 = (1'h0);
  reg [(4'h8):(1'h0)] reg1106 = (1'h0);
  reg [(4'hf):(1'h0)] reg1105 = (1'h0);
  reg [(3'h4):(1'h0)] reg1104 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1103 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1102 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1101 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1100 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1099 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1098 = (1'h0);
  wire [(2'h2):(1'h0)] wire1097;
  assign y = {wire1184,
                 wire1183,
                 reg1182,
                 reg1181,
                 reg1180,
                 reg1179,
                 reg1178,
                 reg1177,
                 reg1176,
                 reg1175,
                 reg1174,
                 reg1173,
                 reg1172,
                 reg1171,
                 reg1170,
                 reg1169,
                 reg1168,
                 reg1167,
                 reg1166,
                 reg1165,
                 reg1164,
                 reg1163,
                 reg1162,
                 reg1161,
                 reg1160,
                 reg1159,
                 reg1158,
                 reg1157,
                 reg1156,
                 reg1155,
                 reg1154,
                 reg1153,
                 reg1152,
                 reg1151,
                 reg1150,
                 reg1149,
                 reg1148,
                 reg1147,
                 reg1146,
                 reg1145,
                 reg1144,
                 reg1143,
                 reg1142,
                 reg1141,
                 reg1140,
                 reg1139,
                 wire1138,
                 wire1137,
                 wire1136,
                 reg1135,
                 reg1134,
                 reg1133,
                 reg1132,
                 reg1131,
                 reg1130,
                 reg1129,
                 reg1128,
                 reg1127,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1123,
                 reg1122,
                 reg1121,
                 reg1120,
                 reg1119,
                 reg1118,
                 wire1117,
                 wire1116,
                 wire1115,
                 wire1114,
                 reg1113,
                 reg1112,
                 reg1111,
                 reg1110,
                 reg1109,
                 reg1108,
                 reg1107,
                 reg1106,
                 reg1105,
                 reg1104,
                 reg1103,
                 reg1102,
                 reg1101,
                 reg1100,
                 reg1099,
                 reg1098,
                 wire1097,
                 (1'h0)};
  assign wire1097 = $signed({(|wire1093),
                        $signed(((~|wire1095) - $unsigned((8'hbd))))});
  always
    @(posedge clk) begin
      reg1098 <= {wire1097[(1'h1):(1'h0)]};
      reg1099 <= wire1092;
      reg1100 <= wire1095;
      if ({{wire1094, ((+(^wire1095)) > reg1099)}})
        begin
          reg1101 <= wire1095;
          reg1102 <= $signed((8'ha9));
          reg1103 <= wire1096[(3'h7):(3'h5)];
          if ((reg1099[(4'ha):(3'h7)] < wire1093))
            begin
              reg1104 <= $signed(reg1101);
            end
          else
            begin
              reg1104 <= (|$signed((&wire1097)));
              reg1105 <= $signed(reg1098[(2'h3):(1'h1)]);
            end
          if (reg1105[(3'h6):(3'h4)])
            begin
              reg1106 <= (reg1101 ?
                  reg1098 : (reg1103 ?
                      ($signed($signed((8'hb4))) ?
                          (reg1104 <= $signed(wire1092)) : {{wire1096}}) : {{$signed((8'ha5)),
                              reg1105[(4'he):(4'hc)]},
                          (wire1093 >= (^reg1098))}));
              reg1107 <= {$signed($signed(reg1099)),
                  $signed((reg1098 == (+wire1092[(1'h1):(1'h0)])))};
            end
          else
            begin
              reg1106 <= $unsigned($unsigned($signed(wire1093[(5'h11):(4'hd)])));
            end
        end
      else
        begin
          if (wire1096)
            begin
              reg1101 <= $signed(($unsigned(reg1102[(1'h1):(1'h0)]) || reg1103[(3'h6):(1'h1)]));
            end
          else
            begin
              reg1101 <= $unsigned($unsigned(((~|wire1092) ^ reg1104)));
              reg1102 <= (~&((($unsigned(reg1106) ?
                      (reg1102 ? (8'h9f) : (8'h9c)) : wire1092) ?
                  {$unsigned(wire1096)} : ((reg1099 ?
                      reg1100 : reg1099) ^~ ((8'hb0) || reg1101))) ~^ ((((8'hb1) >>> wire1096) ?
                  (!reg1106) : reg1105[(1'h0):(1'h0)]) != ((reg1107 ?
                      reg1098 : reg1099) ?
                  wire1096 : $unsigned(reg1105)))));
              reg1103 <= reg1101;
              reg1104 <= $unsigned(wire1092);
              reg1105 <= ((~^$unsigned((~^(wire1092 ?
                  (7'h43) : reg1100)))) >> reg1103[(1'h0):(1'h0)]);
            end
          reg1106 <= $signed((&(-$signed($signed(reg1101)))));
          if ((((reg1101[(2'h3):(1'h0)] ?
                  (^(-reg1102)) : wire1094[(2'h2):(1'h0)]) ?
              $signed((8'h9e)) : (reg1103 ?
                  ((wire1093 ?
                      reg1103 : wire1092) < $signed(wire1093)) : (^~reg1101))) + $signed((~&(+(wire1097 ?
              reg1103 : reg1102))))))
            begin
              reg1107 <= (^~((~{((8'ha2) >> (8'h9e))}) + (~$unsigned((reg1103 ?
                  wire1097 : wire1093)))));
              reg1108 <= {wire1097[(1'h1):(1'h0)]};
              reg1109 <= (~|($unsigned((wire1094[(2'h3):(1'h1)] || (^wire1095))) && ($signed(reg1101[(2'h3):(1'h1)]) ?
                  reg1104[(1'h1):(1'h0)] : {(wire1097 || reg1104)})));
              reg1110 <= $signed($signed(wire1092[(3'h7):(1'h0)]));
            end
          else
            begin
              reg1107 <= (&((((reg1101 ? reg1098 : reg1103) ?
                          (reg1104 ? reg1108 : wire1095) : (~^reg1110)) ?
                      $unsigned(reg1102) : wire1095) ?
                  $unsigned({(reg1106 || (8'had))}) : $signed(((8'hb5) ?
                      (wire1094 ? reg1108 : reg1110) : (~&wire1097)))));
              reg1108 <= $unsigned(reg1103[(4'hc):(4'h8)]);
            end
          reg1111 <= (^~$signed(wire1095[(2'h2):(2'h2)]));
          reg1112 <= reg1102[(3'h5):(1'h1)];
        end
      reg1113 <= reg1111;
    end
  assign wire1114 = (|reg1101);
  assign wire1115 = reg1106[(3'h5):(1'h1)];
  assign wire1116 = (&((|((reg1108 ? reg1104 : reg1109) < (reg1112 ?
                        (8'ha4) : wire1115))) >= ($unsigned((^(8'hb7))) ?
                        $unsigned((reg1102 ?
                            reg1105 : wire1096)) : (reg1109[(1'h1):(1'h1)] ~^ (+reg1107)))));
  assign wire1117 = (~^(!(^reg1105[(3'h5):(1'h1)])));
  always
    @(posedge clk) begin
      if (reg1099[(1'h0):(1'h0)])
        begin
          reg1118 <= ($signed(reg1103[(4'ha):(3'h6)]) ?
              $unsigned(wire1116[(4'hd):(3'h4)]) : ($unsigned((~|$unsigned(reg1099))) - $signed(wire1117)));
          reg1119 <= (7'h42);
        end
      else
        begin
          reg1118 <= (reg1101[(3'h4):(3'h4)] ?
              {$unsigned(((~|reg1112) ?
                      (wire1115 ?
                          (8'hb0) : reg1098) : (reg1106 & reg1106)))} : (7'h40));
          if ((reg1105 + ($unsigned(reg1100) ?
              reg1100[(3'h4):(3'h4)] : {{$unsigned(reg1100), $signed((7'h40))},
                  wire1096})))
            begin
              reg1119 <= ($unsigned((~reg1108)) >> reg1098[(3'h6):(1'h1)]);
            end
          else
            begin
              reg1119 <= ($signed((&$unsigned((reg1112 < wire1114)))) ?
                  (-reg1112[(4'ha):(3'h6)]) : {{reg1107[(1'h0):(1'h0)]},
                      ((~wire1115[(2'h2):(1'h1)]) * ($unsigned(wire1096) ?
                          $signed(reg1101) : $signed(wire1096)))});
              reg1120 <= (($signed({(~|wire1116)}) <= wire1096) ?
                  (({wire1117[(3'h7):(3'h6)]} && {$unsigned((8'h9d)),
                      reg1119[(4'hb):(4'h8)]}) | $signed($signed((reg1108 ?
                      wire1116 : (8'hb7))))) : (wire1117[(3'h6):(3'h4)] ?
                      $signed($signed($unsigned(reg1112))) : (&reg1098)));
              reg1121 <= (!reg1113);
              reg1122 <= $signed($signed($unsigned($signed(reg1099))));
              reg1123 <= $signed(reg1113);
            end
          reg1124 <= (($unsigned(($signed(reg1119) ?
                  {reg1118} : $signed(reg1112))) << $signed(reg1120[(1'h1):(1'h0)])) ?
              (((~|$unsigned((8'hb2))) ^ $signed(((8'hb1) ?
                  wire1094 : wire1117))) & ((~^(reg1111 || reg1112)) ^~ reg1100[(2'h2):(2'h2)])) : (8'hba));
        end
      reg1125 <= reg1124[(1'h0):(1'h0)];
      reg1126 <= reg1102[(2'h3):(2'h3)];
      if ($signed($signed({reg1108,
          (wire1117[(4'he):(3'h4)] ?
              $unsigned(reg1102) : (reg1103 ~^ (8'ha8)))})))
        begin
          if ((($unsigned(((-reg1123) & reg1104[(1'h0):(1'h0)])) & $signed((8'hb6))) >= ($signed({$signed(reg1123)}) < reg1100[(3'h5):(3'h5)])))
            begin
              reg1127 <= $unsigned(reg1124[(1'h1):(1'h1)]);
            end
          else
            begin
              reg1127 <= (!$unsigned(((-(reg1104 != reg1109)) > ((~&wire1093) - reg1103[(2'h3):(2'h2)]))));
              reg1128 <= wire1116;
              reg1129 <= {(reg1119[(3'h5):(1'h0)] ?
                      (-$signed((&reg1099))) : ($unsigned(((8'hb1) ^~ reg1102)) & wire1116[(4'ha):(4'h8)])),
                  (~&reg1103)};
              reg1130 <= ((wire1117 >>> $signed((reg1108 ?
                      reg1103 : wire1095))) ?
                  $signed($signed(wire1097)) : (wire1117 >= (~|((reg1104 < reg1129) ?
                      reg1107[(1'h0):(1'h0)] : (reg1107 == reg1108)))));
              reg1131 <= wire1117;
            end
          reg1132 <= ((~((reg1128 ? (-(8'haf)) : (~reg1101)) ?
              reg1112 : (&$unsigned(reg1125)))) & $signed({(^$unsigned(reg1098))}));
          reg1133 <= reg1131;
          reg1134 <= (!$signed(reg1113));
        end
      else
        begin
          reg1127 <= (reg1102 != $unsigned($unsigned($unsigned({reg1101,
              reg1132}))));
          reg1128 <= $signed({(reg1103[(4'ha):(2'h2)] ~^ (+wire1096)),
              {(~$signed(reg1113))}});
          if ($unsigned(reg1128[(3'h4):(2'h2)]))
            begin
              reg1129 <= reg1105;
              reg1130 <= reg1123;
            end
          else
            begin
              reg1129 <= (!$signed(wire1097[(1'h1):(1'h0)]));
              reg1130 <= $signed($unsigned((({wire1115} ^~ (wire1092 <= reg1111)) | {$unsigned(reg1100)})));
              reg1131 <= {$signed($signed(((wire1096 ?
                      reg1107 : wire1117) | $unsigned(reg1128))))};
            end
          reg1132 <= {reg1100[(4'h9):(1'h1)],
              (((+reg1134) >= ($signed(reg1098) >= reg1131[(3'h6):(3'h5)])) | $unsigned({reg1124[(1'h0):(1'h0)]}))};
        end
      reg1135 <= $unsigned($unsigned((({wire1116, wire1117} ?
              reg1106[(2'h3):(2'h2)] : (reg1100 >> reg1113)) ?
          (&wire1117[(3'h7):(2'h2)]) : ($unsigned(reg1113) ?
              {reg1104, reg1110} : (8'hab)))));
    end
  assign wire1136 = reg1103[(4'hc):(3'h7)];
  assign wire1137 = ((((+{(8'ha0)}) ?
                                ((reg1124 > reg1106) == $unsigned(reg1125)) : reg1122[(4'h8):(3'h6)]) ?
                            $unsigned(reg1108) : (^$signed((~(7'h43))))) ?
                        ((~$signed(reg1098[(3'h5):(3'h4)])) > ($unsigned(reg1120[(2'h2):(1'h0)]) ?
                            $signed((reg1104 ?
                                reg1129 : reg1108)) : $signed((wire1136 ?
                                reg1118 : (7'h41))))) : {(({reg1129,
                                    wire1095} && ((8'ha6) ?
                                    reg1110 : reg1135)) ?
                                $signed(wire1117[(1'h0):(1'h0)]) : wire1116[(2'h3):(2'h2)])});
  assign wire1138 = ($unsigned((&{(~wire1117)})) ?
                        (wire1115[(2'h2):(1'h0)] << (reg1118 ?
                            (-(!reg1128)) : (~|{(8'h9d)}))) : reg1112);
  always
    @(posedge clk) begin
      if (((reg1134[(1'h1):(1'h0)] ?
              (reg1106 ?
                  reg1112[(4'hf):(4'hd)] : (~^(reg1098 ?
                      wire1096 : (8'hae)))) : $unsigned($unsigned((!wire1138)))) ?
          (^~(($signed(wire1115) >= {reg1102, wire1136}) ?
              ((reg1113 != reg1105) ?
                  (reg1098 ~^ reg1105) : $signed((8'hab))) : $unsigned($signed(reg1104)))) : $signed(reg1109[(1'h0):(1'h0)])))
        begin
          if (((^~$signed($unsigned($unsigned(reg1125)))) < $unsigned($signed($unsigned($unsigned(wire1097))))))
            begin
              reg1139 <= (&wire1095[(2'h3):(2'h3)]);
              reg1140 <= reg1112[(5'h10):(4'he)];
              reg1141 <= (+(+(^$signed((reg1133 ? reg1119 : (8'ha5))))));
            end
          else
            begin
              reg1139 <= ($unsigned({(+$signed(reg1099)),
                  $unsigned({wire1137, reg1130})}) & (-($unsigned(wire1114) ?
                  ((~^wire1092) ?
                      (reg1109 ?
                          reg1107 : (8'h9e)) : reg1132) : (reg1141[(4'h9):(3'h4)] ?
                      (reg1112 >>> wire1114) : reg1102[(1'h0):(1'h0)]))));
              reg1140 <= (^~$signed({$signed($unsigned(reg1103))}));
              reg1141 <= reg1139[(4'hc):(4'hb)];
              reg1142 <= {reg1131[(5'h10):(5'h10)], reg1106};
              reg1143 <= $unsigned((~|reg1123[(3'h5):(3'h4)]));
            end
          if (reg1140[(4'ha):(2'h3)])
            begin
              reg1144 <= ((^~reg1119[(3'h4):(2'h2)]) ?
                  $signed($unsigned(wire1116)) : (reg1140 ? reg1107 : reg1100));
              reg1145 <= (($signed(reg1110) ?
                  $signed((wire1096[(1'h1):(1'h1)] < $signed((8'hb7)))) : reg1141[(1'h1):(1'h1)]) ~^ $signed(((reg1144 ?
                      reg1108 : (reg1125 && (8'hb9))) ?
                  (wire1117 ?
                      wire1137[(1'h1):(1'h1)] : $signed(reg1143)) : ($signed(reg1121) ?
                      $unsigned(reg1125) : reg1098[(2'h3):(1'h1)]))));
              reg1146 <= reg1127;
              reg1147 <= $signed((reg1111 ? reg1128[(3'h4):(2'h3)] : reg1107));
            end
          else
            begin
              reg1144 <= wire1117;
            end
        end
      else
        begin
          reg1139 <= reg1109;
          reg1140 <= (~$signed(reg1105));
          reg1141 <= $signed(reg1127[(2'h2):(2'h2)]);
          reg1142 <= reg1134;
        end
      if ((~|$signed($unsigned(({(7'h43)} & $unsigned(reg1112))))))
        begin
          reg1148 <= $signed((~^reg1118));
          reg1149 <= (^((8'hb8) ?
              {({reg1121,
                      wire1116} || reg1130)} : $unsigned($unsigned((reg1099 <= wire1117)))));
          reg1150 <= ($unsigned((((reg1130 | reg1132) ?
                  reg1133[(2'h2):(1'h1)] : reg1128) >> ((-(8'hb0)) ?
                  $unsigned(reg1139) : {reg1098, (8'hb5)}))) ?
              ($unsigned(reg1113[(4'ha):(3'h5)]) && (reg1144 >> ($signed((8'h9d)) ~^ (!reg1142)))) : (^$unsigned(((reg1104 > reg1149) != (~|wire1138)))));
          if ((^~{$unsigned(((reg1146 ^~ reg1149) + {reg1106})),
              $signed((reg1118[(1'h1):(1'h1)] || {reg1121, reg1129}))}))
            begin
              reg1151 <= ({$unsigned((-{reg1105, reg1105})),
                  {(^~reg1145[(4'h9):(2'h2)])}} == $signed($unsigned(((8'hb8) > (reg1103 ?
                  reg1143 : reg1102)))));
              reg1152 <= wire1096;
              reg1153 <= (~wire1092);
              reg1154 <= ((~&reg1108) ?
                  {reg1134[(1'h1):(1'h0)]} : $unsigned(reg1135[(3'h4):(2'h3)]));
              reg1155 <= $signed($unsigned(reg1106[(1'h1):(1'h1)]));
            end
          else
            begin
              reg1151 <= {(~|wire1092[(4'h9):(4'h8)]),
                  $unsigned((!($unsigned((8'ha8)) >> (reg1100 ?
                      wire1097 : (8'hb6)))))};
              reg1152 <= (wire1115 ?
                  (7'h41) : {$signed(((^reg1104) ?
                          ((8'ha3) + reg1147) : $unsigned(reg1151)))});
              reg1153 <= reg1120;
              reg1154 <= wire1097[(1'h0):(1'h0)];
              reg1155 <= wire1117[(4'hf):(3'h6)];
            end
        end
      else
        begin
          reg1148 <= reg1150[(4'he):(2'h3)];
          reg1149 <= $unsigned(reg1141[(1'h0):(1'h0)]);
        end
      if (((+$signed($signed($unsigned(reg1124)))) != (+$signed($unsigned((~&reg1100))))))
        begin
          if ((($unsigned((reg1111[(1'h1):(1'h0)] * {(7'h42)})) >= $signed(({reg1155} ?
              (wire1136 ?
                  (8'haf) : reg1143) : $unsigned(reg1126)))) + $signed({reg1113})))
            begin
              reg1156 <= (^~({{(reg1140 ? wire1092 : (8'hb4)),
                          (wire1115 | reg1106)},
                      reg1121[(4'h9):(3'h7)]} ?
                  reg1149[(1'h0):(1'h0)] : reg1119));
              reg1157 <= $signed(wire1114[(1'h1):(1'h0)]);
              reg1158 <= reg1141;
            end
          else
            begin
              reg1156 <= $unsigned((8'ha5));
              reg1157 <= $unsigned((($signed(reg1123) ?
                  $signed((&reg1100)) : ({(8'h9f)} > (reg1149 ?
                      reg1147 : reg1158))) >= reg1155));
              reg1158 <= reg1123;
              reg1159 <= wire1114;
            end
          reg1160 <= (reg1100[(4'h9):(3'h4)] ?
              $unsigned(reg1146[(1'h1):(1'h1)]) : reg1159[(3'h4):(1'h1)]);
        end
      else
        begin
          if ((($signed(reg1142[(2'h2):(1'h1)]) ?
                  ({$signed((8'hae)), ((8'hb3) ? wire1114 : reg1157)} ?
                      $signed($signed(reg1143)) : (reg1148[(3'h6):(3'h6)] && $signed((8'hac)))) : reg1107[(3'h4):(1'h0)]) ?
              reg1160 : ($unsigned(($unsigned(reg1155) << (^~reg1153))) | (!$unsigned({wire1137,
                  reg1146})))))
            begin
              reg1156 <= reg1154[(4'hb):(3'h7)];
              reg1157 <= {($unsigned({((7'h40) ? wire1095 : reg1155),
                      reg1120}) >= {(~&{reg1106, reg1125}),
                      {(+reg1107), (reg1118 ? wire1115 : (7'h43))}}),
                  reg1103[(2'h2):(1'h0)]};
              reg1158 <= ($signed(reg1139) ?
                  $unsigned(wire1094[(3'h4):(2'h3)]) : $unsigned(((~|$signed(wire1095)) < (reg1131[(4'ha):(3'h6)] ?
                      (reg1101 ? reg1152 : reg1108) : (~^reg1133)))));
            end
          else
            begin
              reg1156 <= wire1115[(1'h0):(1'h0)];
              reg1157 <= reg1122[(4'h8):(1'h0)];
            end
          reg1159 <= (^(~|reg1154[(1'h1):(1'h0)]));
          reg1160 <= (($signed(($signed(reg1113) ?
                      reg1102[(1'h1):(1'h1)] : reg1126[(3'h4):(1'h0)])) ?
                  ($unsigned((reg1140 <= reg1129)) ?
                      $unsigned((reg1152 != (8'hb5))) : reg1152[(4'h8):(2'h2)]) : ($unsigned(((8'had) ?
                      reg1123 : (7'h42))) ^ ((^(8'h9f)) | (reg1112 >> reg1130)))) ?
              wire1114 : reg1110[(5'h11):(2'h2)]);
          reg1161 <= ($signed($unsigned($unsigned(reg1102[(3'h5):(2'h2)]))) | (wire1114 ?
              $signed(((reg1100 ? wire1114 : wire1093) ?
                  (^~reg1132) : (reg1098 ? wire1094 : reg1124))) : wire1095));
        end
      if (reg1099)
        begin
          reg1162 <= $signed(({reg1144[(4'hb):(3'h5)]} ?
              reg1099 : $signed($signed(((8'hab) ? wire1093 : (8'ha4))))));
        end
      else
        begin
          if ($signed($signed((reg1155 << reg1150[(4'h8):(3'h4)]))))
            begin
              reg1162 <= (({reg1156[(2'h3):(1'h1)]} ?
                      (~&reg1141) : reg1143[(1'h0):(1'h0)]) ?
                  ($unsigned($unsigned((reg1129 ? reg1150 : reg1122))) ?
                      $signed(reg1113[(4'hb):(1'h0)]) : $unsigned((+(reg1151 ^~ reg1130)))) : (($signed($unsigned(reg1133)) - (&reg1133[(3'h5):(2'h2)])) ?
                      $signed($signed($signed(reg1144))) : $signed((reg1102[(2'h3):(2'h3)] < (reg1102 ?
                          (8'hbd) : reg1121)))));
              reg1163 <= {(-(+(8'hbc)))};
              reg1164 <= $unsigned(((reg1118[(1'h1):(1'h1)] ?
                  ({wire1136} ?
                      $unsigned(reg1102) : ((8'hbb) | reg1144)) : {wire1136[(2'h2):(1'h1)],
                      $signed((7'h41))}) < (((wire1095 ? reg1134 : reg1151) ?
                  (reg1153 ?
                      reg1130 : reg1159) : $unsigned(reg1123)) << ((8'hbb) ?
                  (~^reg1100) : (8'hb6)))));
            end
          else
            begin
              reg1162 <= $signed(reg1154);
              reg1163 <= reg1144;
              reg1164 <= reg1129;
              reg1165 <= (reg1143[(1'h1):(1'h0)] ?
                  $signed((|reg1139)) : ((-reg1146[(1'h0):(1'h0)]) ?
                      $signed(((reg1122 <= reg1129) >>> (reg1164 + wire1096))) : (reg1105 << (reg1111[(3'h5):(2'h3)] <= $unsigned(reg1141)))));
            end
          if ($unsigned($unsigned($signed(reg1145))))
            begin
              reg1166 <= reg1106[(1'h0):(1'h0)];
              reg1167 <= (reg1145[(2'h3):(2'h3)] * $signed(reg1102[(2'h2):(1'h1)]));
              reg1168 <= reg1135[(4'h9):(1'h0)];
              reg1169 <= (8'ha6);
              reg1170 <= ($signed($unsigned($unsigned(reg1118[(5'h10):(3'h5)]))) >= (reg1169[(3'h5):(3'h5)] ?
                  ((~^(wire1097 ?
                      reg1165 : reg1163)) || reg1104) : wire1093[(5'h12):(1'h1)]));
            end
          else
            begin
              reg1166 <= $unsigned((~|$signed(reg1118)));
              reg1167 <= reg1149[(2'h2):(1'h1)];
            end
          reg1171 <= $signed((~&{$unsigned((reg1143 ? reg1112 : reg1101)),
              ($unsigned(reg1125) ? wire1117 : $unsigned(reg1103))}));
        end
      if ((&reg1135[(4'hf):(4'ha)]))
        begin
          reg1172 <= (reg1124 ~^ wire1136[(3'h4):(3'h4)]);
          reg1173 <= (~^wire1117);
          reg1174 <= ($signed(wire1092) || reg1122[(3'h4):(3'h4)]);
        end
      else
        begin
          reg1172 <= $signed($signed((~|(~&$signed(reg1110)))));
          reg1173 <= ($signed(((&(reg1170 ^ reg1140)) ?
              $signed((8'hac)) : (^~{(8'had),
                  reg1143}))) != $unsigned((-($unsigned(reg1163) ?
              $unsigned((8'hb7)) : reg1161))));
          reg1174 <= $signed(reg1103);
          if (reg1119[(4'hc):(4'hc)])
            begin
              reg1175 <= (|$unsigned($signed(($unsigned(reg1133) >>> (reg1159 >> reg1122)))));
            end
          else
            begin
              reg1175 <= reg1123[(4'h9):(3'h5)];
              reg1176 <= ($signed($signed(({(8'ha6), reg1164} ?
                  ((8'haf) ^ reg1150) : $unsigned(reg1118)))) & $signed((!((reg1105 > reg1147) <= (reg1140 >> reg1122)))));
              reg1177 <= $signed($unsigned(($signed((reg1153 ?
                  reg1169 : reg1139)) != ((reg1172 == reg1128) ?
                  (!reg1143) : $signed(reg1173)))));
              reg1178 <= reg1109[(1'h1):(1'h1)];
              reg1179 <= $signed($signed(reg1176[(3'h7):(3'h4)]));
            end
          if ($unsigned(reg1157))
            begin
              reg1180 <= $unsigned((-reg1123));
              reg1181 <= ($signed(($signed($unsigned(wire1096)) ?
                      ((reg1148 ? reg1161 : reg1107) ?
                          {wire1116,
                              reg1149} : $unsigned((8'hb5))) : reg1180[(2'h3):(2'h2)])) ?
                  $signed({((reg1151 ? (8'hab) : reg1171) * (wire1092 ?
                          reg1154 : reg1173))}) : ((^(~{reg1156,
                      reg1101})) >= reg1159[(2'h3):(1'h1)]));
              reg1182 <= $unsigned((~^(($signed((8'hb4)) || $unsigned(reg1172)) & $unsigned((|reg1148)))));
            end
          else
            begin
              reg1180 <= reg1145;
              reg1181 <= $signed((($signed({reg1130}) ?
                      (((8'ha4) <<< wire1136) && reg1139) : wire1094[(1'h1):(1'h1)]) ?
                  (~^(^(reg1168 ^~ reg1160))) : {({reg1175,
                          reg1163} <= $unsigned(reg1149)),
                      wire1136}));
            end
        end
    end
  assign wire1183 = $signed((reg1124[(3'h4):(1'h1)] ?
                        $unsigned($signed((reg1108 ?
                            wire1116 : wire1096))) : (reg1144[(4'he):(3'h4)] ?
                            (~|$signed((8'ha3))) : (((8'ha6) + reg1168) ?
                                reg1124 : (8'hbd)))));
  assign wire1184 = $signed(((reg1111 ?
                        $signed((-(7'h40))) : ($unsigned(wire1093) ~^ (reg1100 ?
                            reg1144 : (8'hb8)))) >> reg1143[(4'h9):(2'h3)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1299
#( parameter param1322 = {((((+(8'hb1)) >>> ((8'hab) > (8'ha9))) + (-(7'h43))) ? (+(((8'hbb) ? (8'ha2) : (8'ha5)) ? {(8'hb6), (8'h9f)} : (~|(8'hbd)))) : ((((8'hb1) ? (8'hb9) : (8'h9e)) ? ((7'h43) < (8'hbd)) : (-(8'ha5))) ? (((8'hb1) < (8'ha7)) * ((8'hb8) < (8'hb4))) : {((7'h43) ^~ (8'hae)), ((8'haf) ? (8'hab) : (8'hb1))})), (-(({(7'h44)} && {(8'hb1), (8'ha6)}) ? {((8'ha2) ? (8'hb7) : (8'ha8)), (~&(7'h43))} : ((!(8'h9f)) || (8'hb1))))}
, parameter param1323 = (|((!(^(param1322 == param1322))) ? param1322 : (((8'hb0) ? (^param1322) : (~&param1322)) < param1322))) )
(y, clk, wire1304, wire1303, wire1302, wire1301, wire1300);
  output wire [(32'hca):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire1304;
  input wire signed [(5'h15):(1'h0)] wire1303;
  input wire signed [(5'h15):(1'h0)] wire1302;
  input wire signed [(4'ha):(1'h0)] wire1301;
  input wire signed [(4'h8):(1'h0)] wire1300;
  wire signed [(5'h11):(1'h0)] wire1321;
  reg signed [(4'hc):(1'h0)] reg1320 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1319 = (1'h0);
  wire [(4'h8):(1'h0)] wire1318;
  wire signed [(4'he):(1'h0)] wire1317;
  wire signed [(3'h7):(1'h0)] wire1316;
  wire signed [(4'h8):(1'h0)] wire1315;
  wire signed [(5'h15):(1'h0)] wire1314;
  wire signed [(3'h4):(1'h0)] wire1313;
  wire [(4'he):(1'h0)] wire1312;
  wire signed [(3'h4):(1'h0)] wire1311;
  wire signed [(2'h3):(1'h0)] wire1310;
  wire signed [(5'h11):(1'h0)] wire1309;
  wire [(5'h14):(1'h0)] wire1308;
  wire signed [(4'he):(1'h0)] wire1307;
  wire signed [(4'h9):(1'h0)] wire1306;
  wire signed [(4'hf):(1'h0)] wire1305;
  assign y = {wire1321,
                 reg1320,
                 reg1319,
                 wire1318,
                 wire1317,
                 wire1316,
                 wire1315,
                 wire1314,
                 wire1313,
                 wire1312,
                 wire1311,
                 wire1310,
                 wire1309,
                 wire1308,
                 wire1307,
                 wire1306,
                 wire1305,
                 (1'h0)};
  assign wire1305 = $unsigned($signed(($signed(wire1300[(3'h5):(1'h0)]) && $signed(wire1300[(3'h7):(3'h5)]))));
  assign wire1306 = wire1302[(1'h1):(1'h0)];
  assign wire1307 = ($unsigned((~|(^(~^wire1302)))) ?
                        $signed($unsigned((|(wire1304 ?
                            wire1305 : wire1300)))) : $signed($unsigned((wire1301[(2'h2):(1'h1)] && (~&wire1305)))));
  assign wire1308 = {(wire1304[(5'h10):(5'h10)] ?
                            (wire1302 <<< $unsigned((~wire1305))) : $signed({$unsigned(wire1305)}))};
  assign wire1309 = $signed((~|wire1304[(2'h2):(2'h2)]));
  assign wire1310 = wire1303;
  assign wire1311 = (~^$signed({(wire1302 ?
                            $unsigned(wire1307) : (wire1305 >>> wire1301)),
                        wire1301[(4'h9):(2'h2)]}));
  assign wire1312 = $unsigned({wire1305[(3'h6):(2'h3)]});
  assign wire1313 = ($unsigned($unsigned($signed(wire1306))) < (wire1306[(3'h5):(3'h4)] <= $unsigned((wire1305[(3'h4):(1'h0)] ?
                        $signed(wire1305) : ((8'hb0) ? wire1309 : wire1304)))));
  assign wire1314 = wire1311;
  assign wire1315 = {{wire1302[(3'h4):(3'h4)],
                            $signed(((wire1311 >> wire1304) ^~ {wire1301}))},
                        $signed(wire1303)};
  assign wire1316 = (($unsigned({wire1309[(4'hb):(3'h6)]}) ?
                        ((~^$unsigned(wire1312)) || wire1309) : $signed(wire1309)) & $unsigned((~|$unsigned(wire1300))));
  assign wire1317 = {$unsigned($signed(((wire1301 == wire1305) - wire1310[(1'h1):(1'h0)]))),
                        wire1307};
  assign wire1318 = {wire1302, ((^($unsigned((8'hb5)) ^ wire1306)) & (8'hb4))};
  always
    @(posedge clk) begin
      reg1319 <= wire1310;
      reg1320 <= $unsigned($unsigned((($signed(wire1301) ?
              $unsigned(wire1313) : $unsigned(wire1317)) ?
          ($signed(wire1305) ?
              {wire1309} : $signed(wire1309)) : wire1308[(3'h5):(3'h4)])));
    end
  assign wire1321 = ((^~(($signed(wire1315) ?
                            $signed(wire1304) : $signed(wire1305)) ?
                        ($unsigned(wire1306) >= (~^wire1304)) : ((wire1308 ?
                            wire1311 : (8'hac)) > wire1312[(4'hd):(1'h0)]))) * (wire1314[(4'he):(4'ha)] ?
                        wire1305[(4'hf):(1'h1)] : {($signed((8'haa)) <<< (-wire1315)),
                            (^wire1318)}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1222
#( parameter param1291 = ((({{(8'hbe)}, {(7'h42)}} ? {(+(8'hb7)), ((8'hbc) * (8'hba))} : (((8'haf) ? (8'haa) : (8'ha1)) ? ((8'haa) ? (8'h9d) : (7'h43)) : ((8'ha8) != (8'ha8)))) << ({(~|(7'h40))} >>> (((7'h43) > (8'hbc)) ? ((8'ha9) || (7'h41)) : ((8'hb1) | (8'haf))))) > (^~(((~|(8'hbd)) && ((8'hb7) ? (8'ha1) : (8'hbd))) ? ((|(8'ha4)) ? (8'had) : {(8'hb1), (8'hbb)}) : {{(8'hab)}, (^~(8'hb8))})))
, parameter param1292 = ((param1291 ? (((param1291 ? param1291 : param1291) > (param1291 | param1291)) ? ((param1291 & param1291) ? (param1291 ? param1291 : param1291) : (param1291 ? param1291 : param1291)) : ((^param1291) ? ((8'hbb) ~^ param1291) : {param1291})) : param1291) ^ {(param1291 <<< (~|param1291)), {param1291}}) )
(y, clk, wire1227, wire1226, wire1225, wire1224, wire1223);
  output wire [(32'h284):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire1227;
  input wire signed [(3'h6):(1'h0)] wire1226;
  input wire [(4'ha):(1'h0)] wire1225;
  input wire [(4'ha):(1'h0)] wire1224;
  input wire [(5'h10):(1'h0)] wire1223;
  reg [(5'h10):(1'h0)] reg1290 = (1'h0);
  reg [(3'h6):(1'h0)] reg1289 = (1'h0);
  reg [(3'h7):(1'h0)] reg1288 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1287 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1286 = (1'h0);
  reg [(4'ha):(1'h0)] reg1285 = (1'h0);
  reg [(4'ha):(1'h0)] reg1284 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1283 = (1'h0);
  reg [(2'h3):(1'h0)] reg1282 = (1'h0);
  reg [(5'h12):(1'h0)] reg1281 = (1'h0);
  reg [(2'h2):(1'h0)] reg1280 = (1'h0);
  reg [(5'h15):(1'h0)] reg1279 = (1'h0);
  reg [(4'ha):(1'h0)] reg1278 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1277 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1276 = (1'h0);
  reg [(3'h6):(1'h0)] reg1275 = (1'h0);
  reg [(4'h8):(1'h0)] reg1274 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1273 = (1'h0);
  reg [(3'h7):(1'h0)] reg1272 = (1'h0);
  reg [(3'h6):(1'h0)] reg1271 = (1'h0);
  reg [(4'hc):(1'h0)] reg1270 = (1'h0);
  reg [(4'hb):(1'h0)] reg1269 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1268 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1267 = (1'h0);
  reg [(4'ha):(1'h0)] reg1266 = (1'h0);
  reg [(5'h10):(1'h0)] reg1265 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1264 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1263 = (1'h0);
  reg [(2'h3):(1'h0)] reg1262 = (1'h0);
  reg [(4'hb):(1'h0)] reg1261 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1260 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1259 = (1'h0);
  reg [(2'h3):(1'h0)] reg1258 = (1'h0);
  reg [(3'h6):(1'h0)] reg1257 = (1'h0);
  reg [(4'h9):(1'h0)] reg1256 = (1'h0);
  reg [(2'h2):(1'h0)] reg1255 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1254 = (1'h0);
  reg [(2'h3):(1'h0)] reg1253 = (1'h0);
  wire [(4'h9):(1'h0)] wire1252;
  wire [(5'h11):(1'h0)] wire1251;
  reg [(3'h4):(1'h0)] reg1250 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1249 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1248 = (1'h0);
  reg [(2'h3):(1'h0)] reg1247 = (1'h0);
  reg [(4'hd):(1'h0)] reg1246 = (1'h0);
  reg [(4'hd):(1'h0)] reg1245 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1244 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1243 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1242 = (1'h0);
  reg [(5'h11):(1'h0)] reg1241 = (1'h0);
  reg [(4'hf):(1'h0)] reg1240 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1239 = (1'h0);
  reg [(4'hf):(1'h0)] reg1238 = (1'h0);
  reg [(4'h8):(1'h0)] reg1237 = (1'h0);
  reg [(3'h5):(1'h0)] reg1236 = (1'h0);
  reg [(3'h5):(1'h0)] reg1235 = (1'h0);
  reg [(3'h5):(1'h0)] reg1234 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1233 = (1'h0);
  reg [(4'hc):(1'h0)] reg1232 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1231 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1230 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1229 = (1'h0);
  wire [(4'he):(1'h0)] wire1228;
  assign y = {reg1290,
                 reg1289,
                 reg1288,
                 reg1287,
                 reg1286,
                 reg1285,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1281,
                 reg1280,
                 reg1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 reg1275,
                 reg1274,
                 reg1273,
                 reg1272,
                 reg1271,
                 reg1270,
                 reg1269,
                 reg1268,
                 reg1267,
                 reg1266,
                 reg1265,
                 reg1264,
                 reg1263,
                 reg1262,
                 reg1261,
                 reg1260,
                 reg1259,
                 reg1258,
                 reg1257,
                 reg1256,
                 reg1255,
                 reg1254,
                 reg1253,
                 wire1252,
                 wire1251,
                 reg1250,
                 reg1249,
                 reg1248,
                 reg1247,
                 reg1246,
                 reg1245,
                 reg1244,
                 reg1243,
                 reg1242,
                 reg1241,
                 reg1240,
                 reg1239,
                 reg1238,
                 reg1237,
                 reg1236,
                 reg1235,
                 reg1234,
                 reg1233,
                 reg1232,
                 reg1231,
                 reg1230,
                 reg1229,
                 wire1228,
                 (1'h0)};
  assign wire1228 = $signed((~((~^wire1224[(3'h6):(2'h3)]) >> $signed((wire1223 ?
                        wire1223 : (8'hb8))))));
  always
    @(posedge clk) begin
      reg1229 <= ((-$signed({wire1226[(2'h2):(1'h1)],
          $signed(wire1223)})) ^ wire1223);
      if (wire1225)
        begin
          reg1230 <= wire1224;
          reg1231 <= $signed(wire1223);
          reg1232 <= $unsigned(((wire1228[(4'h8):(3'h5)] | ((wire1227 == wire1223) ?
                  wire1225[(3'h5):(2'h3)] : (wire1227 ? (7'h44) : wire1223))) ?
              $signed($unsigned(wire1225[(4'ha):(4'h9)])) : wire1223));
          reg1233 <= $unsigned({wire1227});
          if ($signed($unsigned((reg1229[(2'h3):(1'h1)] ?
              reg1229 : (~&reg1233[(2'h2):(2'h2)])))))
            begin
              reg1234 <= ($unsigned(reg1229[(1'h1):(1'h0)]) ?
                  reg1230 : $signed((8'ha6)));
              reg1235 <= reg1229;
            end
          else
            begin
              reg1234 <= (^~(~|reg1232[(1'h1):(1'h1)]));
              reg1235 <= ((&reg1230[(5'h10):(2'h2)]) != $unsigned(($unsigned($unsigned((8'ha4))) ?
                  (reg1231 ?
                      wire1228 : ((8'hb4) ?
                          reg1229 : wire1226)) : (|$signed(reg1231)))));
              reg1236 <= reg1232;
              reg1237 <= $unsigned(($signed(wire1224) ?
                  wire1225 : (wire1224 >>> wire1226)));
            end
        end
      else
        begin
          if (((~^$signed((~|(reg1233 ? wire1224 : reg1234)))) >> (7'h40)))
            begin
              reg1230 <= reg1233;
              reg1231 <= ($unsigned($signed((reg1230[(2'h2):(1'h1)] ?
                  (reg1231 ? wire1225 : wire1224) : {wire1225,
                      wire1226}))) + $signed(($signed(reg1235[(2'h2):(1'h0)]) < ((reg1235 | reg1236) ?
                  wire1228 : wire1226))));
            end
          else
            begin
              reg1230 <= wire1227;
              reg1231 <= ($unsigned(($unsigned(reg1233) ?
                      reg1229 : $signed((reg1232 || wire1228)))) ?
                  reg1236 : $unsigned({$signed((reg1230 > reg1236)),
                      ((reg1236 ?
                          (7'h41) : reg1231) - (wire1223 && reg1234))}));
            end
        end
      reg1238 <= ({{($unsigned(wire1227) >>> (reg1229 ? reg1236 : wire1226)),
                  (~^((7'h42) ? (7'h41) : reg1229))},
              ({$unsigned(wire1225)} ~^ (+(-reg1234)))} ?
          $unsigned((-$unsigned(reg1237))) : reg1229);
      reg1239 <= reg1235[(2'h2):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg1240 <= {((7'h42) ?
              reg1235[(1'h0):(1'h0)] : (($signed(reg1237) ?
                      (~|wire1228) : wire1228) ?
                  {(reg1230 ? reg1237 : wire1228), reg1229} : wire1227)),
          (reg1232 != $unsigned($signed($unsigned(wire1227))))};
      if ((|{({(reg1235 ? reg1238 : reg1239)} * $signed(reg1240))}))
        begin
          reg1241 <= reg1232;
          reg1242 <= (($unsigned(reg1231[(3'h6):(1'h0)]) & wire1227[(2'h2):(2'h2)]) ?
              $unsigned((!(!$signed((8'hba))))) : reg1236[(3'h4):(2'h3)]);
          reg1243 <= wire1228[(3'h7):(2'h2)];
        end
      else
        begin
          reg1241 <= (8'hb9);
          reg1242 <= {reg1229[(1'h0):(1'h0)]};
          reg1243 <= {(!reg1229[(1'h0):(1'h0)]),
              (wire1227 ?
                  $unsigned(($signed(reg1239) != (|reg1240))) : reg1233[(1'h1):(1'h0)])};
          reg1244 <= ((+$unsigned($signed($unsigned(wire1224)))) ?
              {((reg1234[(2'h2):(1'h1)] ~^ $signed(reg1234)) ?
                      $unsigned((^reg1231)) : reg1234)} : wire1224);
          reg1245 <= ((reg1238[(2'h3):(2'h3)] ?
                  wire1224[(2'h3):(2'h2)] : (8'had)) ?
              (^~(|(&wire1227))) : reg1240[(4'hc):(4'ha)]);
        end
      if ({{(({reg1235, reg1241} ^ $unsigned((8'hb7))) ?
                  (!{(8'hb6)}) : ((wire1226 * reg1236) ?
                      {reg1234, reg1244} : $unsigned(wire1226))),
              (($signed(wire1224) ?
                  wire1223[(4'ha):(2'h3)] : $signed(reg1240)) << $signed($signed((8'ha8))))},
          {(wire1225[(1'h1):(1'h1)] ? wire1227 : $unsigned({reg1233, reg1233})),
              ($signed((wire1227 ?
                  wire1224 : wire1228)) >> $unsigned($unsigned(reg1233)))}})
        begin
          reg1246 <= $signed((reg1243 <<< $signed(reg1241)));
        end
      else
        begin
          reg1246 <= $signed(reg1233[(2'h2):(1'h1)]);
          reg1247 <= (&reg1243[(1'h1):(1'h0)]);
          reg1248 <= (~&((-(~^$unsigned(wire1223))) == (wire1224[(3'h5):(1'h0)] ?
              (8'hb7) : wire1227[(4'hd):(2'h2)])));
          reg1249 <= ($unsigned($signed(reg1247)) ?
              reg1235 : (((^~(-wire1227)) ?
                  ($signed(reg1241) || (wire1225 < reg1236)) : $signed($signed(reg1238))) == $unsigned(reg1245)));
          reg1250 <= wire1225;
        end
    end
  assign wire1251 = $unsigned((((~&$signed((8'ha2))) ^ ($signed(reg1241) ?
                            ((8'hae) ? reg1232 : reg1248) : (~reg1250))) ?
                        ($unsigned($signed(reg1233)) - ({reg1238} + (!reg1241))) : $signed((~^{wire1223,
                            reg1233}))));
  assign wire1252 = ({($unsigned($unsigned(reg1245)) ?
                                (!(wire1227 ?
                                    reg1246 : wire1225)) : $unsigned(reg1235))} ?
                        $signed(reg1250[(1'h0):(1'h0)]) : reg1250[(2'h2):(1'h0)]);
  always
    @(posedge clk) begin
      if ({$unsigned({(((8'hba) ? reg1230 : reg1236) ?
                  reg1241 : {reg1250, (8'hbe)})}),
          reg1238})
        begin
          reg1253 <= $signed(($signed($signed((reg1231 != reg1248))) ?
              reg1229[(2'h3):(2'h3)] : ($unsigned($signed(wire1251)) ?
                  ((~reg1242) ?
                      (wire1251 ? reg1242 : reg1230) : (8'ha5)) : reg1248)));
          reg1254 <= ((~$signed($unsigned(reg1253[(1'h1):(1'h1)]))) > reg1238[(4'hc):(3'h6)]);
          if ($unsigned(reg1243[(1'h0):(1'h0)]))
            begin
              reg1255 <= reg1248;
            end
          else
            begin
              reg1255 <= reg1239;
              reg1256 <= (($signed($signed(reg1249)) ?
                  (~reg1248[(3'h4):(2'h3)]) : {(+$signed(reg1240))}) & reg1255[(1'h0):(1'h0)]);
              reg1257 <= reg1247;
            end
          if (wire1226[(3'h6):(3'h5)])
            begin
              reg1258 <= $unsigned((+((~|$signed(wire1223)) >>> (|reg1238[(4'hf):(2'h3)]))));
              reg1259 <= reg1245;
            end
          else
            begin
              reg1258 <= reg1230[(5'h12):(5'h10)];
              reg1259 <= ($signed((~^reg1242)) ?
                  reg1243 : (((^~$signed(wire1227)) >= ($unsigned((8'hbc)) ?
                          reg1257 : reg1237[(1'h0):(1'h0)])) ?
                      (((&reg1255) & $unsigned((8'hb6))) ?
                          ({reg1230} ?
                              $unsigned(wire1225) : wire1223) : (!{reg1257})) : (($signed(reg1233) >> reg1238) <<< $signed(((8'ha7) << wire1225)))));
              reg1260 <= (7'h40);
              reg1261 <= reg1235;
              reg1262 <= reg1244;
            end
          if (reg1242)
            begin
              reg1263 <= ($unsigned(reg1236) | $unsigned((^~(wire1223[(3'h6):(3'h4)] - ((8'hac) && reg1261)))));
              reg1264 <= $unsigned((^wire1225));
              reg1265 <= reg1253;
            end
          else
            begin
              reg1263 <= $unsigned($unsigned(reg1234));
              reg1264 <= $signed((reg1258[(2'h2):(1'h0)] > (&reg1248)));
              reg1265 <= (-(reg1235[(3'h4):(1'h1)] >= $signed($signed((reg1261 ?
                  reg1255 : reg1262)))));
              reg1266 <= $signed($unsigned($unsigned($unsigned(reg1240[(3'h5):(1'h1)]))));
              reg1267 <= ($unsigned(reg1263) ?
                  (~(reg1245 ?
                      ((&(8'hb2)) >= (&(8'h9e))) : $signed(reg1239))) : {({{reg1263,
                              (8'haa)}} * reg1253[(2'h2):(1'h0)]),
                      ({{(8'hbf)}, reg1236} ?
                          $unsigned(reg1238[(2'h2):(1'h0)]) : $unsigned($signed(wire1223)))});
            end
        end
      else
        begin
          reg1253 <= reg1239;
          if ($unsigned((reg1237 ?
              reg1254 : ($signed($signed(reg1265)) ?
                  (reg1257 ?
                      (~^(8'hbe)) : wire1227[(5'h10):(2'h2)]) : (^~$unsigned(reg1265))))))
            begin
              reg1254 <= (!$signed((-{$signed(reg1245), (reg1235 & reg1243)})));
              reg1255 <= reg1233[(2'h2):(2'h2)];
            end
          else
            begin
              reg1254 <= ((reg1230[(3'h7):(2'h2)] << $signed(((reg1249 | reg1262) ?
                      (reg1231 || reg1254) : wire1228[(3'h5):(3'h4)]))) ?
                  reg1241 : $unsigned($signed((reg1250[(2'h3):(2'h3)] ?
                      (~&(7'h41)) : (reg1230 >>> wire1228)))));
              reg1255 <= (!$unsigned($unsigned(((|reg1248) ?
                  wire1228[(4'ha):(4'ha)] : $unsigned(reg1236)))));
            end
        end
      reg1268 <= (reg1249[(3'h4):(1'h0)] || reg1243);
      if (reg1264)
        begin
          reg1269 <= {wire1226};
          if (reg1260)
            begin
              reg1270 <= (({(8'hb5), (~&$signed((8'haf)))} ?
                      {reg1257[(3'h6):(2'h2)]} : ($signed($unsigned(reg1253)) ?
                          (-(reg1264 ?
                              wire1252 : reg1257)) : {(reg1264 > reg1239),
                              reg1235})) ?
                  (8'hb9) : {$unsigned((~^{reg1269, wire1223})),
                      reg1239[(3'h6):(1'h1)]});
              reg1271 <= wire1225;
              reg1272 <= (reg1242 <= ({{reg1234[(3'h4):(1'h0)]}} >= $signed(reg1246[(1'h1):(1'h0)])));
            end
          else
            begin
              reg1270 <= $signed(reg1269[(3'h6):(2'h3)]);
              reg1271 <= {(reg1253[(2'h3):(2'h2)] ?
                      $signed((+$unsigned(wire1228))) : (wire1228 != $unsigned($unsigned(reg1241)))),
                  {((wire1225[(3'h7):(1'h1)] == ((8'hb2) ?
                          reg1238 : reg1259)) & (~&$signed(reg1239))),
                      reg1248[(4'hb):(4'hb)]}};
              reg1272 <= (8'h9c);
            end
          reg1273 <= $unsigned((^{(^~(reg1253 || reg1264))}));
          reg1274 <= (reg1247[(1'h0):(1'h0)] << $signed({wire1226[(2'h2):(1'h1)]}));
          if (wire1224)
            begin
              reg1275 <= {(+wire1224),
                  $unsigned($unsigned(((reg1255 ?
                      reg1243 : reg1242) <= $unsigned((8'hbb)))))};
              reg1276 <= reg1273;
              reg1277 <= $signed($signed(((reg1266 ?
                  {reg1234,
                      reg1246} : reg1230) ^ $signed(reg1240[(3'h6):(1'h0)]))));
              reg1278 <= {reg1243[(2'h3):(2'h2)]};
              reg1279 <= wire1224;
            end
          else
            begin
              reg1275 <= $signed(wire1224);
              reg1276 <= (reg1259 ?
                  (($signed(reg1248) | (-(reg1257 ? wire1228 : reg1266))) ?
                      reg1233 : (8'ha3)) : {$unsigned(reg1254)});
              reg1277 <= reg1254;
            end
        end
      else
        begin
          if (reg1275[(3'h4):(1'h0)])
            begin
              reg1269 <= (-((-$signed(reg1267)) ?
                  wire1226 : {reg1258[(1'h0):(1'h0)]}));
            end
          else
            begin
              reg1269 <= (^~reg1278[(3'h6):(2'h2)]);
              reg1270 <= reg1230[(1'h0):(1'h0)];
            end
          reg1271 <= $unsigned(((&((reg1230 ? (8'hb8) : reg1264) ?
              wire1223[(4'h9):(1'h0)] : $signed(reg1234))) + reg1277));
        end
      reg1280 <= (reg1235 - $signed(reg1244[(3'h7):(1'h1)]));
    end
  always
    @(posedge clk) begin
      if (reg1253)
        begin
          reg1281 <= $signed((|$signed(reg1278[(1'h0):(1'h0)])));
          reg1282 <= (&(reg1255[(1'h0):(1'h0)] ?
              reg1250[(2'h2):(2'h2)] : reg1231));
          reg1283 <= {reg1269[(4'ha):(4'h8)]};
        end
      else
        begin
          if ($unsigned(reg1265[(4'ha):(2'h2)]))
            begin
              reg1281 <= ($unsigned(reg1242[(4'hb):(4'ha)]) ?
                  (!((~{reg1264, reg1239}) ?
                      $unsigned((|reg1229)) : reg1277)) : (reg1242[(3'h4):(2'h2)] ?
                      $unsigned(({reg1244} ?
                          $unsigned(reg1250) : $signed(reg1270))) : $unsigned(($signed((8'hb2)) > ((8'ha3) ?
                          reg1270 : wire1225)))));
              reg1282 <= ($unsigned($unsigned($unsigned((reg1275 ?
                      reg1236 : wire1228)))) ?
                  ($signed({(reg1236 ? reg1235 : wire1227),
                          (reg1236 ? reg1234 : reg1253)}) ?
                      ({(reg1254 ?
                              wire1225 : reg1243)} ^ reg1242) : $signed(reg1276)) : $signed({{(wire1228 ?
                              reg1250 : reg1264),
                          $signed(reg1282)},
                      {(reg1256 ? reg1235 : reg1265), reg1240}}));
              reg1283 <= reg1234;
              reg1284 <= wire1251[(5'h10):(4'he)];
              reg1285 <= {$signed(reg1281[(5'h11):(4'hf)]), $unsigned(reg1242)};
            end
          else
            begin
              reg1281 <= (({(|(reg1248 + wire1224))} ?
                  (reg1269 >>> (((8'ha8) * reg1240) ^ $unsigned(reg1241))) : {($unsigned(reg1278) ?
                          $unsigned(wire1226) : $unsigned((8'hb4)))}) << $signed($unsigned((reg1261[(4'h8):(4'h8)] || (reg1248 * reg1242)))));
              reg1282 <= $unsigned((+$signed((&((8'hb8) ?
                  reg1242 : wire1224)))));
              reg1283 <= $unsigned(reg1233[(1'h1):(1'h1)]);
            end
        end
      if (({$unsigned(reg1232)} >= (&$signed($signed((8'hb3))))))
        begin
          if ((~^(((~reg1253[(1'h0):(1'h0)]) ?
              ($unsigned(reg1273) ?
                  reg1272[(2'h2):(2'h2)] : $signed(reg1253)) : $signed((reg1244 ?
                  (8'ha0) : reg1265))) >= reg1232)))
            begin
              reg1286 <= reg1237[(3'h7):(3'h5)];
              reg1287 <= (reg1231 << $signed({(|(wire1223 < reg1286))}));
              reg1288 <= $unsigned(($signed($signed($signed((8'ha9)))) ?
                  $unsigned($signed(reg1241)) : (reg1283[(3'h4):(1'h0)] ?
                      reg1284[(3'h4):(1'h1)] : (reg1240[(4'ha):(2'h3)] ?
                          $unsigned(reg1237) : reg1246[(2'h3):(1'h1)]))));
            end
          else
            begin
              reg1286 <= $unsigned(reg1265[(2'h3):(1'h0)]);
              reg1287 <= reg1280[(2'h2):(1'h1)];
              reg1288 <= $signed(($signed($unsigned((reg1264 ?
                  reg1280 : reg1235))) & (!(reg1258[(2'h2):(2'h2)] ?
                  $unsigned((8'hba)) : (reg1255 ? reg1229 : reg1246)))));
            end
          reg1289 <= reg1287[(1'h1):(1'h1)];
          reg1290 <= reg1259[(3'h6):(3'h6)];
        end
      else
        begin
          reg1286 <= reg1275[(3'h6):(3'h5)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1354
#( parameter param1383 = ((~&(~(+((8'hb1) ? (8'hb9) : (8'had))))) ? (((((8'hb6) < (8'ha7)) == ((8'hbe) <<< (8'hbc))) ? (~&(~&(8'hb8))) : ((^(8'hbc)) ^ {(8'ha1)})) || (+(8'h9e))) : (((|{(8'hbb), (8'hab)}) >> ({(8'hb2), (8'haf)} ? {(8'h9d), (7'h42)} : ((7'h40) ? (8'ha6) : (7'h40)))) + (+((^~(8'haf)) ? ((8'hb3) <= (8'hac)) : ((8'haa) ? (8'had) : (8'ha4)))))) )
(y, clk, wire1358, wire1357, wire1356, wire1355);
  output wire [(32'h43):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire1358;
  input wire [(4'h8):(1'h0)] wire1357;
  input wire signed [(4'hb):(1'h0)] wire1356;
  input wire [(5'h11):(1'h0)] wire1355;
  wire signed [(5'h10):(1'h0)] wire1382;
  wire signed [(5'h13):(1'h0)] wire1380;
  wire [(5'h12):(1'h0)] wire1360;
  wire signed [(4'hd):(1'h0)] wire1359;
  assign y = {wire1382, wire1380, wire1360, wire1359, (1'h0)};
  assign wire1359 = $signed(wire1355);
  assign wire1360 = $signed(wire1357);
  module1361 modinst1381 (.wire1365(wire1355), .clk(clk), .y(wire1380), .wire1364(wire1357), .wire1363(wire1360), .wire1362(wire1359));
  assign wire1382 = $signed({(^~wire1356[(2'h2):(2'h2)])});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1361
#( parameter param1378 = ((((-{(8'had), (7'h44)}) ? (-((8'haa) ? (7'h40) : (8'ha7))) : (((8'hac) ? (8'hae) : (8'ha8)) ? ((7'h43) >= (8'ha9)) : (&(8'hb0)))) >> ({((8'hbe) - (8'hbb)), ((7'h42) ? (8'hb9) : (8'hab))} | {{(8'hb7), (8'hb2)}, ((8'haf) ? (8'hbe) : (8'hba))})) ? ((^~(-((8'ha5) ? (8'hbf) : (8'hb0)))) >> ((((8'haf) != (8'hbe)) ? ((8'hb8) <<< (8'ha8)) : {(8'ha9), (8'hbb)}) ? (~^((8'haf) ? (8'hba) : (8'ha2))) : {((8'hb4) ? (8'hb9) : (8'haf))})) : (((((8'ha6) > (8'hbd)) ? (^~(8'hb9)) : ((8'hb7) ? (8'hbd) : (8'hab))) >>> (((8'ha0) || (7'h43)) ? {(8'hb3)} : (~^(8'ha4)))) ? (((~&(8'haf)) | (!(8'hbf))) ? (((8'h9f) >>> (8'ha4)) ? (~&(8'ha0)) : (~^(7'h40))) : {(^(8'hbb))}) : (((^(8'h9f)) ? ((8'ha8) || (8'h9d)) : ((8'hb5) ~^ (8'hae))) ? ((~(7'h42)) >> {(8'hb5)}) : (((8'ha7) ? (8'ha0) : (8'hb6)) != ((7'h40) ? (8'hb3) : (8'haa))))))
, parameter param1379 = (^((((param1378 ? (8'hb2) : param1378) ? (param1378 ? (8'had) : param1378) : param1378) || (~|{param1378})) > ((8'haa) * ((param1378 ? param1378 : param1378) && (param1378 ^~ param1378))))) )
(y, clk, wire1365, wire1364, wire1363, wire1362);
  output wire [(32'h9f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire1365;
  input wire signed [(4'h8):(1'h0)] wire1364;
  input wire [(2'h3):(1'h0)] wire1363;
  input wire signed [(4'hd):(1'h0)] wire1362;
  wire [(5'h13):(1'h0)] wire1377;
  wire signed [(5'h15):(1'h0)] wire1376;
  wire [(5'h11):(1'h0)] wire1375;
  wire [(3'h6):(1'h0)] wire1374;
  reg [(2'h3):(1'h0)] reg1373 = (1'h0);
  reg [(5'h14):(1'h0)] reg1372 = (1'h0);
  reg [(5'h11):(1'h0)] reg1371 = (1'h0);
  reg [(2'h3):(1'h0)] reg1370 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1369 = (1'h0);
  wire [(4'hf):(1'h0)] wire1368;
  wire [(4'h9):(1'h0)] wire1367;
  wire signed [(5'h15):(1'h0)] wire1366;
  assign y = {wire1377,
                 wire1376,
                 wire1375,
                 wire1374,
                 reg1373,
                 reg1372,
                 reg1371,
                 reg1370,
                 reg1369,
                 wire1368,
                 wire1367,
                 wire1366,
                 (1'h0)};
  assign wire1366 = wire1363[(2'h2):(2'h2)];
  assign wire1367 = ($signed(wire1365[(3'h7):(2'h3)]) >>> wire1366);
  assign wire1368 = $unsigned(wire1362[(4'hb):(3'h6)]);
  always
    @(posedge clk) begin
      if ((^(^~(~&(~^{wire1363})))))
        begin
          if ($signed($unsigned({$unsigned(wire1363)})))
            begin
              reg1369 <= {wire1366, wire1363[(1'h1):(1'h0)]};
            end
          else
            begin
              reg1369 <= ({wire1367[(4'h8):(3'h5)]} ?
                  wire1366 : ($unsigned(($signed(wire1364) & (~wire1365))) ?
                      wire1363 : $unsigned((wire1367 ?
                          (~reg1369) : wire1365[(4'hb):(4'hb)]))));
              reg1370 <= wire1368;
              reg1371 <= $signed($signed((({wire1365} ?
                      {wire1367} : ((7'h43) ^~ reg1370)) ?
                  $signed(((8'hb9) <<< reg1370)) : {$signed((8'ha5)),
                      (~wire1366)})));
              reg1372 <= wire1363;
            end
          reg1373 <= wire1367[(3'h4):(3'h4)];
        end
      else
        begin
          reg1369 <= reg1371[(2'h3):(2'h2)];
        end
    end
  assign wire1374 = ($unsigned($signed(wire1367)) ?
                        (8'hbf) : (($signed((8'ha4)) ?
                                reg1369[(2'h3):(1'h1)] : $signed(reg1373)) ?
                            ((wire1365[(4'hc):(3'h4)] ?
                                    reg1373[(2'h2):(1'h0)] : (8'hb2)) ?
                                (8'hb8) : $unsigned((~|wire1363))) : (^~($signed(reg1371) * $signed(wire1362)))));
  assign wire1375 = ($signed({wire1367[(1'h0):(1'h0)],
                        $signed((reg1371 ^ reg1369))}) + $signed(reg1371[(4'ha):(3'h4)]));
  assign wire1376 = (reg1372[(1'h1):(1'h1)] ?
                        ($signed(((~|reg1370) ^ (wire1375 <= reg1369))) ?
                            wire1368[(4'he):(4'h8)] : wire1374) : wire1364);
  assign wire1377 = ((({$signed(wire1362)} >>> ((wire1366 ?
                                wire1365 : reg1370) ?
                            (8'hb3) : $signed(reg1372))) ?
                        $unsigned((~$unsigned(reg1371))) : wire1367) ~^ $unsigned((wire1367[(4'h9):(4'h8)] ?
                        $signed((8'hbd)) : (^~$unsigned((8'ha9))))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1884  (y, clk, wire1888, wire1887, wire1886, wire1885);
  output wire [(32'h85):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire1888;
  input wire [(4'hf):(1'h0)] wire1887;
  input wire signed [(5'h13):(1'h0)] wire1886;
  input wire [(3'h7):(1'h0)] wire1885;
  wire [(2'h3):(1'h0)] wire1902;
  wire [(3'h6):(1'h0)] wire1901;
  wire [(5'h14):(1'h0)] wire1900;
  wire [(2'h3):(1'h0)] wire1899;
  wire signed [(5'h11):(1'h0)] wire1898;
  wire signed [(3'h5):(1'h0)] wire1897;
  wire [(3'h6):(1'h0)] wire1896;
  wire signed [(4'h8):(1'h0)] wire1895;
  wire signed [(5'h11):(1'h0)] wire1894;
  wire signed [(3'h7):(1'h0)] wire1893;
  reg [(3'h6):(1'h0)] reg1892 = (1'h0);
  reg [(4'ha):(1'h0)] reg1891 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1890 = (1'h0);
  wire [(4'ha):(1'h0)] wire1889;
  assign y = {wire1902,
                 wire1901,
                 wire1900,
                 wire1899,
                 wire1898,
                 wire1897,
                 wire1896,
                 wire1895,
                 wire1894,
                 wire1893,
                 reg1892,
                 reg1891,
                 reg1890,
                 wire1889,
                 (1'h0)};
  assign wire1889 = ($signed($unsigned({$unsigned(wire1888), wire1886})) ?
                        $signed(wire1887) : (^$signed(wire1888)));
  always
    @(posedge clk) begin
      reg1890 <= (wire1888[(1'h0):(1'h0)] == (^~wire1886));
      reg1891 <= (8'haf);
      reg1892 <= wire1889;
    end
  assign wire1893 = (^reg1892[(3'h4):(1'h0)]);
  assign wire1894 = (&(^$unsigned((wire1888[(2'h2):(1'h0)] != $signed(reg1891)))));
  assign wire1895 = (~(~^(~|$signed((+(8'hbc))))));
  assign wire1896 = (wire1889 * {$unsigned(wire1895)});
  assign wire1897 = $signed((-wire1887));
  assign wire1898 = (|$signed((wire1893[(3'h6):(3'h5)] ?
                        $signed($unsigned(wire1887)) : $unsigned((wire1889 ?
                            wire1885 : wire1885)))));
  assign wire1899 = $unsigned($signed({(wire1889 | (wire1894 ?
                            wire1887 : wire1896))}));
  assign wire1900 = $signed((~^$unsigned($unsigned($signed(reg1891)))));
  assign wire1901 = ((~wire1900[(1'h1):(1'h1)]) > reg1892[(1'h1):(1'h1)]);
  assign wire1902 = $unsigned($unsigned($signed($unsigned((&wire1887)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1760
#( parameter param1876 = ((7'h40) ? ((-{(~(8'hb8)), ((8'ha6) ? (8'had) : (7'h42))}) ? ({((8'hac) >>> (8'hb0))} ? ((~|(8'hae)) ? {(8'ha5), (8'hb7)} : (~|(8'ha1))) : (((8'h9f) ? (8'hb2) : (8'h9c)) ? (^~(8'had)) : (8'ha9))) : ((((8'haf) ? (8'hbb) : (8'hb1)) ? ((8'ha1) ^~ (8'ha8)) : ((8'hae) ? (8'hb7) : (8'ha8))) ? (8'hb7) : (((8'hb1) >>> (8'h9d)) ? ((7'h40) >>> (8'hab)) : ((8'h9f) ^ (8'hba))))) : {((|((8'hb8) ? (8'hac) : (7'h43))) ? (8'ha4) : (((8'ha0) ? (8'hb0) : (8'hbc)) ? (~|(8'hbe)) : (^~(8'hb4)))), (^~(!(~&(8'hae))))})
, parameter param1877 = (((~param1876) ? (param1876 ? ({param1876, param1876} >> (8'h9c)) : (~&(param1876 ? param1876 : param1876))) : param1876) - (-((~(~param1876)) < ((~^param1876) ? param1876 : {param1876, param1876})))) )
(y, clk, wire1761, wire1762, wire1763, wire1764, wire1765);
  output wire [(32'h34e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire1761;
  input wire [(5'h10):(1'h0)] wire1762;
  input wire [(5'h10):(1'h0)] wire1763;
  input wire signed [(5'h12):(1'h0)] wire1764;
  input wire [(5'h15):(1'h0)] wire1765;
  wire signed [(5'h11):(1'h0)] wire1875;
  wire signed [(4'ha):(1'h0)] wire1874;
  wire [(5'h12):(1'h0)] wire1873;
  reg [(4'he):(1'h0)] reg1872 = (1'h0);
  reg [(2'h3):(1'h0)] reg1871 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1870 = (1'h0);
  reg [(4'h9):(1'h0)] reg1869 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1868 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1867 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1866 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1865 = (1'h0);
  reg [(5'h10):(1'h0)] reg1864 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1863 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1862 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1861 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1860 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1859 = (1'h0);
  reg [(3'h7):(1'h0)] reg1858 = (1'h0);
  reg [(4'hf):(1'h0)] reg1857 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1856 = (1'h0);
  reg [(5'h12):(1'h0)] reg1855 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1854 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1853 = (1'h0);
  reg [(5'h11):(1'h0)] reg1852 = (1'h0);
  reg [(3'h6):(1'h0)] reg1851 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1850 = (1'h0);
  reg [(5'h12):(1'h0)] reg1849 = (1'h0);
  reg [(2'h3):(1'h0)] reg1848 = (1'h0);
  reg [(3'h5):(1'h0)] reg1847 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire1846;
  wire [(4'hc):(1'h0)] wire1845;
  wire signed [(3'h5):(1'h0)] wire1844;
  reg signed [(5'h10):(1'h0)] reg1843 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1842 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1841 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1840 = (1'h0);
  reg [(2'h3):(1'h0)] reg1839 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1838 = (1'h0);
  reg [(2'h3):(1'h0)] reg1837 = (1'h0);
  reg [(2'h3):(1'h0)] reg1836 = (1'h0);
  reg [(4'hd):(1'h0)] reg1835 = (1'h0);
  reg [(4'hd):(1'h0)] reg1834 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire1833;
  wire signed [(4'ha):(1'h0)] wire1832;
  wire [(4'h9):(1'h0)] wire1831;
  wire signed [(3'h6):(1'h0)] wire1830;
  wire [(3'h5):(1'h0)] wire1829;
  wire [(4'hd):(1'h0)] wire1827;
  wire [(4'h9):(1'h0)] wire1766;
  wire signed [(5'h13):(1'h0)] wire1767;
  wire signed [(3'h4):(1'h0)] wire1768;
  reg [(2'h3):(1'h0)] reg1769 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1770 = (1'h0);
  reg [(4'he):(1'h0)] reg1771 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1772 = (1'h0);
  reg [(5'h11):(1'h0)] reg1773 = (1'h0);
  reg [(2'h3):(1'h0)] reg1774 = (1'h0);
  reg [(5'h14):(1'h0)] reg1775 = (1'h0);
  reg [(4'ha):(1'h0)] reg1776 = (1'h0);
  reg [(3'h5):(1'h0)] reg1777 = (1'h0);
  reg [(2'h2):(1'h0)] reg1778 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1779 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1780 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1781 = (1'h0);
  reg [(5'h12):(1'h0)] reg1782 = (1'h0);
  reg [(5'h15):(1'h0)] reg1783 = (1'h0);
  reg [(3'h6):(1'h0)] reg1784 = (1'h0);
  reg [(5'h13):(1'h0)] reg1785 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1786 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1787 = (1'h0);
  reg [(5'h14):(1'h0)] reg1788 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1789 = (1'h0);
  reg [(3'h7):(1'h0)] reg1790 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1791 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire1813;
  assign y = {wire1875,
                 wire1874,
                 wire1873,
                 reg1872,
                 reg1871,
                 reg1870,
                 reg1869,
                 reg1868,
                 reg1867,
                 reg1866,
                 reg1865,
                 reg1864,
                 reg1863,
                 reg1862,
                 reg1861,
                 reg1860,
                 reg1859,
                 reg1858,
                 reg1857,
                 reg1856,
                 reg1855,
                 reg1854,
                 reg1853,
                 reg1852,
                 reg1851,
                 reg1850,
                 reg1849,
                 reg1848,
                 reg1847,
                 wire1846,
                 wire1845,
                 wire1844,
                 reg1843,
                 reg1842,
                 reg1841,
                 reg1840,
                 reg1839,
                 reg1838,
                 reg1837,
                 reg1836,
                 reg1835,
                 reg1834,
                 wire1833,
                 wire1832,
                 wire1831,
                 wire1830,
                 wire1829,
                 wire1827,
                 wire1766,
                 wire1767,
                 wire1768,
                 reg1769,
                 reg1770,
                 reg1771,
                 reg1772,
                 reg1773,
                 reg1774,
                 reg1775,
                 reg1776,
                 reg1777,
                 reg1778,
                 reg1779,
                 reg1780,
                 reg1781,
                 reg1782,
                 reg1783,
                 reg1784,
                 reg1785,
                 reg1786,
                 reg1787,
                 reg1788,
                 reg1789,
                 reg1790,
                 reg1791,
                 wire1813,
                 (1'h0)};
  assign wire1766 = (wire1765 ?
                        (wire1764[(3'h7):(2'h2)] | (((8'hb9) * wire1763[(4'hc):(1'h0)]) <= wire1765)) : wire1762);
  assign wire1767 = (($signed(wire1766[(3'h5):(1'h1)]) ?
                        (wire1763[(3'h4):(1'h1)] ^ wire1763) : (&wire1763)) - ({{(wire1761 ?
                                wire1766 : wire1764),
                            (|wire1766)},
                        (~^$signed(wire1764))} <<< (^wire1763)));
  assign wire1768 = wire1761;
  always
    @(posedge clk) begin
      reg1769 <= (wire1766 > {wire1763[(3'h7):(3'h7)]});
      if ($unsigned(({reg1769[(2'h2):(2'h2)]} ?
          wire1761[(2'h2):(1'h1)] : (-({wire1768} ?
              (&reg1769) : (+wire1764))))))
        begin
          reg1770 <= ({(&$signed(wire1764)),
              ($signed(wire1764[(3'h5):(2'h3)]) >>> $signed((~(8'ha3))))} != wire1763[(4'h9):(1'h1)]);
          reg1771 <= $unsigned(wire1768);
          if ($unsigned((&{(8'ha5)})))
            begin
              reg1772 <= $signed($signed($signed(((wire1761 && wire1762) ?
                  (wire1766 ? wire1763 : wire1762) : (+wire1767)))));
              reg1773 <= wire1768[(2'h2):(1'h0)];
              reg1774 <= $unsigned(((reg1772[(1'h0):(1'h0)] ?
                  wire1768 : (8'hb2)) == reg1769[(2'h3):(1'h0)]));
              reg1775 <= $unsigned((~^$unsigned((reg1769 ?
                  reg1769[(2'h2):(1'h0)] : wire1761[(3'h4):(1'h1)]))));
              reg1776 <= $unsigned(wire1763);
            end
          else
            begin
              reg1772 <= $unsigned(($unsigned(wire1763[(4'hc):(1'h1)]) ?
                  wire1765 : $unsigned(((wire1763 ? wire1761 : reg1773) ?
                      reg1775 : $signed(wire1762)))));
            end
          reg1777 <= (($signed(wire1767) - (({reg1774} ?
                  $unsigned((8'haa)) : reg1775[(2'h2):(2'h2)]) < {wire1761})) ?
              (^$signed((((7'h43) ?
                  reg1769 : reg1774) > $unsigned(reg1771)))) : ((~&(8'haa)) ?
                  reg1771[(3'h5):(3'h5)] : (+$unsigned((wire1768 ^~ reg1776)))));
          reg1778 <= (~&(-(((reg1773 >= reg1774) << (wire1763 > reg1769)) | $signed((^~wire1765)))));
        end
      else
        begin
          reg1770 <= reg1775;
          reg1771 <= $signed({wire1765[(2'h3):(1'h1)]});
          reg1772 <= $unsigned((&((~^(wire1767 ? wire1766 : wire1765)) ?
              wire1762[(4'hb):(3'h5)] : (reg1769[(1'h0):(1'h0)] ^ (reg1776 & reg1771)))));
          reg1773 <= reg1777[(2'h3):(1'h0)];
        end
      if ((8'h9f))
        begin
          if ((wire1763 ? reg1774 : reg1774))
            begin
              reg1779 <= ((reg1775[(4'hc):(2'h3)] ?
                      (($unsigned(reg1770) + $signed(reg1774)) ?
                          $signed($unsigned((7'h41))) : wire1766) : (reg1775[(5'h14):(5'h11)] << ((!reg1777) != (!wire1761)))) ?
                  reg1778[(1'h1):(1'h0)] : wire1766[(3'h7):(1'h1)]);
            end
          else
            begin
              reg1779 <= $unsigned(($signed(((|reg1773) ?
                  {reg1773,
                      reg1770} : $signed(reg1771))) != $signed(reg1776[(3'h6):(2'h2)])));
              reg1780 <= $unsigned(((~(7'h41)) ?
                  $signed($signed((wire1764 + wire1762))) : $unsigned(reg1769)));
              reg1781 <= (^~$signed((~wire1767)));
              reg1782 <= $signed($unsigned(($signed(reg1777[(1'h0):(1'h0)]) <<< wire1761)));
              reg1783 <= reg1773[(3'h4):(1'h0)];
            end
          reg1784 <= (+(~^$unsigned($unsigned(wire1763))));
          reg1785 <= $signed(reg1777);
          reg1786 <= (8'hb1);
          reg1787 <= wire1762;
        end
      else
        begin
          reg1779 <= (((~$unsigned((~|reg1773))) ?
              (-($unsigned((8'ha1)) ? (~&reg1785) : reg1779)) : (!((~^(8'ha9)) ?
                  (reg1785 ?
                      reg1785 : reg1780) : reg1777))) >> (reg1769[(1'h0):(1'h0)] ?
              (+wire1767[(4'hb):(1'h0)]) : reg1783));
          reg1780 <= $signed(reg1779[(4'h8):(3'h7)]);
          reg1781 <= $unsigned(reg1778[(2'h2):(2'h2)]);
          reg1782 <= ((wire1765 <<< reg1778) ?
              reg1785[(4'hd):(2'h3)] : ((~|((reg1785 ? reg1772 : reg1787) ?
                      $unsigned(reg1785) : {reg1777})) ?
                  reg1773[(3'h7):(2'h2)] : $unsigned(wire1762)));
        end
      if ($signed($unsigned((&$signed($signed(reg1771))))))
        begin
          if (($unsigned((~$unsigned($signed(wire1767)))) ?
              {reg1773[(3'h6):(3'h6)],
                  {{{(8'hbd)}, (^wire1762)},
                      $unsigned((+reg1783))}} : ($unsigned(reg1771) ?
                  (+reg1784[(3'h5):(2'h3)]) : {(-wire1761),
                      (-$unsigned(wire1767))})))
            begin
              reg1788 <= reg1783[(2'h2):(1'h1)];
              reg1789 <= $signed(($unsigned(((~^reg1771) >> reg1774)) >>> (8'ha1)));
            end
          else
            begin
              reg1788 <= (reg1773 ?
                  ((~|reg1779[(3'h5):(3'h4)]) ?
                      reg1787[(4'he):(1'h1)] : (wire1763[(3'h7):(3'h6)] <<< $signed((reg1771 ?
                          reg1781 : (8'ha8))))) : reg1783);
              reg1789 <= {(8'ha7), wire1761};
              reg1790 <= $unsigned($unsigned((($signed(wire1765) || (|wire1764)) ~^ $signed(reg1776[(3'h4):(2'h3)]))));
            end
        end
      else
        begin
          if ({((8'ha2) ?
                  ((-(reg1783 <<< reg1787)) * (reg1773 - $unsigned(reg1786))) : {((wire1761 < wire1763) != reg1782)}),
              (reg1773 | wire1768[(2'h3):(2'h3)])})
            begin
              reg1788 <= $signed((reg1773 * (~&{(reg1773 ? wire1763 : reg1783),
                  $unsigned((8'hb7))})));
              reg1789 <= (|reg1776);
              reg1790 <= $unsigned((^~wire1766));
              reg1791 <= $signed($signed($unsigned((reg1772 > ((8'ha9) != wire1768)))));
            end
          else
            begin
              reg1788 <= wire1762[(2'h3):(1'h0)];
              reg1789 <= (reg1770[(4'h9):(3'h7)] <= wire1767);
              reg1790 <= (8'hb0);
              reg1791 <= ($signed((|(~reg1775))) < ($unsigned($unsigned($signed((8'hb1)))) | $unsigned(reg1770[(2'h2):(1'h0)])));
            end
        end
    end
  module1792 modinst1814 (wire1813, clk, reg1788, reg1786, reg1776, wire1762, wire1767);
  module1815 modinst1828 (wire1827, clk, reg1780, wire1762, reg1782, wire1765);
  assign wire1829 = $signed($signed((reg1778[(2'h2):(1'h1)] ?
                        ((^~wire1762) ? (!reg1776) : wire1767) : {(~|reg1788),
                            (reg1790 ? wire1762 : wire1768)})));
  assign wire1830 = (~|$signed(((+$signed(reg1786)) ~^ $unsigned((reg1783 ?
                        (8'ha3) : (7'h41))))));
  assign wire1831 = $unsigned(wire1813[(1'h0):(1'h0)]);
  assign wire1832 = (^~reg1774[(1'h1):(1'h1)]);
  assign wire1833 = {(~&$unsigned((~&$signed(reg1773)))),
                        reg1772[(3'h6):(3'h6)]};
  always
    @(posedge clk) begin
      if (wire1813[(2'h3):(2'h3)])
        begin
          if ($unsigned($signed($signed(((wire1832 < (8'ha5)) ?
              $signed((8'hb2)) : (8'ha4))))))
            begin
              reg1834 <= reg1771;
              reg1835 <= reg1834[(4'ha):(4'h8)];
            end
          else
            begin
              reg1834 <= (|$unsigned(($signed(reg1777) != ((wire1763 <= (8'hb3)) <<< ((8'hbc) ?
                  reg1784 : reg1784)))));
              reg1835 <= reg1777[(2'h3):(2'h2)];
              reg1836 <= (~&reg1782[(3'h7):(3'h7)]);
            end
        end
      else
        begin
          reg1834 <= $signed(reg1769[(2'h2):(2'h2)]);
        end
      reg1837 <= wire1768[(1'h0):(1'h0)];
      if ({$signed((|{(8'hab), wire1764}))})
        begin
          reg1838 <= reg1769[(2'h3):(2'h3)];
          reg1839 <= ((reg1783 << reg1834) ?
              (~&$unsigned(((~|reg1782) ?
                  wire1763[(4'hb):(4'hb)] : (reg1777 << (8'ha6))))) : $signed($signed(($unsigned((8'hab)) + (!reg1770)))));
        end
      else
        begin
          if ($unsigned(($signed($signed(reg1790[(2'h3):(2'h2)])) && $unsigned((+(reg1781 ?
              reg1776 : (8'hb1)))))))
            begin
              reg1838 <= $signed(wire1765);
              reg1839 <= ($signed(reg1787[(4'h9):(1'h0)]) ?
                  $unsigned($unsigned(wire1764[(4'hd):(3'h6)])) : (8'hae));
              reg1840 <= (^{(8'hb9)});
              reg1841 <= $signed((~^wire1830));
              reg1842 <= $signed($unsigned((|(reg1791[(3'h5):(1'h1)] ?
                  wire1762 : ((8'had) * (8'ha0))))));
            end
          else
            begin
              reg1838 <= (-(-$signed($signed($unsigned((8'hb7))))));
            end
        end
      reg1843 <= ({(~^$unsigned($signed(reg1783))),
              ({$unsigned(reg1780),
                  wire1767[(5'h12):(4'he)]} >> reg1780[(5'h14):(4'he)])} ?
          reg1834[(4'h8):(3'h4)] : ({((wire1764 ? wire1765 : (8'ha7)) ?
                      {(8'h9e)} : $unsigned(reg1787))} ?
              reg1774 : {(~^wire1829[(2'h2):(2'h2)])}));
    end
  assign wire1844 = $unsigned(((^~{((8'hae) ? reg1841 : wire1813),
                            $unsigned(wire1827)}) ?
                        (reg1835 >>> (~&(reg1789 ?
                            (8'hb5) : (8'ha6)))) : (reg1836[(2'h3):(1'h1)] ?
                            $signed(wire1761) : reg1786[(4'he):(2'h2)])));
  assign wire1845 = $unsigned(($signed({{reg1837}, (~reg1842)}) ?
                        {((wire1761 | wire1764) ?
                                {reg1780, wire1827} : (reg1790 ?
                                    reg1789 : reg1786)),
                            $unsigned($unsigned(reg1780))} : (~|((wire1813 ?
                                wire1764 : (8'ha3)) ?
                            (wire1761 ~^ (8'haf)) : reg1785[(3'h5):(2'h3)]))));
  assign wire1846 = (^$unsigned({$unsigned(wire1829[(2'h2):(2'h2)]), (8'hbe)}));
  always
    @(posedge clk) begin
      reg1847 <= (reg1843[(3'h6):(3'h5)] && $signed($signed((wire1761 ?
          wire1831 : (|reg1838)))));
      reg1848 <= $unsigned((~|((&$signed(reg1771)) || $unsigned((+wire1767)))));
    end
  always
    @(posedge clk) begin
      reg1849 <= {reg1780[(1'h1):(1'h0)], wire1830};
      reg1850 <= reg1838[(1'h1):(1'h1)];
      reg1851 <= (!((&wire1763[(4'he):(4'h8)]) ?
          reg1779[(2'h2):(1'h0)] : $unsigned((&(^~reg1786)))));
      reg1852 <= $signed(($signed(reg1840[(2'h2):(1'h0)]) ?
          ($unsigned((^reg1770)) ?
              (~^{(8'hab), reg1834}) : {reg1836}) : (reg1769 ?
              ($signed(reg1784) ?
                  (wire1845 != reg1785) : (!(8'ha0))) : ((wire1833 << reg1835) && (!reg1776)))));
      if ($unsigned({((reg1770 > (reg1781 ?
              reg1785 : (8'h9f))) >>> (^~$signed(reg1839))),
          (((wire1830 || (8'ha0)) ? (|wire1831) : wire1844) ?
              (wire1845[(4'hb):(4'ha)] >>> ((8'ha5) ?
                  reg1772 : reg1788)) : $unsigned(reg1791[(3'h5):(1'h0)]))}))
        begin
          reg1853 <= (((7'h40) >= (((reg1850 ? reg1774 : reg1848) ?
              (+reg1791) : $signed((7'h44))) || {(reg1849 ^~ reg1841),
              $unsigned(reg1784)})) && ((($signed(wire1830) ?
                  (reg1780 ?
                      reg1780 : wire1845) : (~^reg1790)) >> (^~(wire1829 > reg1770))) ?
              wire1767[(2'h3):(1'h1)] : reg1842));
          if ((&(reg1786 ? (~(~|wire1813)) : (~&(+reg1839)))))
            begin
              reg1854 <= reg1770[(4'hc):(2'h2)];
              reg1855 <= reg1771[(3'h4):(1'h0)];
            end
          else
            begin
              reg1854 <= (&($signed((&(reg1849 || reg1781))) || (+({reg1771} ?
                  $signed((8'hbd)) : ((7'h40) && reg1835)))));
              reg1855 <= $unsigned($signed(reg1849[(2'h3):(1'h1)]));
            end
          reg1856 <= reg1785;
          reg1857 <= (7'h40);
          if ({(7'h41),
              $signed((reg1778[(1'h1):(1'h0)] ?
                  (+wire1833) : $unsigned(wire1830[(3'h6):(1'h0)])))})
            begin
              reg1858 <= $signed(({wire1768[(2'h3):(2'h2)]} ?
                  reg1838 : ((reg1851[(1'h1):(1'h1)] >>> $unsigned(wire1764)) >> $unsigned((reg1785 && reg1790)))));
              reg1859 <= {$signed((&$unsigned(wire1767[(4'ha):(3'h5)]))),
                  reg1791[(5'h11):(2'h3)]};
              reg1860 <= (wire1845[(2'h3):(2'h3)] ?
                  reg1786[(4'hf):(3'h6)] : reg1777[(3'h4):(1'h0)]);
              reg1861 <= reg1836;
            end
          else
            begin
              reg1858 <= ($unsigned(reg1790[(2'h3):(1'h1)]) ?
                  $unsigned(reg1779[(2'h3):(2'h3)]) : wire1764[(5'h11):(4'hd)]);
              reg1859 <= $unsigned({reg1842[(4'hf):(4'hf)],
                  ($signed(reg1788) ?
                      $signed($signed(wire1832)) : $unsigned((reg1785 ^ (8'hae))))});
              reg1860 <= $unsigned((-{reg1776}));
              reg1861 <= {(wire1830 ~^ (&$signed((reg1837 ?
                      reg1784 : (8'ha2)))))};
              reg1862 <= (8'ha7);
            end
        end
      else
        begin
          if (($signed($signed(reg1775)) ~^ reg1840[(1'h1):(1'h0)]))
            begin
              reg1853 <= $signed(($unsigned($unsigned((reg1839 ?
                      wire1762 : (8'hbb)))) ?
                  (reg1777[(1'h0):(1'h0)] ?
                      $unsigned(wire1765[(2'h2):(1'h0)]) : reg1776) : (~&reg1780)));
              reg1854 <= reg1849[(4'he):(4'h9)];
              reg1855 <= ($signed((&wire1762[(5'h10):(3'h7)])) ?
                  (^$unsigned(reg1770[(4'h8):(4'h8)])) : ((reg1835[(3'h5):(2'h2)] ?
                      reg1837[(2'h3):(1'h1)] : $unsigned($signed(reg1850))) >>> {({(8'ha3),
                          reg1860} & $unsigned((8'ha1)))}));
            end
          else
            begin
              reg1853 <= (reg1776 || (~^(reg1853 << $unsigned($signed(reg1854)))));
              reg1854 <= wire1763[(3'h7):(2'h3)];
              reg1855 <= $unsigned($signed(reg1834[(4'h9):(3'h4)]));
              reg1856 <= {reg1836[(1'h1):(1'h1)], (8'hac)};
              reg1857 <= (reg1840 != ((((^reg1782) != (reg1853 ?
                      reg1858 : reg1842)) ?
                  {(+reg1782), $signed(reg1851)} : ($unsigned(reg1855) ?
                      reg1835[(3'h4):(1'h0)] : (|reg1782))) ~^ ({((8'ha9) ?
                          (8'hb1) : (8'ha6)),
                      (reg1780 ? wire1844 : (8'ha5))} ?
                  (~^(~(8'ha3))) : (~&$unsigned(wire1831)))));
            end
          if ((($unsigned((wire1833[(4'hd):(3'h7)] != $unsigned(wire1765))) ?
                  $signed($signed(reg1770[(4'ha):(2'h2)])) : reg1861) ?
              ($signed($unsigned((reg1840 == wire1845))) < ($unsigned(wire1844) ?
                  ($unsigned(reg1848) ?
                      reg1782 : (wire1768 >>> reg1835)) : {((8'hb2) ?
                          wire1762 : (8'hb0))})) : (wire1833 != (~|$unsigned($signed(reg1854))))))
            begin
              reg1858 <= ((^((-{reg1787}) <= (!$unsigned(wire1831)))) ?
                  $unsigned(reg1784[(3'h6):(2'h3)]) : $signed($unsigned(reg1840[(2'h2):(2'h2)])));
              reg1859 <= (((^~(~reg1785[(4'h9):(4'h9)])) ?
                  reg1862 : $unsigned(wire1844)) || $unsigned($signed(reg1837[(1'h0):(1'h0)])));
              reg1860 <= (~^(-reg1854));
            end
          else
            begin
              reg1858 <= $signed(reg1843);
            end
          reg1861 <= {wire1846};
          if ($signed({{reg1860}}))
            begin
              reg1862 <= ($unsigned(($signed((~&reg1860)) == $unsigned($unsigned((8'hb1))))) ~^ ((8'ha1) | wire1845[(4'h8):(3'h4)]));
            end
          else
            begin
              reg1862 <= $signed((((&(reg1851 != (7'h40))) ?
                  (8'ha8) : wire1827[(3'h5):(2'h2)]) <<< (&(^$unsigned(reg1782)))));
              reg1863 <= $unsigned((reg1791[(2'h3):(2'h2)] ^ $signed($unsigned($unsigned(reg1781)))));
              reg1864 <= (~^$signed(reg1836));
              reg1865 <= $signed($unsigned({{$unsigned(reg1791)},
                  (reg1851[(2'h3):(2'h3)] + reg1776)}));
            end
        end
    end
  always
    @(posedge clk) begin
      if ((-(!reg1835[(1'h0):(1'h0)])))
        begin
          reg1866 <= $unsigned($signed(reg1842));
          if ($signed($signed(($unsigned($signed(reg1837)) ?
              wire1844[(1'h0):(1'h0)] : ($signed(reg1834) ?
                  $signed(reg1840) : (|reg1851))))))
            begin
              reg1867 <= reg1784;
              reg1868 <= $unsigned(($signed(($signed(reg1854) | ((8'ha9) ?
                  wire1844 : reg1851))) > reg1863[(4'hd):(4'ha)]));
              reg1869 <= $signed({$signed(({(8'hb3)} ?
                      reg1861 : (wire1767 <<< reg1848)))});
              reg1870 <= (wire1761[(3'h7):(3'h5)] ?
                  (~^(wire1763[(4'hf):(3'h4)] ~^ ((|wire1762) ?
                      ((8'hb6) * reg1851) : $unsigned(reg1838)))) : ((^~$signed($unsigned(reg1780))) ?
                      reg1780 : reg1849[(3'h5):(2'h3)]));
            end
          else
            begin
              reg1867 <= ((-($signed(((8'hbf) ?
                  reg1854 : reg1770)) * reg1784[(3'h5):(3'h4)])) ^ reg1787);
              reg1868 <= (reg1855 ? (8'hbc) : wire1764);
              reg1869 <= (reg1772[(3'h6):(3'h4)] * (reg1849[(5'h12):(3'h5)] >= $unsigned((reg1854[(1'h0):(1'h0)] ?
                  (-reg1870) : {(8'hb4), (8'hab)}))));
            end
        end
      else
        begin
          if ($signed({(reg1839[(1'h0):(1'h0)] ~^ wire1765[(4'hf):(4'h8)])}))
            begin
              reg1866 <= $signed((wire1765 ?
                  $signed(reg1849[(4'h9):(1'h1)]) : (-reg1837[(2'h3):(2'h2)])));
              reg1867 <= $signed((!$unsigned((~$unsigned((8'h9f))))));
              reg1868 <= reg1850[(1'h1):(1'h1)];
              reg1869 <= wire1765[(3'h6):(3'h5)];
            end
          else
            begin
              reg1866 <= (^~$signed(reg1850[(4'h9):(2'h2)]));
              reg1867 <= $unsigned(($unsigned($unsigned(wire1833)) ?
                  (&reg1867) : $unsigned((!wire1829[(2'h2):(1'h1)]))));
              reg1868 <= (!reg1785);
              reg1869 <= reg1777;
            end
          reg1870 <= $signed($unsigned($unsigned(((8'ha2) ?
              wire1830 : {reg1840}))));
          reg1871 <= (reg1773 <= {wire1767[(4'hc):(3'h7)]});
          reg1872 <= $unsigned(reg1788);
        end
    end
  assign wire1873 = ($signed(($unsigned(reg1771) >>> wire1833[(2'h3):(2'h3)])) ^ (($signed(reg1852[(2'h3):(1'h0)]) && (+{reg1872})) ?
                        ((~(^reg1853)) ?
                            reg1772[(4'hf):(4'ha)] : (reg1870 ?
                                (reg1838 << (7'h43)) : reg1854[(1'h0):(1'h0)])) : reg1775[(3'h7):(2'h3)]));
  assign wire1874 = $signed((~&$signed(((~reg1834) != {(8'ha0)}))));
  assign wire1875 = ((({(&reg1858), {reg1866, wire1762}} ?
                            (^~{reg1867,
                                reg1849}) : $unsigned((~|reg1840))) + wire1830[(3'h5):(2'h3)]) ?
                        {{$unsigned((~&reg1836))},
                            (&(8'hbc))} : ((reg1835[(4'h8):(1'h1)] << reg1835[(4'hd):(3'h5)]) - $signed(reg1853[(3'h7):(2'h2)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1567
#( parameter param1756 = (((|{((8'hb7) ^~ (7'h41)), ((7'h40) || (8'hba))}) ? ((-((8'h9c) ? (8'hb7) : (8'had))) > (~|{(7'h42), (8'ha3)})) : ((!(-(8'hba))) ? {((8'h9d) & (8'hb4))} : (((7'h40) || (7'h44)) ? ((8'hb4) != (8'ha9)) : ((7'h42) ? (8'hab) : (8'ha5))))) ? ((((&(8'ha2)) ^ (~^(8'hae))) ? (((8'had) - (7'h40)) ? ((8'ha5) ^ (8'ha9)) : ((7'h44) ? (8'hae) : (8'ha5))) : (^((8'hb8) ~^ (8'ha6)))) ? {(((8'hac) ? (8'hbf) : (8'hbd)) ? ((8'hb7) ? (8'ha5) : (8'hac)) : {(8'ha3), (8'ha8)}), {((8'h9d) ? (8'hb1) : (8'hbe)), (8'ha9)}} : ({((8'ha4) - (8'ha3))} ? ({(8'ha3)} ? (~|(8'ha9)) : ((8'had) == (8'hab))) : (((8'ha5) ? (8'h9e) : (8'ha3)) & (-(8'ha8))))) : (((((8'ha5) ? (8'h9f) : (8'haa)) >> ((8'ha7) ? (8'hac) : (8'hb1))) ? (((8'ha7) ? (8'ha4) : (8'haf)) ? ((7'h42) ? (8'hb5) : (8'hb7)) : ((8'had) << (7'h42))) : (((8'ha8) ~^ (8'ha6)) ^ (+(8'hb2)))) > ((~|(!(8'hb3))) ? (^~{(8'haa)}) : (((8'hb7) ? (8'hae) : (8'ha3)) ? ((8'hb5) >= (8'hbf)) : ((8'hb0) <<< (8'haf)))))) )
(y, clk, wire1568, wire1569, wire1570, wire1571, wire1572);
  output wire [(32'h211):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire1568;
  input wire signed [(4'hd):(1'h0)] wire1569;
  input wire signed [(5'h14):(1'h0)] wire1570;
  input wire signed [(5'h11):(1'h0)] wire1571;
  input wire [(5'h15):(1'h0)] wire1572;
  wire signed [(4'h8):(1'h0)] wire1755;
  wire signed [(2'h2):(1'h0)] wire1754;
  wire [(5'h14):(1'h0)] wire1753;
  wire signed [(2'h3):(1'h0)] wire1752;
  wire [(3'h7):(1'h0)] wire1750;
  reg [(4'h8):(1'h0)] reg1725 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1724 = (1'h0);
  reg [(3'h7):(1'h0)] reg1723 = (1'h0);
  reg [(4'hb):(1'h0)] reg1722 = (1'h0);
  reg [(4'ha):(1'h0)] reg1721 = (1'h0);
  reg [(4'he):(1'h0)] reg1720 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1719 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1718 = (1'h0);
  reg [(3'h6):(1'h0)] reg1717 = (1'h0);
  reg [(5'h11):(1'h0)] reg1716 = (1'h0);
  reg [(4'ha):(1'h0)] reg1715 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire1673;
  wire signed [(4'hf):(1'h0)] wire1600;
  wire signed [(4'hf):(1'h0)] wire1599;
  wire signed [(4'hd):(1'h0)] wire1598;
  wire signed [(4'he):(1'h0)] wire1597;
  wire [(4'hf):(1'h0)] wire1596;
  wire signed [(4'ha):(1'h0)] wire1595;
  wire signed [(3'h4):(1'h0)] wire1594;
  wire [(5'h11):(1'h0)] wire1593;
  wire signed [(4'hf):(1'h0)] wire1592;
  wire signed [(5'h14):(1'h0)] wire1591;
  wire signed [(4'hd):(1'h0)] wire1589;
  reg [(5'h13):(1'h0)] reg1675 = (1'h0);
  reg [(5'h13):(1'h0)] reg1676 = (1'h0);
  reg [(5'h11):(1'h0)] reg1677 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1678 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1679 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1680 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1681 = (1'h0);
  reg [(3'h6):(1'h0)] reg1682 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1683 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1684 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1685 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1686 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire1713;
  assign y = {wire1755,
                 wire1754,
                 wire1753,
                 wire1752,
                 wire1750,
                 reg1725,
                 reg1724,
                 reg1723,
                 reg1722,
                 reg1721,
                 reg1720,
                 reg1719,
                 reg1718,
                 reg1717,
                 reg1716,
                 reg1715,
                 wire1673,
                 wire1600,
                 wire1599,
                 wire1598,
                 wire1597,
                 wire1596,
                 wire1595,
                 wire1594,
                 wire1593,
                 wire1592,
                 wire1591,
                 wire1589,
                 reg1675,
                 reg1676,
                 reg1677,
                 reg1678,
                 reg1679,
                 reg1680,
                 reg1681,
                 reg1682,
                 reg1683,
                 reg1684,
                 reg1685,
                 reg1686,
                 wire1713,
                 (1'h0)};
  module1573 modinst1590 (.wire1578(wire1569), .wire1574(wire1568), .wire1576(wire1570), .wire1577(wire1572), .y(wire1589), .clk(clk), .wire1575(wire1571));
  assign wire1591 = $signed(wire1572[(4'h8):(2'h3)]);
  assign wire1592 = ({$unsigned(wire1570[(4'h8):(4'h8)]),
                        ($signed((wire1589 ? wire1571 : wire1572)) ?
                            {(8'hb0)} : $signed($unsigned(wire1570)))} ^~ ((wire1572 == {$signed(wire1571),
                            ((7'h43) ? wire1570 : wire1572)}) ?
                        $unsigned(((wire1571 ?
                            wire1571 : (8'ha1)) > wire1591)) : wire1572[(4'ha):(1'h1)]));
  assign wire1593 = $unsigned($unsigned((8'ha6)));
  assign wire1594 = wire1571;
  assign wire1595 = $unsigned({wire1569[(4'hb):(2'h3)],
                        wire1593[(4'h9):(4'h8)]});
  assign wire1596 = $signed($unsigned($unsigned($unsigned((wire1591 ?
                        wire1570 : wire1571)))));
  assign wire1597 = (+(wire1596 ^~ (!$unsigned(wire1569[(4'hc):(4'h8)]))));
  assign wire1598 = wire1592[(1'h1):(1'h1)];
  assign wire1599 = (wire1595 || ((wire1592[(2'h3):(2'h3)] ?
                            (wire1589 ?
                                (~(8'hac)) : $signed(wire1571)) : $unsigned(((8'had) ?
                                wire1595 : wire1572))) ?
                        $signed(wire1597[(4'ha):(3'h7)]) : wire1569));
  assign wire1600 = $signed($signed((+$signed($unsigned(wire1596)))));
  module1601 modinst1674 (.wire1604(wire1589), .wire1602(wire1600), .y(wire1673), .wire1603(wire1592), .wire1606(wire1593), .clk(clk), .wire1605(wire1594));
  always
    @(posedge clk) begin
      reg1675 <= wire1600[(4'hf):(2'h2)];
      reg1676 <= $unsigned($signed($signed(wire1594)));
      if ($unsigned($unsigned($unsigned($signed($unsigned((8'hb6)))))))
        begin
          reg1677 <= (!$unsigned((wire1572[(5'h15):(2'h2)] ?
              ($signed((8'hb5)) ?
                  (~wire1594) : wire1569[(4'hb):(4'h8)]) : {wire1591})));
          reg1678 <= (8'hb5);
          reg1679 <= (wire1572[(3'h7):(2'h3)] >> (8'hb5));
          if (($unsigned({$unsigned(wire1593[(3'h6):(2'h2)]),
                  ((-wire1594) != reg1677[(5'h10):(4'he)])}) ?
              wire1597[(3'h5):(1'h1)] : {wire1597}))
            begin
              reg1680 <= wire1571[(3'h4):(3'h4)];
              reg1681 <= $unsigned(($signed($signed((7'h40))) ?
                  ((+$unsigned((8'hbf))) ?
                      $unsigned(wire1599[(4'hc):(4'hc)]) : (+(wire1598 ?
                          reg1680 : wire1589))) : (-$signed(reg1676))));
              reg1682 <= reg1677[(4'ha):(4'h9)];
            end
          else
            begin
              reg1680 <= $signed(((wire1589[(4'h8):(1'h1)] * wire1572[(2'h2):(1'h0)]) ?
                  $unsigned($signed(reg1682[(2'h3):(2'h2)])) : $unsigned((+(|wire1596)))));
              reg1681 <= wire1595[(4'ha):(1'h0)];
              reg1682 <= wire1597[(1'h0):(1'h0)];
              reg1683 <= (-$signed(($signed((+(8'ha5))) ^~ $unsigned($unsigned(reg1678)))));
              reg1684 <= (reg1677[(2'h2):(1'h0)] ?
                  {wire1572[(2'h2):(1'h0)], wire1599} : $unsigned((+wire1572)));
            end
          reg1685 <= $unsigned((~&reg1677));
        end
      else
        begin
          reg1677 <= ((8'hbc) >> $unsigned(reg1677[(3'h6):(3'h4)]));
          reg1678 <= $signed(($unsigned(reg1675[(2'h3):(2'h2)]) ?
              (8'hb1) : ((~&$unsigned(reg1677)) - $signed((wire1598 ?
                  (8'hb9) : reg1677)))));
        end
      reg1686 <= (~^{(+(~^(-wire1569)))});
    end
  module1687 modinst1714 (.wire1688(wire1589), .y(wire1713), .wire1691(reg1679), .clk(clk), .wire1690(reg1675), .wire1692(wire1673), .wire1689(reg1680));
  always
    @(posedge clk) begin
      if (reg1685)
        begin
          reg1715 <= $signed(wire1568[(4'he):(4'hd)]);
          if ((&(8'ha3)))
            begin
              reg1716 <= reg1685;
            end
          else
            begin
              reg1716 <= reg1679;
              reg1717 <= reg1686;
            end
          if (({reg1683[(2'h2):(1'h1)]} << reg1684[(2'h2):(1'h1)]))
            begin
              reg1718 <= (reg1682[(3'h4):(2'h3)] * {($signed((~&wire1572)) ?
                      $unsigned($unsigned(reg1685)) : (&wire1596))});
              reg1719 <= ({wire1597[(3'h6):(1'h1)]} >>> (({$unsigned(reg1716),
                  (|reg1683)} * (-(wire1572 << (8'h9f)))) << ((wire1594[(3'h4):(2'h2)] ?
                  reg1718 : $signed(reg1676)) | wire1572[(1'h1):(1'h0)])));
              reg1720 <= $unsigned((~|($unsigned({wire1591, wire1673}) ?
                  (8'ha2) : (~wire1596))));
              reg1721 <= ((reg1719[(2'h3):(1'h1)] ?
                      $signed({(wire1673 >> (8'ha0)),
                          $signed(reg1675)}) : (!$signed(((8'hab) ?
                          reg1680 : (8'ha2))))) ?
                  $unsigned({reg1718}) : wire1570);
            end
          else
            begin
              reg1718 <= $signed(reg1719[(3'h4):(2'h2)]);
              reg1719 <= wire1592[(2'h2):(2'h2)];
              reg1720 <= ($unsigned(($unsigned(reg1716) ?
                  $signed((^~wire1595)) : reg1682[(3'h5):(2'h3)])) != $signed(wire1596));
              reg1721 <= {$signed((!$signed(wire1713[(4'he):(3'h5)]))),
                  (~^wire1599[(1'h1):(1'h0)])};
              reg1722 <= reg1685[(3'h5):(1'h0)];
            end
          if ($signed((~|reg1675[(4'he):(1'h1)])))
            begin
              reg1723 <= $unsigned(wire1597);
            end
          else
            begin
              reg1723 <= reg1717[(2'h3):(2'h2)];
            end
        end
      else
        begin
          reg1715 <= ({$unsigned($signed($signed((8'hb1)))),
              $unsigned($signed({wire1599, reg1721}))} & ($signed((~(reg1716 ?
              reg1681 : wire1713))) != ({reg1685,
              (~^wire1589)} >>> wire1600[(1'h0):(1'h0)])));
          reg1716 <= $unsigned({(((reg1676 >= reg1684) <<< reg1723[(1'h1):(1'h0)]) ?
                  reg1715[(4'ha):(3'h7)] : {(wire1570 ^~ reg1683),
                      (reg1678 ? (7'h40) : reg1719)}),
              reg1683[(3'h4):(1'h0)]});
          if ($unsigned(wire1599))
            begin
              reg1717 <= (wire1571 ^~ reg1723);
              reg1718 <= $signed({(8'hb5),
                  (($unsigned(reg1684) ?
                          reg1715[(3'h4):(3'h4)] : (reg1678 ?
                              reg1719 : wire1593)) ?
                      ((+(8'hbd)) ?
                          reg1679[(3'h7):(1'h0)] : $unsigned((7'h41))) : (reg1719 ?
                          $signed(wire1571) : $signed(wire1673)))});
              reg1719 <= ($unsigned($signed((wire1599[(3'h7):(2'h2)] | (~|reg1715)))) + ((~&reg1679) << {wire1597}));
              reg1720 <= $signed(reg1676[(1'h0):(1'h0)]);
            end
          else
            begin
              reg1717 <= $unsigned(((reg1680 ?
                      {$signed(wire1568),
                          (reg1681 ? (8'hb6) : (8'hbd))} : ((&wire1592) ?
                          wire1597 : (~(8'haf)))) ?
                  ((7'h43) ^ reg1682[(3'h5):(2'h3)]) : (reg1679 > $signed((~^reg1716)))));
            end
        end
      reg1724 <= {(+reg1683), (-reg1681[(4'h8):(4'h8)])};
      reg1725 <= ((~&(((reg1717 ? reg1685 : reg1679) - (^~(8'hb8))) ?
          {$unsigned(reg1721)} : ({wire1589,
              (8'hb1)} + (wire1571 < reg1724)))) >> $signed(($signed($unsigned(wire1570)) <= reg1684)));
    end
  module1726 modinst1751 (wire1750, clk, reg1721, reg1718, reg1724, reg1720);
  assign wire1752 = ((reg1678 || reg1715) ?
                        $unsigned((~^(^~$unsigned(reg1725)))) : (8'haa));
  assign wire1753 = ((reg1719 & wire1572) ?
                        $signed(($signed($signed(reg1676)) ?
                            $unsigned((~^reg1678)) : (wire1596[(4'ha):(3'h5)] ?
                                wire1673 : ((8'hb1) ~^ reg1677)))) : $unsigned(wire1673));
  assign wire1754 = {$unsigned($unsigned((~|(|wire1569)))), $signed(reg1684)};
  assign wire1755 = (~^wire1597[(3'h5):(1'h0)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1435
#( parameter param1554 = ({({((7'h44) < (8'hb4))} ? ({(8'ha3)} >> ((8'hb4) ^~ (8'ha5))) : ((^(8'hba)) - (!(8'ha8)))), ((8'h9e) ? (!((8'hbc) ? (8'hb3) : (8'hb8))) : (((8'haa) > (8'hb1)) != ((8'ha4) ? (8'ha2) : (8'haa))))} < (~(^~{(!(8'ha4)), ((8'hb5) ? (7'h43) : (8'ha7))})))
, parameter param1555 = (param1554 - (&(param1554 - param1554))) )
(y, clk, wire1440, wire1439, wire1438, wire1437, wire1436);
  output wire [(32'h77):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire1440;
  input wire [(5'h14):(1'h0)] wire1439;
  input wire [(5'h10):(1'h0)] wire1438;
  input wire [(5'h12):(1'h0)] wire1437;
  input wire [(3'h7):(1'h0)] wire1436;
  wire [(4'hb):(1'h0)] wire1553;
  wire signed [(4'hb):(1'h0)] wire1551;
  wire [(4'h8):(1'h0)] wire1499;
  reg [(3'h6):(1'h0)] reg1498 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire1497;
  wire [(4'hd):(1'h0)] wire1496;
  wire [(3'h4):(1'h0)] wire1495;
  wire [(4'hc):(1'h0)] wire1493;
  reg signed [(4'hd):(1'h0)] reg1444 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1443 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire1442;
  wire [(4'h9):(1'h0)] wire1441;
  assign y = {wire1553,
                 wire1551,
                 wire1499,
                 reg1498,
                 wire1497,
                 wire1496,
                 wire1495,
                 wire1493,
                 reg1444,
                 reg1443,
                 wire1442,
                 wire1441,
                 (1'h0)};
  assign wire1441 = wire1439[(1'h0):(1'h0)];
  assign wire1442 = wire1436[(2'h3):(1'h1)];
  always
    @(posedge clk) begin
      reg1443 <= ($signed((7'h40)) == $signed($signed(wire1438)));
      reg1444 <= (~^(-wire1441[(1'h0):(1'h0)]));
    end
  module1445 modinst1494 (.wire1449(wire1441), .clk(clk), .wire1446(wire1438), .wire1448(wire1440), .wire1447(wire1436), .y(wire1493));
  assign wire1495 = (wire1442[(1'h1):(1'h1)] ?
                        $unsigned(wire1436) : $unsigned($unsigned(wire1439[(3'h4):(1'h0)])));
  assign wire1496 = $signed($signed($unsigned($signed((~^reg1443)))));
  assign wire1497 = ($signed(wire1438[(4'hc):(4'h8)]) ?
                        $signed($signed({(wire1440 ? reg1443 : wire1442),
                            (&wire1440)})) : $unsigned($signed(((8'hba) < $signed(wire1441)))));
  always
    @(posedge clk) begin
      reg1498 <= (!$signed($signed($unsigned(reg1443))));
    end
  assign wire1499 = ((~^$unsigned(($unsigned(wire1439) && (reg1498 <<< wire1442)))) >>> $unsigned((^~reg1498[(3'h4):(2'h2)])));
  module1500 modinst1552 (wire1551, clk, wire1493, wire1497, wire1439, wire1436);
  assign wire1553 = {reg1443, (^(^~{wire1493[(4'h8):(4'h8)]}))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1500
#( parameter param1549 = ((~^(~^{((8'ha1) && (8'hb6)), (~^(8'ha5))})) ? ((8'hbc) ^ (-(&(^(8'ha1))))) : (((((8'hb9) == (7'h42)) | ((8'ha0) ? (8'hb0) : (8'hbd))) ? ((~(7'h44)) * {(8'h9e)}) : ((~(7'h40)) ? ((7'h43) ? (8'hb6) : (8'haf)) : ((8'ha2) > (8'hae)))) <<< {{(|(8'h9e))}}))
, parameter param1550 = (param1549 >= param1549) )
(y, clk, wire1504, wire1503, wire1502, wire1501);
  output wire [(32'h1da):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire1504;
  input wire [(5'h15):(1'h0)] wire1503;
  input wire signed [(5'h14):(1'h0)] wire1502;
  input wire signed [(3'h5):(1'h0)] wire1501;
  wire signed [(4'hc):(1'h0)] wire1548;
  wire signed [(5'h11):(1'h0)] wire1547;
  wire [(5'h11):(1'h0)] wire1546;
  reg signed [(4'hb):(1'h0)] reg1545 = (1'h0);
  reg [(4'hb):(1'h0)] reg1544 = (1'h0);
  reg [(3'h7):(1'h0)] reg1543 = (1'h0);
  reg [(4'h8):(1'h0)] reg1542 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1541 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1540 = (1'h0);
  reg [(4'ha):(1'h0)] reg1539 = (1'h0);
  reg [(5'h14):(1'h0)] reg1538 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1537 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1536 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1535 = (1'h0);
  reg [(5'h10):(1'h0)] reg1534 = (1'h0);
  reg [(2'h3):(1'h0)] reg1533 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1532 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1531 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1530 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1529 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1528 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1527 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1526 = (1'h0);
  reg [(3'h4):(1'h0)] reg1525 = (1'h0);
  reg [(4'hb):(1'h0)] reg1524 = (1'h0);
  reg [(2'h2):(1'h0)] reg1523 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1522 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1521 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1520 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1519 = (1'h0);
  reg [(2'h2):(1'h0)] reg1518 = (1'h0);
  reg [(4'hc):(1'h0)] reg1517 = (1'h0);
  reg [(5'h14):(1'h0)] reg1516 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1515 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1514 = (1'h0);
  reg [(3'h6):(1'h0)] reg1513 = (1'h0);
  reg [(5'h10):(1'h0)] reg1512 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1511 = (1'h0);
  reg [(2'h3):(1'h0)] reg1510 = (1'h0);
  reg [(3'h5):(1'h0)] reg1509 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire1508;
  reg [(4'h8):(1'h0)] reg1507 = (1'h0);
  wire [(2'h3):(1'h0)] wire1506;
  wire [(2'h3):(1'h0)] wire1505;
  assign y = {wire1548,
                 wire1547,
                 wire1546,
                 reg1545,
                 reg1544,
                 reg1543,
                 reg1542,
                 reg1541,
                 reg1540,
                 reg1539,
                 reg1538,
                 reg1537,
                 reg1536,
                 reg1535,
                 reg1534,
                 reg1533,
                 reg1532,
                 reg1531,
                 reg1530,
                 reg1529,
                 reg1528,
                 reg1527,
                 reg1526,
                 reg1525,
                 reg1524,
                 reg1523,
                 reg1522,
                 reg1521,
                 reg1520,
                 reg1519,
                 reg1518,
                 reg1517,
                 reg1516,
                 reg1515,
                 reg1514,
                 reg1513,
                 reg1512,
                 reg1511,
                 reg1510,
                 reg1509,
                 wire1508,
                 reg1507,
                 wire1506,
                 wire1505,
                 (1'h0)};
  assign wire1505 = wire1503[(5'h15):(4'he)];
  assign wire1506 = (-wire1501[(3'h4):(1'h1)]);
  always
    @(posedge clk) begin
      reg1507 <= wire1504[(4'h8):(3'h6)];
    end
  assign wire1508 = $signed((((-{wire1505}) ?
                        ({wire1503, (8'hbf)} ?
                            $unsigned((7'h44)) : $signed(wire1504)) : wire1504[(2'h2):(1'h0)]) >> (8'h9d)));
  always
    @(posedge clk) begin
      reg1509 <= wire1508;
      if ((^(8'hac)))
        begin
          if ($unsigned((!((&(8'h9f)) || (((8'ha0) ?
              wire1501 : wire1508) & $unsigned(wire1504))))))
            begin
              reg1510 <= (~^$signed(((~^$unsigned(reg1509)) ?
                  (~$unsigned(wire1508)) : ((wire1506 ?
                      wire1505 : wire1504) <<< wire1505[(1'h1):(1'h1)]))));
              reg1511 <= (wire1501[(2'h3):(2'h3)] << reg1509[(3'h4):(1'h1)]);
            end
          else
            begin
              reg1510 <= wire1508[(3'h4):(1'h1)];
              reg1511 <= (wire1503 ? reg1510 : {wire1503});
              reg1512 <= wire1506;
              reg1513 <= (~^{(8'hb5),
                  (($signed((7'h44)) || (reg1507 ^~ (7'h40))) ?
                      ({(8'ha7)} | $unsigned(reg1510)) : ((wire1502 >>> reg1510) && reg1509))});
              reg1514 <= wire1504[(1'h0):(1'h0)];
            end
          if ($signed((wire1501[(1'h0):(1'h0)] ?
              (~{{(8'hac)}}) : ($unsigned((reg1512 ?
                  (8'hb8) : (8'hba))) || (^wire1505[(2'h3):(2'h2)])))))
            begin
              reg1515 <= (reg1511[(2'h2):(1'h1)] ?
                  {wire1503,
                      wire1506[(1'h0):(1'h0)]} : (~|(^$signed($signed(reg1513)))));
              reg1516 <= (wire1502[(4'h9):(1'h0)] >> (~^{(&reg1515),
                  reg1514[(2'h2):(1'h1)]}));
              reg1517 <= $unsigned(($signed(($signed(reg1515) + $unsigned(reg1514))) && (8'hb1)));
              reg1518 <= $unsigned($unsigned($signed($signed({reg1509}))));
              reg1519 <= $unsigned($unsigned(({(+wire1504),
                      reg1510[(1'h0):(1'h0)]} ?
                  $signed($signed(wire1501)) : (-{reg1514}))));
            end
          else
            begin
              reg1515 <= reg1509;
              reg1516 <= (~(wire1504[(2'h3):(2'h2)] ~^ ((!((7'h41) ?
                      reg1513 : (8'hbf))) ?
                  reg1507[(3'h5):(3'h4)] : $signed($unsigned(reg1512)))));
            end
          if (reg1515[(4'ha):(1'h1)])
            begin
              reg1520 <= $signed(reg1510);
              reg1521 <= ((^~(({reg1520} ?
                          $signed(wire1501) : $unsigned(reg1512)) ?
                      (wire1501[(1'h1):(1'h1)] ?
                          (!(8'hbc)) : {reg1507}) : $unsigned((reg1517 ?
                          reg1520 : wire1502)))) ?
                  (((wire1501 ?
                          $signed(reg1518) : (wire1508 & wire1506)) - reg1519[(2'h3):(2'h2)]) ?
                      $unsigned((8'hb9)) : (({reg1514, (7'h41)} ?
                          (reg1515 ?
                              reg1511 : wire1505) : reg1509) | (~&$signed(reg1509)))) : reg1516);
            end
          else
            begin
              reg1520 <= (($signed({reg1519,
                      $unsigned(wire1501)}) | wire1508[(5'h12):(5'h11)]) ?
                  (((|$unsigned(wire1504)) < (~|$unsigned(reg1510))) ?
                      (~&($unsigned(wire1502) ?
                          {wire1504, reg1521} : (reg1515 ?
                              reg1518 : reg1518))) : reg1511[(3'h4):(2'h3)]) : wire1502[(4'hf):(1'h1)]);
              reg1521 <= ($unsigned(wire1504[(2'h2):(1'h1)]) ?
                  (8'ha6) : {{reg1516[(4'hf):(2'h2)]},
                      $signed($unsigned(wire1501[(3'h4):(3'h4)]))});
              reg1522 <= reg1509;
              reg1523 <= ((($signed($signed(wire1505)) ?
                      $signed((8'hba)) : ((reg1509 ?
                          wire1504 : wire1503) > {reg1512})) ?
                  ((|(~^(8'hb3))) ?
                      $unsigned((-reg1512)) : {reg1512[(1'h0):(1'h0)],
                          reg1510}) : $signed($signed((reg1507 && wire1504)))) | $signed(wire1505));
              reg1524 <= wire1508;
            end
          reg1525 <= {reg1521[(2'h2):(1'h1)], ($unsigned(reg1515) ~^ (8'hbd))};
          reg1526 <= $signed(reg1517[(2'h2):(1'h1)]);
        end
      else
        begin
          reg1510 <= $signed(($signed((reg1510[(2'h3):(1'h0)] & $unsigned(reg1522))) << (((reg1521 != (8'hbb)) ?
              (reg1512 ? reg1522 : reg1517) : ((8'ha2) ?
                  reg1510 : (8'ha4))) ^ reg1514)));
          reg1511 <= $unsigned($unsigned($unsigned((reg1521[(1'h1):(1'h0)] ?
              (&reg1512) : (wire1505 <<< wire1504)))));
        end
    end
  always
    @(posedge clk) begin
      reg1527 <= $signed(reg1521[(1'h0):(1'h0)]);
      if (wire1504)
        begin
          reg1528 <= (!reg1516);
          reg1529 <= $unsigned(reg1511[(3'h5):(3'h5)]);
          if ((~$signed((wire1505[(1'h1):(1'h1)] ?
              reg1511[(2'h3):(2'h2)] : ((reg1520 * wire1505) ?
                  wire1502 : (reg1524 ? reg1518 : wire1503))))))
            begin
              reg1530 <= reg1510;
              reg1531 <= $unsigned($unsigned({{(reg1529 ? reg1525 : reg1517),
                      reg1516[(1'h1):(1'h0)]}}));
              reg1532 <= $signed($signed(((((8'haa) ?
                  wire1501 : wire1502) >>> {wire1502}) >= {wire1502})));
              reg1533 <= {$unsigned(reg1528[(2'h3):(1'h0)]),
                  $signed((reg1524 ?
                      {reg1512[(1'h0):(1'h0)]} : ($unsigned(reg1521) ~^ reg1523[(2'h2):(1'h0)])))};
              reg1534 <= (~(reg1521[(1'h1):(1'h0)] * ((-$signed(reg1522)) >> ((reg1509 ?
                      (8'hbc) : reg1512) ?
                  wire1502[(5'h14):(4'hb)] : (reg1519 - reg1517)))));
            end
          else
            begin
              reg1530 <= (((($signed(reg1510) < (!reg1532)) ?
                      $signed((wire1508 <= wire1508)) : $unsigned({reg1534})) ?
                  reg1523[(1'h0):(1'h0)] : (~|(wire1508[(3'h4):(1'h1)] ?
                      $unsigned((8'ha8)) : $signed(reg1520)))) ^ reg1517);
              reg1531 <= reg1520[(3'h5):(3'h4)];
              reg1532 <= ($unsigned(((+$unsigned(reg1532)) ~^ (|wire1508))) ?
                  {($signed(reg1514[(2'h3):(1'h0)]) ?
                          (-{reg1513, reg1523}) : (~&(~reg1510)))} : wire1508);
              reg1533 <= wire1508;
            end
        end
      else
        begin
          if (((^~($unsigned((reg1511 ?
                  reg1531 : reg1524)) || reg1510[(1'h1):(1'h0)])) ?
              (($signed(((8'hb8) ? reg1515 : reg1534)) ?
                      reg1511 : $signed(reg1516)) ?
                  $unsigned($signed({wire1501})) : $signed(((~reg1507) >>> (^~wire1502)))) : (reg1512 ?
                  (~$signed(reg1530)) : (reg1511[(1'h0):(1'h0)] ?
                      reg1517 : ((wire1504 ? reg1517 : reg1511) ?
                          reg1513 : wire1504[(3'h5):(2'h2)])))))
            begin
              reg1528 <= $signed($signed($signed({$signed(wire1504)})));
              reg1529 <= $signed(reg1523[(1'h0):(1'h0)]);
            end
          else
            begin
              reg1528 <= reg1530[(4'he):(2'h3)];
            end
          reg1530 <= reg1518;
          reg1531 <= wire1503[(4'he):(3'h4)];
          reg1532 <= reg1534[(2'h3):(1'h1)];
          reg1533 <= reg1522[(4'hc):(2'h3)];
        end
      reg1535 <= ($signed(wire1506) ?
          reg1522 : ((((8'hbb) < $signed(wire1501)) || $unsigned($signed(wire1501))) ?
              wire1501 : ($signed($signed(wire1506)) ?
                  wire1501 : reg1521[(2'h2):(1'h1)])));
    end
  always
    @(posedge clk) begin
      reg1536 <= ((~^reg1513) <= (-(($signed(reg1535) ?
          $unsigned(reg1511) : reg1518[(1'h0):(1'h0)]) >>> (reg1521[(2'h2):(1'h0)] ?
          $signed(reg1518) : $unsigned(reg1522)))));
      reg1537 <= (~&$unsigned((reg1523[(1'h0):(1'h0)] ?
          wire1508 : (reg1531 ^~ (reg1517 << reg1510)))));
      if (((~&$unsigned($unsigned(((8'hba) ? reg1514 : (8'ha0))))) ?
          reg1514 : wire1501[(2'h2):(1'h1)]))
        begin
          reg1538 <= $signed(reg1513);
          reg1539 <= ((($unsigned($unsigned(reg1523)) ^ reg1530[(5'h12):(4'he)]) >> (|$signed((reg1511 + wire1505)))) ~^ (8'hab));
          reg1540 <= (8'haa);
          if (wire1508[(1'h0):(1'h0)])
            begin
              reg1541 <= {reg1515,
                  $unsigned((|(reg1512 ^ (reg1533 ? reg1531 : wire1502))))};
              reg1542 <= ($signed($unsigned(((+(8'ha3)) ?
                      (reg1507 ? wire1503 : reg1539) : ((8'hab) ?
                          (8'had) : (8'hae))))) ?
                  ((reg1538 ?
                      $signed($signed(reg1533)) : (~&$signed(reg1531))) > ({{reg1517},
                          (8'hac)} ?
                      {(reg1518 | reg1521)} : reg1518[(2'h2):(2'h2)])) : $signed((((~reg1536) ?
                          wire1504[(3'h5):(2'h2)] : $signed((8'ha8))) ?
                      (~|(~&reg1520)) : {(~^reg1530), (8'hbd)})));
              reg1543 <= ($signed($signed($unsigned((reg1520 ?
                      reg1516 : wire1503)))) ?
                  reg1519[(2'h2):(1'h1)] : ((~wire1501) | (+((~^reg1519) <= reg1523))));
              reg1544 <= $signed((&wire1501[(1'h1):(1'h1)]));
            end
          else
            begin
              reg1541 <= reg1531[(3'h6):(3'h6)];
              reg1542 <= (8'hb3);
              reg1543 <= {$signed({(^~reg1533)}), reg1533[(1'h1):(1'h1)]};
              reg1544 <= (|(&(({(8'hb6)} >>> (|(8'haf))) | $signed(reg1518))));
            end
        end
      else
        begin
          reg1538 <= ($signed(((reg1526 ^ (reg1517 >> reg1510)) || $signed({reg1534,
                  reg1532}))) ?
              (8'hb3) : (($signed($unsigned(reg1538)) <<< reg1529[(5'h11):(4'h9)]) ?
                  $signed((~{reg1537, reg1534})) : ($unsigned((^~wire1501)) ?
                      ((^reg1543) ?
                          {reg1511,
                              (8'hb2)} : (wire1501 || reg1544)) : {((8'hb4) ?
                              (8'hbc) : reg1540)})));
          if ($unsigned(reg1538[(4'he):(1'h0)]))
            begin
              reg1539 <= reg1536[(4'hf):(3'h6)];
              reg1540 <= ((!$signed((8'hbd))) ?
                  reg1540[(4'h8):(3'h6)] : reg1522[(3'h7):(1'h1)]);
              reg1541 <= reg1514[(1'h1):(1'h1)];
              reg1542 <= ($unsigned((reg1523[(2'h2):(1'h0)] ?
                      reg1513[(1'h0):(1'h0)] : reg1517[(2'h2):(2'h2)])) ?
                  $signed($unsigned(reg1531)) : ($unsigned(((8'had) << $signed(reg1539))) + reg1544[(1'h1):(1'h0)]));
            end
          else
            begin
              reg1539 <= $unsigned(wire1508[(2'h3):(2'h2)]);
              reg1540 <= {((-$unsigned((^reg1532))) ?
                      ((|(reg1533 ? reg1536 : reg1511)) ?
                          ((+reg1521) <<< (reg1538 ?
                              reg1522 : reg1526)) : wire1503) : reg1519),
                  (7'h44)};
              reg1541 <= $unsigned($signed(wire1505));
              reg1542 <= reg1544;
            end
          reg1543 <= (^~reg1523);
          reg1544 <= reg1523[(2'h2):(2'h2)];
          reg1545 <= reg1532[(1'h0):(1'h0)];
        end
    end
  assign wire1546 = (reg1528[(1'h0):(1'h0)] & ({((-reg1526) << {reg1538}),
                        $unsigned($unsigned(reg1521))} >>> (~{wire1501})));
  assign wire1547 = reg1544;
  assign wire1548 = ((8'h9f) & wire1506[(1'h1):(1'h1)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1445  (y, clk, wire1449, wire1448, wire1447, wire1446);
  output wire [(32'h20f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire1449;
  input wire [(4'ha):(1'h0)] wire1448;
  input wire [(3'h7):(1'h0)] wire1447;
  input wire signed [(5'h10):(1'h0)] wire1446;
  wire [(3'h6):(1'h0)] wire1492;
  wire signed [(4'h8):(1'h0)] wire1491;
  wire [(4'h8):(1'h0)] wire1490;
  wire [(4'ha):(1'h0)] wire1489;
  wire signed [(5'h11):(1'h0)] wire1488;
  wire [(4'ha):(1'h0)] wire1487;
  wire signed [(5'h10):(1'h0)] wire1486;
  wire [(4'he):(1'h0)] wire1485;
  wire [(4'h8):(1'h0)] wire1484;
  wire [(4'h9):(1'h0)] wire1483;
  wire [(3'h6):(1'h0)] wire1482;
  wire [(5'h15):(1'h0)] wire1481;
  wire signed [(2'h2):(1'h0)] wire1480;
  reg [(3'h7):(1'h0)] reg1479 = (1'h0);
  reg [(3'h5):(1'h0)] reg1478 = (1'h0);
  reg [(5'h13):(1'h0)] reg1477 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1476 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1475 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1474 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1473 = (1'h0);
  reg [(4'ha):(1'h0)] reg1472 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1471 = (1'h0);
  wire [(5'h14):(1'h0)] wire1470;
  reg signed [(5'h13):(1'h0)] reg1469 = (1'h0);
  reg [(5'h15):(1'h0)] reg1468 = (1'h0);
  reg [(5'h15):(1'h0)] reg1467 = (1'h0);
  reg [(4'he):(1'h0)] reg1466 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1465 = (1'h0);
  reg [(5'h10):(1'h0)] reg1464 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1463 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1462 = (1'h0);
  wire [(5'h11):(1'h0)] wire1461;
  reg signed [(2'h3):(1'h0)] reg1460 = (1'h0);
  reg [(5'h12):(1'h0)] reg1459 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1458 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1457 = (1'h0);
  reg [(5'h15):(1'h0)] reg1456 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1455 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1454 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1453 = (1'h0);
  reg [(5'h12):(1'h0)] reg1452 = (1'h0);
  wire [(2'h2):(1'h0)] wire1451;
  reg [(5'h12):(1'h0)] reg1450 = (1'h0);
  assign y = {wire1492,
                 wire1491,
                 wire1490,
                 wire1489,
                 wire1488,
                 wire1487,
                 wire1486,
                 wire1485,
                 wire1484,
                 wire1483,
                 wire1482,
                 wire1481,
                 wire1480,
                 reg1479,
                 reg1478,
                 reg1477,
                 reg1476,
                 reg1475,
                 reg1474,
                 reg1473,
                 reg1472,
                 reg1471,
                 wire1470,
                 reg1469,
                 reg1468,
                 reg1467,
                 reg1466,
                 reg1465,
                 reg1464,
                 reg1463,
                 reg1462,
                 wire1461,
                 reg1460,
                 reg1459,
                 reg1458,
                 reg1457,
                 reg1456,
                 reg1455,
                 reg1454,
                 reg1453,
                 reg1452,
                 wire1451,
                 reg1450,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1450 <= (^({($signed((8'hb9)) >= (wire1448 ? wire1447 : wire1447)),
              wire1446} ?
          $unsigned(((8'hab) != wire1446[(4'he):(4'h9)])) : (($unsigned((8'hb2)) ?
                  $signed(wire1448) : (^~wire1446)) ?
              {(~&(8'haa)), (|wire1447)} : (|{wire1448, wire1449}))));
    end
  assign wire1451 = wire1449[(3'h6):(2'h3)];
  always
    @(posedge clk) begin
      if ($unsigned((wire1447 == (wire1446 ?
          $unsigned(wire1446) : $signed($signed(wire1448))))))
        begin
          if (($signed(reg1450) ^ (wire1447[(3'h7):(3'h6)] ?
              {$signed((reg1450 ? wire1446 : wire1449)),
                  (wire1448 ?
                      (reg1450 ^~ (8'ha7)) : (reg1450 ?
                          (7'h44) : reg1450))} : (wire1451 + {{(8'hb4),
                      (7'h40)},
                  wire1448}))))
            begin
              reg1452 <= wire1446[(1'h0):(1'h0)];
              reg1453 <= $signed(reg1452);
              reg1454 <= (wire1451 ? reg1453[(5'h13):(4'hf)] : (8'hb0));
            end
          else
            begin
              reg1452 <= $unsigned(wire1449[(3'h4):(2'h2)]);
              reg1453 <= ($unsigned(wire1449[(3'h5):(2'h3)]) & reg1452[(4'he):(4'hb)]);
              reg1454 <= {(~&((wire1447[(3'h7):(1'h1)] ?
                      wire1451 : $unsigned(wire1449)) != wire1449)),
                  (reg1453 >= wire1451[(1'h1):(1'h0)])};
              reg1455 <= ((8'ha2) ^~ (^~(|wire1448)));
            end
          reg1456 <= ((~^$unsigned(($unsigned(wire1449) ?
              (8'hac) : wire1446[(3'h5):(1'h0)]))) <<< $signed((~|{reg1455,
              {wire1451}})));
          reg1457 <= (reg1452 >= ($signed({$signed(reg1453),
                  (wire1446 || wire1448)}) ?
              ($unsigned(reg1454) ?
                  reg1456[(4'hb):(3'h6)] : (((8'hac) << reg1452) != $unsigned(wire1448))) : (reg1455[(1'h1):(1'h1)] ?
                  ({reg1452,
                      (8'ha5)} ^ (^~reg1450)) : (~^wire1447[(3'h4):(3'h4)]))));
          if ($signed($signed(($signed((wire1448 ?
              reg1455 : wire1447)) > reg1452))))
            begin
              reg1458 <= (~&wire1447);
              reg1459 <= ((-reg1450[(4'hf):(4'hc)]) >= (~|reg1450));
            end
          else
            begin
              reg1458 <= reg1459[(4'hb):(1'h0)];
              reg1459 <= (wire1448 ?
                  wire1447 : ((~$unsigned(reg1453)) ~^ (reg1456 >= $signed($signed(reg1457)))));
              reg1460 <= wire1448;
            end
        end
      else
        begin
          reg1452 <= $unsigned($unsigned($unsigned((|$unsigned(reg1458)))));
        end
    end
  assign wire1461 = (reg1454 ?
                        (~&reg1458) : (reg1458 ?
                            reg1455[(4'hc):(4'h8)] : ($unsigned((8'hb7)) ?
                                (reg1460[(2'h3):(2'h3)] >= (!reg1458)) : reg1450[(3'h7):(1'h0)])));
  always
    @(posedge clk) begin
      if ($signed({((((8'h9c) ? reg1458 : reg1458) ?
                  $unsigned(reg1452) : reg1456) ?
              $signed({reg1459, wire1449}) : (+$signed(reg1457))),
          (~&reg1458)}))
        begin
          reg1462 <= ($signed(($unsigned((8'ha3)) ?
              ((8'ha1) ?
                  $signed(reg1460) : (&wire1446)) : (!reg1460[(2'h3):(1'h0)]))) <= reg1454);
          if (reg1459)
            begin
              reg1463 <= $signed($signed(wire1461[(4'h9):(1'h1)]));
            end
          else
            begin
              reg1463 <= reg1460;
            end
          reg1464 <= (reg1452 || $signed($signed(((|(7'h41)) * wire1461))));
          if ({reg1463, reg1462})
            begin
              reg1465 <= wire1451[(1'h1):(1'h0)];
            end
          else
            begin
              reg1465 <= $signed(($signed($signed((^~reg1465))) ?
                  (+reg1454[(2'h2):(2'h2)]) : ($signed(reg1456) ?
                      {(wire1448 >>> (8'hb2)),
                          (reg1459 ?
                              reg1450 : wire1451)} : $signed($unsigned(reg1457)))));
              reg1466 <= (^($unsigned((reg1465[(1'h0):(1'h0)] + ((7'h43) <= wire1451))) ?
                  reg1463[(2'h2):(1'h1)] : $unsigned((reg1457[(2'h3):(1'h0)] - $unsigned(wire1448)))));
            end
        end
      else
        begin
          reg1462 <= (+($unsigned($unsigned(reg1456[(3'h5):(2'h2)])) ?
              (&($signed(reg1460) ?
                  $signed((8'h9d)) : wire1451[(1'h0):(1'h0)])) : ($signed(((8'hb9) ?
                      reg1466 : wire1461)) ?
                  $unsigned((reg1457 == reg1453)) : reg1463[(3'h5):(1'h1)])));
          reg1463 <= $signed(((~|$signed(reg1450[(5'h12):(3'h7)])) - {reg1454[(1'h1):(1'h0)],
              reg1455}));
          reg1464 <= $unsigned($signed((((reg1456 && reg1466) ?
              {(8'ha9), reg1458} : reg1454) >>> $unsigned((reg1464 ?
              reg1458 : reg1456)))));
          reg1465 <= reg1458[(3'h4):(2'h3)];
          reg1466 <= {$signed(wire1461[(3'h4):(1'h0)]), (8'hb5)};
        end
      reg1467 <= reg1466[(4'h9):(4'h8)];
      reg1468 <= wire1451;
      reg1469 <= $unsigned($signed($unsigned($signed(reg1454[(4'h8):(2'h3)]))));
    end
  assign wire1470 = $signed((+$unsigned({reg1464})));
  always
    @(posedge clk) begin
      if (reg1452)
        begin
          reg1471 <= reg1454[(2'h2):(2'h2)];
          if (reg1469[(5'h11):(1'h0)])
            begin
              reg1472 <= $unsigned(($unsigned($signed((|wire1447))) - ((wire1448 && (!(8'hb8))) ?
                  wire1451 : (~&$signed(wire1449)))));
            end
          else
            begin
              reg1472 <= (($signed((^~$unsigned(reg1460))) ?
                      (($signed(reg1466) ?
                          reg1471[(3'h6):(3'h5)] : {reg1466}) >= ((~^(8'haa)) ?
                          (reg1464 & reg1457) : reg1466)) : (reg1457 + (reg1458 ^~ (wire1449 && reg1472)))) ?
                  reg1452[(1'h0):(1'h0)] : ((^{{(8'had)}, (^reg1456)}) ?
                      {$unsigned(((8'ha4) || wire1447))} : $signed((~^((8'hb5) <<< reg1471)))));
              reg1473 <= wire1449;
              reg1474 <= $signed((!(~^reg1456[(4'he):(2'h2)])));
              reg1475 <= reg1466[(4'hc):(1'h1)];
            end
          reg1476 <= (((^~reg1458) == reg1473[(4'hc):(2'h2)]) ?
              $signed(wire1451[(1'h1):(1'h0)]) : ($signed(((reg1452 < wire1448) ?
                  {reg1471} : (^~wire1451))) >> ($unsigned($unsigned((8'hbb))) >> ((reg1475 ?
                      wire1461 : (8'ha3)) ?
                  $unsigned(wire1470) : (~|(8'ha9))))));
          if ((wire1451[(1'h0):(1'h0)] ?
              $signed((~|((reg1463 ? reg1463 : (8'hbf)) ?
                  {(8'h9d)} : (-reg1463)))) : (reg1460 << reg1472)))
            begin
              reg1477 <= reg1456;
              reg1478 <= $unsigned((((-(wire1447 ? wire1461 : reg1469)) ?
                      reg1462 : $unsigned($unsigned(reg1454))) ?
                  (&(wire1447[(2'h2):(2'h2)] ?
                      $signed(reg1471) : (7'h44))) : wire1447[(2'h3):(1'h0)]));
              reg1479 <= $signed((8'had));
            end
          else
            begin
              reg1477 <= reg1471;
              reg1478 <= reg1465[(1'h1):(1'h0)];
              reg1479 <= reg1464[(4'h8):(3'h7)];
            end
        end
      else
        begin
          reg1471 <= $signed($unsigned({reg1462,
              ((reg1478 ? reg1452 : (8'h9c)) + (+reg1467))}));
          if ((+reg1456[(3'h6):(3'h6)]))
            begin
              reg1472 <= $unsigned(reg1459);
              reg1473 <= {{reg1456[(4'hc):(3'h7)],
                      (({reg1474} - {reg1457, (8'ha3)}) ?
                          ($signed(reg1471) ?
                              (^~(8'hbc)) : (&reg1457)) : reg1456)},
                  $unsigned(reg1463)};
              reg1474 <= (&(({reg1455[(3'h4):(1'h0)],
                  {reg1460, reg1468}} * {$signed(reg1468),
                  {wire1446, reg1457}}) ~^ $signed(reg1453)));
              reg1475 <= $unsigned((~|reg1452));
            end
          else
            begin
              reg1472 <= (({((7'h41) ? (~^reg1456) : (-reg1453))} + reg1462) ?
                  (^~$signed((^wire1461[(1'h0):(1'h0)]))) : (^~$signed(($signed((8'ha2)) ?
                      (reg1460 > wire1448) : (~&reg1479)))));
            end
        end
    end
  assign wire1480 = $signed($unsigned(($unsigned(reg1479[(2'h2):(2'h2)]) ?
                        reg1460[(2'h2):(1'h0)] : reg1468)));
  assign wire1481 = reg1459[(3'h7):(1'h1)];
  assign wire1482 = reg1463;
  assign wire1483 = (^$unsigned($signed($signed({wire1482}))));
  assign wire1484 = ($unsigned($signed(($unsigned(reg1453) ?
                            reg1471 : $signed((8'ha5))))) ?
                        $unsigned(reg1452[(4'hf):(1'h0)]) : reg1479);
  assign wire1485 = (8'hbb);
  assign wire1486 = ((8'hbe) ?
                        (8'ha4) : (^~(((reg1464 > reg1473) + $unsigned(wire1482)) ?
                            reg1477[(4'hd):(4'h9)] : $signed((~|wire1447)))));
  assign wire1487 = $unsigned($signed((reg1475[(1'h1):(1'h1)] ?
                        $unsigned((8'ha7)) : ($signed(reg1475) ?
                            reg1471 : $unsigned(reg1472)))));
  assign wire1488 = reg1471;
  assign wire1489 = (!reg1468);
  assign wire1490 = (reg1454 != (-($signed((~reg1454)) >= ($signed(reg1465) ?
                        $unsigned(reg1456) : $signed(reg1476)))));
  assign wire1491 = reg1456[(3'h5):(2'h2)];
  assign wire1492 = (8'hab);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1726  (y, clk, wire1730, wire1729, wire1728, wire1727);
  output wire [(32'hdc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire1730;
  input wire [(4'hf):(1'h0)] wire1729;
  input wire [(2'h3):(1'h0)] wire1728;
  input wire [(4'he):(1'h0)] wire1727;
  wire [(3'h7):(1'h0)] wire1749;
  reg [(3'h5):(1'h0)] reg1748 = (1'h0);
  reg [(4'h8):(1'h0)] reg1747 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire1746;
  reg signed [(4'he):(1'h0)] reg1745 = (1'h0);
  reg [(3'h6):(1'h0)] reg1744 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1743 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1742 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1741 = (1'h0);
  reg [(5'h10):(1'h0)] reg1740 = (1'h0);
  reg [(5'h13):(1'h0)] reg1739 = (1'h0);
  reg [(5'h14):(1'h0)] reg1738 = (1'h0);
  reg [(3'h6):(1'h0)] reg1737 = (1'h0);
  reg [(5'h14):(1'h0)] reg1736 = (1'h0);
  reg [(4'ha):(1'h0)] reg1735 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1734 = (1'h0);
  reg [(4'hc):(1'h0)] reg1733 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1732 = (1'h0);
  reg [(4'he):(1'h0)] reg1731 = (1'h0);
  assign y = {wire1749,
                 reg1748,
                 reg1747,
                 wire1746,
                 reg1745,
                 reg1744,
                 reg1743,
                 reg1742,
                 reg1741,
                 reg1740,
                 reg1739,
                 reg1738,
                 reg1737,
                 reg1736,
                 reg1735,
                 reg1734,
                 reg1733,
                 reg1732,
                 reg1731,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1731 <= wire1730;
      reg1732 <= wire1728;
      reg1733 <= (({$signed($unsigned(reg1731))} ? (~wire1730) : (^wire1728)) ?
          wire1729 : (&$unsigned(wire1727[(3'h7):(3'h6)])));
      reg1734 <= ((({(wire1728 >>> wire1727)} | reg1731) ?
              $unsigned((~&{wire1729, reg1732})) : wire1727[(1'h1):(1'h1)]) ?
          ({(reg1731 == reg1731)} <<< wire1727) : ($unsigned((reg1733[(3'h5):(2'h2)] ?
                  $signed((8'h9f)) : (wire1727 ~^ wire1729))) ?
              ($signed(reg1731[(3'h5):(3'h5)]) >= ((wire1727 ?
                  reg1733 : reg1732) ^ (reg1731 ?
                  wire1730 : reg1732))) : reg1731[(1'h1):(1'h0)]));
    end
  always
    @(posedge clk) begin
      if ($signed((^~$signed($unsigned((^~reg1734))))))
        begin
          reg1735 <= ($signed($signed(((reg1732 <= (8'h9d)) ?
                  (+(7'h41)) : $unsigned(wire1730)))) ?
              $signed($signed(({reg1732, wire1729} | (reg1734 ?
                  wire1727 : reg1734)))) : $signed($signed({wire1728,
                  (^~reg1734)})));
          reg1736 <= (($signed(reg1733[(4'h8):(3'h4)]) ?
                  ($unsigned((wire1729 << wire1727)) ?
                      reg1733 : reg1733[(1'h0):(1'h0)]) : $signed($signed($unsigned(wire1727)))) ?
              (wire1729 + reg1735) : reg1733);
          reg1737 <= ((-($signed({wire1727}) ?
              (reg1733 ^ (reg1732 ? reg1731 : (8'hac))) : {(reg1734 ?
                      reg1733 : wire1727),
                  $signed(reg1733)})) * ($signed(((wire1727 ?
                  wire1727 : (8'hbc)) ?
              ((8'ha3) <<< (7'h42)) : wire1730)) + (wire1730 ?
              $signed((~&reg1735)) : $signed({reg1734}))));
          reg1738 <= wire1728;
          if ($unsigned(((^~(((8'hac) ? (8'ha0) : wire1727) ~^ (wire1730 ?
                  (8'hbd) : (8'h9e)))) ?
              (!(-$signed(reg1737))) : reg1733[(2'h2):(1'h1)])))
            begin
              reg1739 <= (reg1733 ?
                  ($signed(((^reg1731) ? (+wire1730) : reg1733)) ?
                      (~^$unsigned((reg1733 ?
                          reg1731 : wire1728))) : (({reg1732,
                              wire1728} >= $signed(reg1732)) ?
                          reg1735[(3'h4):(2'h3)] : $unsigned((wire1730 + wire1727)))) : (-((reg1732[(3'h6):(3'h5)] ?
                      {reg1731} : $unsigned(reg1731)) >>> reg1735)));
            end
          else
            begin
              reg1739 <= reg1733[(4'hb):(4'ha)];
              reg1740 <= reg1733[(3'h6):(1'h1)];
              reg1741 <= reg1733[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg1735 <= reg1736[(4'h9):(3'h6)];
          reg1736 <= $signed((($signed(reg1734) ? (+(-reg1732)) : reg1735) ?
              $signed((((8'hb7) >>> reg1731) ?
                  {reg1738} : (wire1730 ? wire1728 : reg1733))) : reg1738));
          reg1737 <= reg1731[(4'hd):(4'h8)];
          reg1738 <= $unsigned($signed(($unsigned((+reg1733)) ?
              (~^(&reg1741)) : {reg1740})));
        end
      reg1742 <= (~|reg1741[(2'h3):(1'h1)]);
      reg1743 <= (!($signed(((|wire1728) * (~|reg1742))) != wire1728));
      reg1744 <= wire1729[(1'h1):(1'h1)];
      reg1745 <= reg1737[(2'h3):(2'h3)];
    end
  assign wire1746 = $signed(wire1729[(1'h1):(1'h0)]);
  always
    @(posedge clk) begin
      reg1747 <= (8'hb5);
      reg1748 <= (($unsigned(reg1744[(3'h6):(3'h6)]) ?
          {$signed((8'hbd))} : (~$signed((wire1727 || (8'hb9))))) - (~&reg1743[(3'h4):(3'h4)]));
    end
  assign wire1749 = reg1732[(3'h6):(1'h1)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1687  (y, clk, wire1692, wire1691, wire1690, wire1689, wire1688);
  output wire [(32'hff):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire1692;
  input wire signed [(4'hd):(1'h0)] wire1691;
  input wire signed [(5'h13):(1'h0)] wire1690;
  input wire signed [(4'hb):(1'h0)] wire1689;
  input wire signed [(4'h8):(1'h0)] wire1688;
  wire signed [(5'h15):(1'h0)] wire1712;
  wire [(3'h7):(1'h0)] wire1711;
  wire [(2'h2):(1'h0)] wire1710;
  wire signed [(4'he):(1'h0)] wire1709;
  wire [(5'h15):(1'h0)] wire1708;
  reg [(5'h12):(1'h0)] reg1707 = (1'h0);
  reg [(3'h7):(1'h0)] reg1706 = (1'h0);
  reg [(3'h6):(1'h0)] reg1705 = (1'h0);
  reg [(4'he):(1'h0)] reg1704 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1703 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1702 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1701 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1700 = (1'h0);
  wire [(4'hc):(1'h0)] wire1699;
  wire signed [(4'hb):(1'h0)] wire1698;
  wire signed [(5'h13):(1'h0)] wire1697;
  wire [(2'h2):(1'h0)] wire1696;
  wire [(4'hd):(1'h0)] wire1695;
  wire signed [(4'hc):(1'h0)] wire1694;
  wire [(2'h2):(1'h0)] wire1693;
  assign y = {wire1712,
                 wire1711,
                 wire1710,
                 wire1709,
                 wire1708,
                 reg1707,
                 reg1706,
                 reg1705,
                 reg1704,
                 reg1703,
                 reg1702,
                 reg1701,
                 reg1700,
                 wire1699,
                 wire1698,
                 wire1697,
                 wire1696,
                 wire1695,
                 wire1694,
                 wire1693,
                 (1'h0)};
  assign wire1693 = $unsigned($signed(({(wire1689 - (8'hb0)),
                            (wire1688 ? wire1692 : (8'ha8))} ?
                        wire1690 : {(wire1688 ? (8'hbd) : wire1690)})));
  assign wire1694 = ($signed({wire1688[(1'h1):(1'h0)]}) ?
                        (~|wire1691) : wire1688[(1'h1):(1'h0)]);
  assign wire1695 = (wire1689[(3'h4):(3'h4)] + wire1690[(4'h9):(2'h3)]);
  assign wire1696 = $unsigned(((|wire1690) ?
                        wire1690[(5'h13):(4'hc)] : wire1694));
  assign wire1697 = $signed((8'hb7));
  assign wire1698 = ((|(&({wire1690} ^ wire1695))) ?
                        $unsigned($unsigned(wire1692[(1'h0):(1'h0)])) : wire1692);
  assign wire1699 = (wire1690[(4'h9):(2'h2)] - ($signed(wire1694) + $unsigned((&$unsigned((8'ha3))))));
  always
    @(posedge clk) begin
      reg1700 <= {$signed(wire1698),
          ((~^(-(~^(7'h42)))) ?
              wire1691[(4'h8):(1'h1)] : $unsigned(((&wire1695) ?
                  wire1690[(5'h10):(4'h8)] : $unsigned(wire1689))))};
      reg1701 <= $unsigned((wire1698[(4'hb):(1'h1)] == ({$unsigned(wire1695)} ?
          $unsigned((wire1689 ? wire1691 : (8'hb8))) : $signed(wire1691))));
      reg1702 <= $unsigned(wire1690[(5'h10):(4'ha)]);
      reg1703 <= $signed((8'haa));
      if (((|reg1700[(4'hb):(3'h5)]) ?
          ((^(wire1691[(2'h3):(2'h2)] ? reg1703 : (|wire1690))) == ((wire1696 ?
              $unsigned(reg1701) : $unsigned(wire1693)) & (|{wire1690,
              (8'hb1)}))) : (((wire1695 ? reg1702 : (reg1703 <= (8'hbf))) ?
              {$signed(wire1688),
                  reg1703} : ($signed(wire1696) ^ wire1691[(4'ha):(4'h9)])) < ($signed($signed((8'had))) || (~&wire1697)))))
        begin
          if (wire1694[(3'h4):(2'h2)])
            begin
              reg1704 <= (^$signed($unsigned(wire1692[(4'ha):(3'h6)])));
              reg1705 <= $unsigned(wire1688[(1'h0):(1'h0)]);
              reg1706 <= ($signed($unsigned((~|(reg1705 ?
                  wire1694 : (8'ha7))))) || (8'ha0));
              reg1707 <= $unsigned(reg1703);
            end
          else
            begin
              reg1704 <= ({(&reg1702),
                      $unsigned({(+wire1699), (wire1694 * reg1705)})} ?
                  $signed($signed(wire1695)) : (wire1694 >= (7'h42)));
              reg1705 <= ($signed($signed(reg1704[(2'h2):(1'h0)])) >> ((+(8'hb7)) >> (~$unsigned($signed((8'hbf))))));
              reg1706 <= (wire1699 + $unsigned((($unsigned(reg1701) || $unsigned(wire1689)) ?
                  (~|$signed(wire1697)) : (~&((8'ha6) ? (8'hb2) : (8'hb5))))));
            end
        end
      else
        begin
          reg1704 <= $signed(reg1707);
          reg1705 <= $signed(($signed((~$signed(wire1699))) || (&wire1692[(4'h8):(3'h5)])));
          reg1706 <= (8'hb2);
        end
    end
  assign wire1708 = $unsigned(((wire1691[(4'hd):(4'h8)] < (-reg1700)) >= {$signed({reg1707})}));
  assign wire1709 = (~^$signed(wire1695[(1'h1):(1'h1)]));
  assign wire1710 = $unsigned(wire1688);
  assign wire1711 = $signed($unsigned($unsigned($signed(reg1701[(4'h8):(3'h7)]))));
  assign wire1712 = ((wire1699[(1'h0):(1'h0)] ?
                        {wire1694,
                            ($signed(wire1699) ?
                                (wire1697 ?
                                    reg1705 : wire1689) : (!reg1704))} : $signed($unsigned((wire1698 ?
                            wire1696 : (8'h9e))))) - (wire1694[(3'h7):(1'h1)] ~^ (~reg1700[(2'h2):(2'h2)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1601
#( parameter param1671 = (7'h40)
, parameter param1672 = (((param1671 ? (param1671 << {(8'hae), param1671}) : (~^param1671)) ? (({param1671, param1671} * (param1671 ^~ param1671)) ? {param1671} : ((param1671 ? param1671 : param1671) ? (^~(8'ha2)) : {param1671})) : {{(+param1671), param1671}, param1671}) ? (((param1671 ? (param1671 == param1671) : ((8'haa) | param1671)) ^~ ((param1671 << (7'h41)) ~^ (-param1671))) ? (|((~|param1671) > (+param1671))) : ((~&((8'hb9) ? (8'hbc) : param1671)) ? {(^~param1671)} : (^{param1671}))) : ((&((param1671 || param1671) ? param1671 : param1671)) - ((^~(param1671 && param1671)) ? ({(8'hb8), param1671} ? ((8'hbd) <<< param1671) : (param1671 ? (8'hb2) : param1671)) : {(param1671 ? param1671 : param1671), {param1671, param1671}}))) )
(y, clk, wire1606, wire1605, wire1604, wire1603, wire1602);
  output wire [(32'h285):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire1606;
  input wire [(3'h4):(1'h0)] wire1605;
  input wire signed [(4'hb):(1'h0)] wire1604;
  input wire signed [(4'hf):(1'h0)] wire1603;
  input wire signed [(3'h7):(1'h0)] wire1602;
  wire [(5'h14):(1'h0)] wire1670;
  reg [(4'ha):(1'h0)] reg1669 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1668 = (1'h0);
  reg [(4'h8):(1'h0)] reg1667 = (1'h0);
  reg [(5'h10):(1'h0)] reg1666 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire1665;
  wire signed [(3'h4):(1'h0)] wire1664;
  wire [(4'h8):(1'h0)] wire1663;
  wire [(2'h3):(1'h0)] wire1662;
  wire signed [(4'hf):(1'h0)] wire1661;
  wire signed [(4'h9):(1'h0)] wire1660;
  wire signed [(4'hc):(1'h0)] wire1659;
  reg [(4'ha):(1'h0)] reg1658 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1657 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1656;
  reg [(3'h6):(1'h0)] reg1655 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1654 = (1'h0);
  reg [(5'h12):(1'h0)] reg1653 = (1'h0);
  reg [(4'ha):(1'h0)] reg1652 = (1'h0);
  reg [(4'hc):(1'h0)] reg1651 = (1'h0);
  reg [(3'h6):(1'h0)] reg1650 = (1'h0);
  reg [(3'h4):(1'h0)] reg1649 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1648 = (1'h0);
  reg [(3'h4):(1'h0)] reg1647 = (1'h0);
  reg [(5'h11):(1'h0)] reg1646 = (1'h0);
  reg [(5'h10):(1'h0)] reg1645 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1644 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1643 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1642 = (1'h0);
  reg [(2'h3):(1'h0)] reg1641 = (1'h0);
  reg [(5'h10):(1'h0)] reg1640 = (1'h0);
  reg [(4'hf):(1'h0)] reg1639 = (1'h0);
  reg [(3'h5):(1'h0)] reg1638 = (1'h0);
  reg [(3'h4):(1'h0)] reg1637 = (1'h0);
  reg [(3'h5):(1'h0)] reg1636 = (1'h0);
  reg [(2'h2):(1'h0)] reg1635 = (1'h0);
  reg [(4'ha):(1'h0)] reg1634 = (1'h0);
  reg [(4'he):(1'h0)] reg1633 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1632 = (1'h0);
  reg [(3'h5):(1'h0)] reg1631 = (1'h0);
  reg [(5'h14):(1'h0)] reg1630 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1629 = (1'h0);
  reg [(3'h7):(1'h0)] reg1628 = (1'h0);
  reg [(5'h14):(1'h0)] reg1627 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1626 = (1'h0);
  reg [(4'h9):(1'h0)] reg1625 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire1624;
  wire signed [(4'hb):(1'h0)] wire1623;
  wire [(4'h8):(1'h0)] wire1622;
  reg signed [(5'h10):(1'h0)] reg1621 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1620 = (1'h0);
  reg [(5'h12):(1'h0)] reg1619 = (1'h0);
  reg [(3'h4):(1'h0)] reg1618 = (1'h0);
  reg [(4'he):(1'h0)] reg1617 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1616 = (1'h0);
  reg [(3'h4):(1'h0)] reg1615 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1614 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1613 = (1'h0);
  reg [(4'hc):(1'h0)] reg1612 = (1'h0);
  wire [(4'he):(1'h0)] wire1611;
  wire [(3'h4):(1'h0)] wire1610;
  reg [(3'h6):(1'h0)] reg1609 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1608 = (1'h0);
  reg [(4'ha):(1'h0)] reg1607 = (1'h0);
  assign y = {wire1670,
                 reg1669,
                 reg1668,
                 reg1667,
                 reg1666,
                 wire1665,
                 wire1664,
                 wire1663,
                 wire1662,
                 wire1661,
                 wire1660,
                 wire1659,
                 reg1658,
                 reg1657,
                 wire1656,
                 reg1655,
                 reg1654,
                 reg1653,
                 reg1652,
                 reg1651,
                 reg1650,
                 reg1649,
                 reg1648,
                 reg1647,
                 reg1646,
                 reg1645,
                 reg1644,
                 reg1643,
                 reg1642,
                 reg1641,
                 reg1640,
                 reg1639,
                 reg1638,
                 reg1637,
                 reg1636,
                 reg1635,
                 reg1634,
                 reg1633,
                 reg1632,
                 reg1631,
                 reg1630,
                 reg1629,
                 reg1628,
                 reg1627,
                 reg1626,
                 reg1625,
                 wire1624,
                 wire1623,
                 wire1622,
                 reg1621,
                 reg1620,
                 reg1619,
                 reg1618,
                 reg1617,
                 reg1616,
                 reg1615,
                 reg1614,
                 reg1613,
                 reg1612,
                 wire1611,
                 wire1610,
                 reg1609,
                 reg1608,
                 reg1607,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1607 <= ($unsigned(($signed({wire1602,
              wire1602}) != ($unsigned(wire1603) >= (~|wire1606)))) ?
          wire1604[(4'h9):(3'h4)] : (8'hb5));
      reg1608 <= (^(-wire1603[(3'h5):(1'h1)]));
      reg1609 <= $signed(wire1602[(3'h7):(2'h3)]);
    end
  assign wire1610 = $unsigned(($signed((reg1609[(3'h5):(1'h1)] ?
                            wire1602[(1'h1):(1'h0)] : wire1602[(2'h3):(1'h0)])) ?
                        (&(wire1604 ?
                            ((8'h9f) && wire1605) : {wire1605,
                                wire1605})) : wire1606[(3'h4):(2'h2)]));
  assign wire1611 = (($unsigned(({reg1608} && $signed(wire1603))) || ((~^$unsigned(wire1603)) ?
                        reg1607 : wire1610)) - {reg1608,
                        ($signed((~&(8'ha9))) * ((reg1609 ?
                                wire1605 : wire1604) ?
                            $unsigned(wire1610) : $unsigned((8'hbc))))});
  always
    @(posedge clk) begin
      if (($unsigned(wire1602[(2'h2):(1'h0)]) ?
          wire1603[(3'h6):(2'h3)] : (&(8'h9d))))
        begin
          reg1612 <= {(($unsigned(reg1608[(3'h6):(3'h4)]) ~^ ((wire1604 ?
                      wire1610 : wire1602) & (~wire1602))) ?
                  {reg1609,
                      (&(reg1609 ?
                          wire1603 : wire1610))} : reg1609[(1'h0):(1'h0)])};
        end
      else
        begin
          if (wire1606[(1'h0):(1'h0)])
            begin
              reg1612 <= reg1608[(3'h7):(3'h6)];
              reg1613 <= $signed({((!reg1607[(4'ha):(3'h6)]) ^~ (-$unsigned(wire1606))),
                  wire1603[(4'h9):(3'h6)]});
              reg1614 <= wire1611;
              reg1615 <= (wire1610[(1'h1):(1'h0)] ?
                  wire1604[(3'h7):(2'h2)] : (wire1610 ?
                      wire1605[(2'h3):(1'h0)] : {$signed($unsigned((8'ha3))),
                          ($unsigned(reg1612) - (wire1610 && wire1602))}));
              reg1616 <= wire1602[(3'h6):(3'h5)];
            end
          else
            begin
              reg1612 <= ((&{(wire1602[(1'h1):(1'h0)] ?
                      $signed(wire1603) : $unsigned(reg1616)),
                  (|(wire1604 != reg1609))}) <<< wire1605);
            end
          reg1617 <= (~|($signed((wire1602[(2'h3):(2'h3)] ^~ reg1612)) ?
              $unsigned((wire1604 << {(8'hae),
                  wire1603})) : $signed(($signed(reg1609) > {reg1616,
                  reg1615}))));
          reg1618 <= reg1609[(1'h1):(1'h1)];
          reg1619 <= (reg1608 ? reg1618 : wire1610);
          reg1620 <= $unsigned($unsigned(wire1610[(2'h3):(1'h0)]));
        end
      reg1621 <= $unsigned(reg1620);
    end
  assign wire1622 = $unsigned(reg1607);
  assign wire1623 = $signed($unsigned(wire1611));
  assign wire1624 = wire1610;
  always
    @(posedge clk) begin
      if ({$signed((~{reg1609, {wire1605, reg1613}})), (8'hbf)})
        begin
          reg1625 <= (reg1609[(3'h6):(1'h0)] ?
              $signed($signed(wire1610)) : $signed(reg1615[(1'h0):(1'h0)]));
          if ($signed($unsigned($signed((reg1621 || $unsigned((8'h9d)))))))
            begin
              reg1626 <= {reg1616[(3'h4):(2'h3)], reg1625[(1'h0):(1'h0)]};
              reg1627 <= $signed({$unsigned(wire1604), wire1611});
              reg1628 <= (^reg1608[(1'h1):(1'h1)]);
              reg1629 <= {(|({((8'hb5) ? reg1613 : reg1616)} << ((+wire1624) ?
                      (wire1623 ? reg1607 : reg1613) : reg1617)))};
              reg1630 <= reg1629;
            end
          else
            begin
              reg1626 <= (({reg1619[(3'h7):(3'h4)],
                  reg1627} == $unsigned({$signed(reg1615)})) && $unsigned(wire1603));
              reg1627 <= $unsigned(($unsigned((-(reg1616 ?
                  wire1624 : reg1617))) == reg1621[(3'h6):(1'h1)]));
              reg1628 <= $signed(($signed(wire1602[(1'h1):(1'h1)]) ^~ (($unsigned(reg1608) ?
                      wire1603[(4'h9):(1'h0)] : wire1603) ?
                  ((reg1613 ? (8'hb8) : reg1621) ?
                      (reg1612 ?
                          reg1609 : wire1624) : reg1619[(4'hf):(4'hb)]) : reg1626)));
              reg1629 <= $unsigned($signed(wire1606));
            end
          reg1631 <= $signed((7'h42));
          if ($signed((wire1603 * (^~reg1613[(3'h4):(2'h2)]))))
            begin
              reg1632 <= reg1614[(3'h6):(3'h5)];
              reg1633 <= {reg1632[(4'h9):(3'h7)]};
              reg1634 <= (^~{(8'hba),
                  (wire1604[(3'h7):(1'h0)] ?
                      ($unsigned(wire1606) ?
                          reg1614 : $unsigned(reg1612)) : reg1614)});
              reg1635 <= $unsigned(((~^($unsigned(reg1612) > (reg1630 + wire1606))) ?
                  reg1607 : $signed(($signed(reg1613) << $signed(reg1608)))));
            end
          else
            begin
              reg1632 <= (-wire1611);
              reg1633 <= (+$signed(((|reg1629[(1'h1):(1'h0)]) ?
                  {reg1614,
                      ((8'ha0) ?
                          (8'hbf) : reg1614)} : reg1617[(3'h5):(1'h1)])));
              reg1634 <= reg1626;
              reg1635 <= (wire1604 != ({(!reg1621), {reg1613}} ?
                  reg1613 : reg1632));
            end
        end
      else
        begin
          reg1625 <= (^{$unsigned(reg1614[(1'h0):(1'h0)]), wire1610});
        end
      reg1636 <= ($signed((&(~&{wire1610,
          wire1605}))) ~^ ((reg1616 == (reg1609 > (+(7'h40)))) ?
          ($signed((reg1629 >>> reg1625)) ?
              reg1631[(1'h1):(1'h1)] : reg1612[(1'h0):(1'h0)]) : $signed({$signed(reg1629),
              (wire1603 << reg1625)})));
    end
  always
    @(posedge clk) begin
      if (((+(reg1631 ^ reg1615)) ? wire1605 : $signed((~^reg1613))))
        begin
          if ({(7'h42)})
            begin
              reg1637 <= $unsigned(reg1636[(1'h1):(1'h1)]);
              reg1638 <= $signed($unsigned({$signed({reg1636})}));
              reg1639 <= (((|{$unsigned(wire1624)}) ?
                  (^$signed((reg1613 ?
                      reg1638 : reg1615))) : (8'hb4)) == wire1622[(3'h6):(3'h5)]);
              reg1640 <= {$unsigned((7'h44)),
                  (^(($signed(wire1623) << $signed(reg1638)) + $unsigned((wire1602 >= reg1639))))};
              reg1641 <= (reg1615 ?
                  (|$unsigned(reg1608[(3'h6):(3'h5)])) : {(~$signed((reg1633 ^ (8'ha1)))),
                      reg1628[(3'h6):(2'h2)]});
            end
          else
            begin
              reg1637 <= (^~wire1606[(4'h9):(3'h4)]);
              reg1638 <= $unsigned(reg1616[(4'hc):(2'h3)]);
              reg1639 <= (~(8'ha3));
            end
          reg1642 <= (|(&(($signed(reg1638) ^~ (reg1609 ?
              reg1614 : wire1602)) ^~ $signed(reg1641[(2'h3):(2'h2)]))));
          if ((((8'hbe) >>> $signed($signed((reg1636 >= reg1617)))) >> reg1619[(4'hf):(4'hf)]))
            begin
              reg1643 <= (wire1622[(3'h7):(3'h4)] || ($unsigned($unsigned((reg1616 ?
                      wire1605 : wire1602))) ?
                  {(((8'hbe) > reg1638) ?
                          (reg1638 ? reg1617 : reg1626) : {(8'hb5), (8'h9e)}),
                      $signed((wire1611 ?
                          reg1629 : reg1616))} : $unsigned($unsigned((reg1617 < reg1621)))));
            end
          else
            begin
              reg1643 <= reg1627;
              reg1644 <= ($signed($signed($unsigned((~|wire1624)))) ?
                  reg1609[(2'h2):(1'h0)] : reg1616);
            end
        end
      else
        begin
          if (((^wire1623) ?
              (reg1617[(3'h6):(2'h3)] < $unsigned(($signed(reg1641) ?
                  reg1628 : (reg1638 ?
                      reg1613 : (8'hab))))) : {(^reg1621[(4'hb):(2'h2)]),
                  $unsigned($unsigned({reg1612, reg1607}))}))
            begin
              reg1637 <= ($unsigned({($unsigned(reg1614) ?
                      reg1629 : reg1614[(3'h4):(1'h0)]),
                  $signed(reg1644[(4'hc):(2'h2)])}) != ((-reg1608) ?
                  reg1641 : (^reg1644)));
            end
          else
            begin
              reg1637 <= {(reg1642 ~^ (8'hab)),
                  ((($unsigned((8'ha1)) == $signed(reg1631)) >= ({(8'ha2),
                          reg1626} & (reg1643 ? reg1626 : wire1602))) ?
                      {(^~$signed(reg1644))} : (((reg1616 ?
                              reg1630 : wire1606) + reg1632[(1'h0):(1'h0)]) ?
                          $unsigned((^wire1604)) : reg1636))};
            end
          reg1638 <= $unsigned($unsigned($unsigned(reg1629[(3'h4):(1'h1)])));
          if (((!$signed($unsigned($unsigned((8'h9f))))) ?
              (({$unsigned((8'ha1)), reg1629} >= (reg1638[(2'h3):(1'h1)] ?
                      $unsigned((8'ha6)) : {reg1636})) ?
                  (7'h42) : $unsigned($unsigned((reg1631 && reg1639)))) : ($signed(reg1636) ?
                  ({wire1624} ?
                      $unsigned(wire1623[(3'h4):(3'h4)]) : (!$signed(reg1629))) : (8'ha8))))
            begin
              reg1639 <= $signed($signed($signed(reg1643)));
            end
          else
            begin
              reg1639 <= reg1621[(1'h0):(1'h0)];
              reg1640 <= (-(~|({reg1641} | reg1627[(4'hc):(2'h2)])));
              reg1641 <= $unsigned(reg1634[(3'h5):(3'h5)]);
              reg1642 <= $unsigned(reg1612);
              reg1643 <= ((($signed((reg1607 ? reg1625 : reg1616)) ?
                  ($signed((8'ha9)) ? reg1631 : (~^wire1603)) : ({reg1616,
                          (8'had)} ?
                      $signed((7'h41)) : reg1631)) <<< ((~$unsigned(wire1602)) & {((8'hbe) * (8'hab)),
                  (wire1610 << reg1643)})) + ($signed($unsigned($unsigned(reg1626))) >> $unsigned(reg1642)));
            end
          reg1644 <= (|(((^(-reg1639)) == (-reg1612[(1'h0):(1'h0)])) ?
              (~^(reg1640[(4'he):(4'hc)] ?
                  (wire1605 | (8'haa)) : reg1612)) : (reg1613 <<< ({(8'ha6)} && $unsigned(reg1618)))));
        end
      if ($signed($signed(wire1603[(4'hd):(4'hb)])))
        begin
          reg1645 <= $unsigned((8'h9d));
          reg1646 <= ((&(((reg1608 ? reg1620 : reg1618) ?
                  (reg1642 ? reg1620 : (8'hb2)) : reg1633[(4'h9):(3'h6)]) ?
              $signed((!reg1612)) : {$signed(reg1635)})) >= ((reg1631[(2'h3):(2'h2)] < $unsigned(wire1604[(3'h7):(3'h7)])) <<< (wire1604 ?
              (8'hbe) : (reg1634 ? $signed(reg1637) : $unsigned(reg1642)))));
          reg1647 <= (^reg1629[(3'h7):(1'h0)]);
        end
      else
        begin
          reg1645 <= (|(~^$signed(($unsigned(reg1614) ?
              $signed((8'ha0)) : ((8'ha5) ^ wire1611)))));
          if (wire1622)
            begin
              reg1646 <= (reg1626 < $signed((((-reg1647) ?
                      (reg1620 >= reg1644) : $unsigned((8'ha4))) ?
                  $unsigned((reg1633 >>> reg1638)) : {$unsigned(reg1636)})));
              reg1647 <= reg1629;
              reg1648 <= $signed((~&(-(8'ha7))));
              reg1649 <= wire1622[(1'h0):(1'h0)];
              reg1650 <= {{((((8'ha9) ? wire1610 : (8'h9f)) < (+wire1624)) ?
                          ((reg1608 > reg1640) == reg1634[(4'h8):(1'h1)]) : wire1604)},
                  $signed(wire1605[(3'h4):(3'h4)])};
            end
          else
            begin
              reg1646 <= $unsigned((+(wire1611[(4'ha):(3'h7)] <= $signed(((8'hac) >>> wire1604)))));
            end
        end
      reg1651 <= ({($signed(((8'haf) ^ wire1622)) ?
                  $signed($unsigned(reg1614)) : reg1632)} ?
          (~^({((8'hb7) ? wire1622 : reg1615),
              $unsigned(reg1614)} || ({reg1628} >>> $unsigned(reg1648)))) : ($unsigned((^~(8'hab))) ?
              reg1608 : $unsigned($unsigned((reg1607 | wire1602)))));
      if ($unsigned(wire1611[(4'hd):(1'h0)]))
        begin
          reg1652 <= ($signed(((!(8'hb9)) >>> wire1611)) ?
              (reg1649[(1'h0):(1'h0)] ?
                  $unsigned((((8'ha9) >> reg1639) && (wire1611 == reg1609))) : wire1623) : ($unsigned(((reg1629 ?
                  reg1616 : reg1633) * (reg1625 ~^ wire1623))) * {$signed((wire1610 ?
                      wire1623 : reg1646)),
                  (+reg1637[(2'h3):(1'h1)])}));
          reg1653 <= {reg1633[(4'hd):(4'hb)]};
        end
      else
        begin
          reg1652 <= (($signed($unsigned(reg1648[(1'h0):(1'h0)])) ?
                  (8'haa) : reg1625) ?
              $signed((({(7'h42)} * $signed((7'h44))) < $unsigned($unsigned(reg1636)))) : reg1650);
          reg1653 <= (($unsigned((^~(reg1620 ?
                  reg1642 : (8'hb3)))) | ((~|((8'hb7) ?
                  (8'haf) : reg1642)) == $signed({wire1624}))) ?
              $unsigned(reg1635[(2'h2):(1'h1)]) : (~&($unsigned($signed(reg1637)) > (^{reg1630,
                  reg1641}))));
          reg1654 <= ((^~reg1652[(3'h4):(2'h2)]) ~^ reg1607);
        end
      reg1655 <= ($unsigned(reg1653[(4'hc):(4'h8)]) ?
          reg1608[(3'h4):(2'h3)] : reg1629);
    end
  assign wire1656 = (|$unsigned(reg1615[(2'h2):(1'h1)]));
  always
    @(posedge clk) begin
      reg1657 <= wire1622;
      reg1658 <= wire1602;
    end
  assign wire1659 = {reg1625[(3'h7):(2'h2)]};
  assign wire1660 = reg1635[(2'h2):(1'h1)];
  assign wire1661 = $signed(({reg1632, (|{reg1655, reg1612})} ?
                        {((reg1652 + wire1605) && (~&reg1650))} : (-(8'hba))));
  assign wire1662 = (+(+(|$unsigned((~(8'ha3))))));
  assign wire1663 = (($signed(($unsigned(wire1603) < (reg1642 + reg1629))) < ($signed(reg1652[(3'h4):(3'h4)]) > ($signed(wire1602) || reg1640))) ?
                        reg1631 : wire1606);
  assign wire1664 = reg1636[(2'h2):(2'h2)];
  assign wire1665 = $signed(({$unsigned((&wire1606)), reg1655} <<< reg1618));
  always
    @(posedge clk) begin
      reg1666 <= {((^$signed($signed(reg1637))) < ((reg1636 < (reg1648 ?
                  wire1603 : reg1635)) ?
              ($signed(reg1640) > $unsigned((8'hbc))) : $signed({(8'ha3)})))};
      reg1667 <= ($signed(wire1606) >= ((8'ha4) ^~ $unsigned($signed(reg1635[(2'h2):(2'h2)]))));
      reg1668 <= (reg1654 ? (8'ha8) : wire1624[(1'h1):(1'h0)]);
      reg1669 <= $signed(reg1651[(1'h0):(1'h0)]);
    end
  assign wire1670 = reg1636[(1'h1):(1'h1)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1573
#( parameter param1587 = ((~{(&{(8'hba), (8'hbd)})}) ? (((((8'hb8) > (8'hac)) <<< (&(7'h44))) >> {((8'had) ? (8'hbc) : (8'hba)), ((8'ha3) ? (8'haa) : (8'haa))}) >>> ((((8'hb4) <<< (8'haa)) << ((8'hb0) << (8'h9e))) << ((!(8'ha8)) != ((8'hab) ? (8'ha2) : (8'hb6))))) : (~&(+((-(7'h43)) + ((8'hae) != (8'haa))))))
, parameter param1588 = {((({param1587} ? param1587 : (param1587 <<< param1587)) ? (((8'hbd) | param1587) ? (param1587 <= param1587) : {param1587, param1587}) : (^~((8'h9c) > param1587))) ? param1587 : (^~({param1587, param1587} != param1587))), (+param1587)} )
(y, clk, wire1578, wire1577, wire1576, wire1575, wire1574);
  output wire [(32'h5e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire1578;
  input wire [(5'h12):(1'h0)] wire1577;
  input wire [(4'hc):(1'h0)] wire1576;
  input wire signed [(5'h10):(1'h0)] wire1575;
  input wire [(3'h5):(1'h0)] wire1574;
  wire signed [(4'h9):(1'h0)] wire1586;
  wire signed [(3'h7):(1'h0)] wire1585;
  wire [(5'h15):(1'h0)] wire1584;
  wire [(3'h6):(1'h0)] wire1583;
  wire [(3'h7):(1'h0)] wire1582;
  wire signed [(4'h9):(1'h0)] wire1581;
  wire [(4'he):(1'h0)] wire1580;
  wire signed [(5'h14):(1'h0)] wire1579;
  assign y = {wire1586,
                 wire1585,
                 wire1584,
                 wire1583,
                 wire1582,
                 wire1581,
                 wire1580,
                 wire1579,
                 (1'h0)};
  assign wire1579 = $unsigned((!((wire1577[(4'hc):(3'h6)] ?
                            (wire1576 ^ wire1577) : $signed((8'hb5))) ?
                        $signed((wire1576 ?
                            (8'hbd) : wire1577)) : {wire1577})));
  assign wire1580 = $signed(wire1574);
  assign wire1581 = ((+$unsigned((~|wire1580[(4'hb):(4'h9)]))) ~^ (~&($signed((~wire1578)) ?
                        $unsigned($signed((8'hb0))) : $signed($unsigned(wire1575)))));
  assign wire1582 = (($unsigned((wire1577[(5'h11):(1'h0)] <<< wire1578)) ^ (^~(|(wire1577 ?
                        (8'ha3) : (8'hb4))))) >> $unsigned((($unsigned((8'ha6)) ?
                            $signed(wire1574) : $signed(wire1576)) ?
                        wire1580 : (8'hab))));
  assign wire1583 = wire1575[(2'h3):(1'h0)];
  assign wire1584 = (~wire1574);
  assign wire1585 = wire1577;
  assign wire1586 = (^~wire1584);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1815
#( parameter param1825 = ({(((~&(8'haf)) ? ((8'h9e) ? (7'h42) : (8'hb2)) : {(8'h9f)}) ? (|(-(8'h9c))) : (8'h9d)), (((~(8'ha8)) ? ((7'h43) ^ (8'h9d)) : ((8'hae) ^ (8'haf))) ? {{(8'hb5), (8'hb2)}, (8'hbe)} : (((8'hbd) ? (7'h41) : (8'ha3)) ~^ ((8'haa) ? (8'had) : (8'h9e))))} && {(((8'h9c) ? ((7'h42) & (8'ha9)) : ((8'ha1) | (8'haa))) ? {(-(8'hb3)), (!(8'h9e))} : {(~|(8'ha8)), ((8'hb0) ? (8'hba) : (8'haa))})})
, parameter param1826 = (((^~{(param1825 | param1825)}) != (~^{param1825})) >> param1825) )
(y, clk, wire1819, wire1818, wire1817, wire1816);
  output wire [(32'h53):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire1819;
  input wire signed [(4'ha):(1'h0)] wire1818;
  input wire [(5'h12):(1'h0)] wire1817;
  input wire [(2'h2):(1'h0)] wire1816;
  wire signed [(5'h11):(1'h0)] wire1824;
  wire signed [(4'he):(1'h0)] wire1823;
  wire signed [(4'hd):(1'h0)] wire1822;
  wire signed [(5'h15):(1'h0)] wire1821;
  wire [(5'h11):(1'h0)] wire1820;
  assign y = {wire1824, wire1823, wire1822, wire1821, wire1820, (1'h0)};
  assign wire1820 = wire1817;
  assign wire1821 = ($unsigned((wire1819[(3'h5):(2'h2)] ?
                        ((^~wire1818) ?
                            ((8'had) ?
                                (8'haa) : wire1820) : (&wire1818)) : wire1816[(1'h0):(1'h0)])) + ($signed($signed($unsigned((8'hac)))) ?
                        wire1816[(1'h0):(1'h0)] : (((8'ha2) ?
                            (wire1820 ? wire1819 : wire1816) : (wire1818 ?
                                wire1819 : wire1819)) >>> $unsigned((wire1817 & wire1816)))));
  assign wire1822 = wire1818;
  assign wire1823 = ((wire1817[(1'h1):(1'h0)] ?
                        wire1818 : wire1821) == wire1819[(3'h4):(3'h4)]);
  assign wire1824 = (wire1818 > wire1817);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1792  (y, clk, wire1797, wire1796, wire1795, wire1794, wire1793);
  output wire [(32'h97):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire1797;
  input wire [(5'h10):(1'h0)] wire1796;
  input wire signed [(4'ha):(1'h0)] wire1795;
  input wire [(4'hd):(1'h0)] wire1794;
  input wire signed [(4'h9):(1'h0)] wire1793;
  wire signed [(4'hd):(1'h0)] wire1812;
  wire [(2'h2):(1'h0)] wire1811;
  wire signed [(4'he):(1'h0)] wire1810;
  wire [(4'hf):(1'h0)] wire1809;
  wire [(4'h8):(1'h0)] wire1808;
  wire signed [(4'hd):(1'h0)] wire1807;
  wire signed [(4'ha):(1'h0)] wire1806;
  wire [(3'h5):(1'h0)] wire1805;
  wire signed [(2'h3):(1'h0)] wire1804;
  wire [(4'ha):(1'h0)] wire1803;
  wire [(4'hf):(1'h0)] wire1802;
  wire signed [(4'hf):(1'h0)] wire1801;
  wire signed [(4'hf):(1'h0)] wire1800;
  wire signed [(3'h5):(1'h0)] wire1799;
  wire [(3'h7):(1'h0)] wire1798;
  assign y = {wire1812,
                 wire1811,
                 wire1810,
                 wire1809,
                 wire1808,
                 wire1807,
                 wire1806,
                 wire1805,
                 wire1804,
                 wire1803,
                 wire1802,
                 wire1801,
                 wire1800,
                 wire1799,
                 wire1798,
                 (1'h0)};
  assign wire1798 = $signed(((+wire1796) + wire1795[(1'h1):(1'h0)]));
  assign wire1799 = (($signed(wire1798) < (~$signed((~^wire1798)))) << ({{wire1796},
                            wire1795} ?
                        $signed(wire1795[(4'h8):(3'h6)]) : $unsigned($unsigned((wire1798 >>> wire1794)))));
  assign wire1800 = ((wire1796 ^ wire1799) ~^ ($signed($signed((+wire1793))) - ($unsigned({wire1797,
                        wire1799}) * (~&wire1799))));
  assign wire1801 = wire1793[(3'h6):(1'h1)];
  assign wire1802 = $unsigned((wire1800[(4'ha):(2'h3)] ?
                        {$signed($signed(wire1801))} : (~&({wire1795} << $unsigned(wire1800)))));
  assign wire1803 = ((!{(wire1799[(1'h0):(1'h0)] | $signed(wire1802)),
                            {wire1797}}) ?
                        wire1800 : $signed((($unsigned(wire1797) ?
                            wire1795 : $signed(wire1799)) || (8'hab))));
  assign wire1804 = (~{wire1796[(3'h4):(2'h2)]});
  assign wire1805 = (!($signed($unsigned($unsigned(wire1794))) >> {$signed(wire1800[(3'h6):(3'h5)])}));
  assign wire1806 = ({$unsigned((&(wire1805 < wire1796)))} & wire1800[(3'h7):(2'h2)]);
  assign wire1807 = {wire1801[(1'h0):(1'h0)],
                        (wire1796 * (((~^wire1802) > $signed(wire1796)) <<< {wire1794}))};
  assign wire1808 = ($signed(wire1801) ?
                        wire1807 : $signed($signed((wire1806 ?
                            wire1796 : (wire1800 ? wire1807 : wire1799)))));
  assign wire1809 = (-wire1801);
  assign wire1810 = {{($unsigned((-wire1796)) ?
                                $signed($signed(wire1801)) : ((+wire1807) ?
                                    $signed((8'ha0)) : (wire1808 ?
                                        wire1796 : wire1795)))}};
  assign wire1811 = wire1800;
  assign wire1812 = $unsigned({(($unsigned(wire1800) < wire1797) || $signed({wire1806,
                            wire1807}))});
endmodule