(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param4582 = (+{(((~&(8'ha7)) == ((8'hb5) ? (8'h9e) : (8'hb1))) ? ((~&(7'h44)) << (^~(8'haa))) : (~&{(7'h41)}))}) )
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h52):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire4;
  input wire signed [(5'h13):(1'h0)] wire3;
  input wire signed [(5'h18):(1'h0)] wire2;
  input wire signed [(5'h13):(1'h0)] wire1;
  input wire [(5'h14):(1'h0)] wire0;
  wire [(5'h12):(1'h0)] wire4581;
  wire [(5'h10):(1'h0)] wire4579;
  reg [(5'h19):(1'h0)] reg4578 = (1'h0);
  reg [(5'h12):(1'h0)] reg4577 = (1'h0);
  wire [(3'h4):(1'h0)] wire4575;
  assign y = {wire4581, wire4579, reg4578, reg4577, wire4575, (1'h0)};
  module5 modinst4576 (wire4575, clk, wire2, wire3, wire0, wire4);
  always
    @(posedge clk) begin
      reg4577 <= wire3;
      reg4578 <= (reg4577 > wire1[(4'h9):(4'h8)]);
    end
  module4117 modinst4580 (wire4579, clk, wire4, wire2, wire3, reg4578);
  assign wire4581 = $unsigned($unsigned($unsigned(wire4575[(1'h0):(1'h0)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module5  (y, clk, wire9, wire8, wire7, wire6);
  output wire [(32'h742):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire9;
  input wire signed [(3'h7):(1'h0)] wire8;
  input wire [(5'h14):(1'h0)] wire7;
  input wire [(4'hd):(1'h0)] wire6;
  reg [(5'h16):(1'h0)] reg4574 = (1'h0);
  reg [(5'h16):(1'h0)] reg4573 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4572 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4571 = (1'h0);
  reg [(5'h11):(1'h0)] reg4570 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire4569;
  reg signed [(2'h2):(1'h0)] reg4568 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg4567 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4566 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar4565 = (1'h0);
  reg [(3'h4):(1'h0)] reg4564 = (1'h0);
  reg [(5'h1a):(1'h0)] reg4563 = (1'h0);
  reg [(5'h17):(1'h0)] reg4562 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4561 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4560 = (1'h0);
  reg [(3'h4):(1'h0)] reg4559 = (1'h0);
  reg [(5'h16):(1'h0)] forvar4558 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire4557;
  wire signed [(5'h18):(1'h0)] wire4556;
  reg signed [(2'h2):(1'h0)] reg4555 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg4554 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4553 = (1'h0);
  reg [(5'h12):(1'h0)] reg4552 = (1'h0);
  reg [(5'h18):(1'h0)] reg4551 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg4550 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4549 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4548 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4547 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4546 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4545 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4544 = (1'h0);
  wire [(2'h2):(1'h0)] wire4542;
  reg signed [(5'h10):(1'h0)] reg4541 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg4540 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4539 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4538 = (1'h0);
  reg [(2'h3):(1'h0)] reg4537 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg4536 = (1'h0);
  reg [(5'h18):(1'h0)] reg4535 = (1'h0);
  reg [(5'h1a):(1'h0)] reg4534 = (1'h0);
  reg [(2'h3):(1'h0)] reg4533 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4532 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4531 = (1'h0);
  reg [(5'h13):(1'h0)] reg4530 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg4529 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar4528 = (1'h0);
  reg [(5'h19):(1'h0)] reg4527 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg4526 = (1'h0);
  reg [(5'h11):(1'h0)] reg4525 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4524 = (1'h0);
  reg [(4'h9):(1'h0)] reg4523 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg4522 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4521 = (1'h0);
  reg [(4'he):(1'h0)] reg4520 = (1'h0);
  reg [(3'h4):(1'h0)] reg4519 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4518 = (1'h0);
  reg [(2'h3):(1'h0)] reg4517 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4516 = (1'h0);
  reg [(5'h14):(1'h0)] reg4515 = (1'h0);
  reg [(5'h18):(1'h0)] reg4514 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4513 = (1'h0);
  reg [(5'h12):(1'h0)] reg4512 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4511 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4510 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4509 = (1'h0);
  reg [(4'he):(1'h0)] reg4508 = (1'h0);
  reg [(5'h19):(1'h0)] forvar4507 = (1'h0);
  reg [(5'h13):(1'h0)] reg4506 = (1'h0);
  reg [(5'h1a):(1'h0)] reg4505 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4504 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4503 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4502 = (1'h0);
  reg [(4'h8):(1'h0)] reg4501 = (1'h0);
  reg [(3'h7):(1'h0)] reg4500 = (1'h0);
  reg [(4'h9):(1'h0)] reg4499 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4498 = (1'h0);
  reg [(4'he):(1'h0)] reg4497 = (1'h0);
  reg [(4'hf):(1'h0)] reg4496 = (1'h0);
  reg [(5'h1a):(1'h0)] reg4495 = (1'h0);
  wire [(5'h14):(1'h0)] wire4494;
  wire signed [(4'hd):(1'h0)] wire4493;
  wire [(4'hc):(1'h0)] wire4492;
  reg signed [(3'h4):(1'h0)] reg4491 = (1'h0);
  reg [(5'h12):(1'h0)] reg4490 = (1'h0);
  reg [(5'h11):(1'h0)] reg4489 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4488 = (1'h0);
  wire [(5'h19):(1'h0)] wire4487;
  wire [(5'h14):(1'h0)] wire4447;
  reg [(4'hf):(1'h0)] reg16 = (1'h0);
  reg [(5'h12):(1'h0)] reg15 = (1'h0);
  reg [(5'h11):(1'h0)] reg14 = (1'h0);
  reg [(5'h17):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg12 = (1'h0);
  reg [(5'h1a):(1'h0)] reg11 = (1'h0);
  wire signed [(5'h19):(1'h0)] wire10;
  wire signed [(3'h6):(1'h0)] wire4449;
  wire [(4'hb):(1'h0)] wire4451;
  wire [(5'h13):(1'h0)] wire4453;
  reg [(5'h18):(1'h0)] reg4454 = (1'h0);
  reg [(5'h12):(1'h0)] reg4455 = (1'h0);
  reg [(5'h14):(1'h0)] reg4456 = (1'h0);
  reg [(5'h17):(1'h0)] forvar4457 = (1'h0);
  reg [(5'h14):(1'h0)] forvar4458 = (1'h0);
  reg [(5'h11):(1'h0)] reg4459 = (1'h0);
  reg [(3'h7):(1'h0)] reg4460 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg4461 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4462 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4463 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4464 = (1'h0);
  reg [(4'hd):(1'h0)] reg4465 = (1'h0);
  reg [(5'h16):(1'h0)] reg4466 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4467 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4468 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4469 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4470 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4471 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg4472 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4473 = (1'h0);
  reg [(2'h2):(1'h0)] reg4474 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4475 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4476 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg4477 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg4478 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg4479 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4480 = (1'h0);
  reg [(4'hd):(1'h0)] reg4481 = (1'h0);
  reg [(3'h5):(1'h0)] reg4482 = (1'h0);
  reg [(4'hd):(1'h0)] reg4483 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg4484 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire4485;
  assign y = {reg4574,
                 reg4573,
                 reg4572,
                 reg4571,
                 reg4570,
                 wire4569,
                 reg4568,
                 reg4567,
                 reg4566,
                 forvar4565,
                 reg4564,
                 reg4563,
                 reg4562,
                 reg4561,
                 forvar4560,
                 reg4559,
                 forvar4558,
                 wire4557,
                 wire4556,
                 reg4555,
                 reg4554,
                 reg4553,
                 reg4552,
                 reg4551,
                 reg4550,
                 reg4549,
                 forvar4548,
                 forvar4547,
                 forvar4546,
                 reg4545,
                 reg4544,
                 wire4542,
                 reg4541,
                 reg4540,
                 reg4539,
                 reg4538,
                 reg4537,
                 reg4536,
                 reg4535,
                 reg4534,
                 reg4533,
                 reg4532,
                 reg4531,
                 reg4530,
                 reg4529,
                 forvar4528,
                 reg4527,
                 reg4526,
                 reg4525,
                 forvar4524,
                 reg4523,
                 reg4522,
                 reg4521,
                 reg4520,
                 reg4519,
                 forvar4518,
                 reg4517,
                 forvar4516,
                 reg4515,
                 reg4514,
                 reg4513,
                 reg4512,
                 reg4511,
                 reg4510,
                 forvar4509,
                 reg4508,
                 forvar4507,
                 reg4506,
                 reg4505,
                 forvar4504,
                 forvar4503,
                 forvar4502,
                 reg4501,
                 reg4500,
                 reg4499,
                 reg4498,
                 reg4497,
                 reg4496,
                 reg4495,
                 wire4494,
                 wire4493,
                 wire4492,
                 reg4491,
                 reg4490,
                 reg4489,
                 forvar4488,
                 wire4487,
                 wire4447,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 wire10,
                 wire4449,
                 wire4451,
                 wire4453,
                 reg4454,
                 reg4455,
                 reg4456,
                 forvar4457,
                 forvar4458,
                 reg4459,
                 reg4460,
                 reg4461,
                 reg4462,
                 reg4463,
                 forvar4464,
                 reg4465,
                 reg4466,
                 reg4467,
                 reg4468,
                 forvar4469,
                 reg4470,
                 reg4471,
                 reg4472,
                 reg4473,
                 reg4474,
                 reg4475,
                 reg4476,
                 reg4477,
                 reg4478,
                 reg4479,
                 forvar4480,
                 reg4481,
                 reg4482,
                 reg4483,
                 reg4484,
                 wire4485,
                 (1'h0)};
  assign wire10 = $unsigned(wire8);
  always
    @(posedge clk) begin
      reg11 <= wire10[(3'h4):(2'h3)];
      reg12 <= (-(|$unsigned((~(^wire10)))));
      reg13 <= reg12;
      reg14 <= {($unsigned(((reg13 >> wire10) ? (~&wire8) : "")) ?
              wire10[(3'h4):(2'h3)] : {(((7'h45) ?
                      (8'hb4) : wire9) ^ (wire9 <= reg13))})};
      reg15 <= wire6;
      reg16 <= ({reg13, reg11[(1'h0):(1'h0)]} ?
          ((^~{$unsigned(reg14)}) ?
              {(-$signed(reg13)),
                  $unsigned((wire10 ?
                      reg15 : wire10))} : $signed(wire8[(1'h1):(1'h1)])) : wire7);
    end
  module17 modinst4448 (wire4447, clk, wire7, wire10, reg14, reg12, reg11);
  module1483 modinst4450 (.wire1485(wire10), .wire1486(reg14), .wire1487(reg15), .clk(clk), .wire1484(reg11), .y(wire4449));
  module93 modinst4452 (.y(wire4451), .wire97(wire7), .clk(clk), .wire94(wire6), .wire96(reg13), .wire95(reg15));
  assign wire4453 = (8'hbc);
  always
    @(posedge clk) begin
      reg4454 <= (^~(~(!reg16[(4'hd):(1'h0)])));
      reg4455 <= wire4451[(4'hb):(2'h3)];
      reg4456 = ((("tNiqIua1ekHlGSsDJP37QY" ^ reg15) > (^reg13[(4'hc):(3'h7)])) ^~ ("bXUzk1H2vyvnbepdA" ?
          (^~(~&(^reg15))) : ""));
      for (forvar4457 = (1'h0); (forvar4457 < (3'h4)); forvar4457 = (forvar4457 + (1'h1)))
        begin
          for (forvar4458 = (1'h0); (forvar4458 < (3'h4)); forvar4458 = (forvar4458 + (1'h1)))
            begin
              reg4459 <= {(|(8'haa)), wire4447};
              reg4460 <= $signed(((("ZIQ4Mm6h" && $unsigned(reg4459)) ?
                      "4KLGNRClFt0PzkcPmC3P4vn" : reg16[(2'h3):(1'h1)]) ?
                  "lbM95U79x8WktqqQMvOmi" : "DNc4OvKwQLMqZsLAzCP"));
              reg4461 <= wire4447;
              reg4462 <= ({(({reg4456} & (~|reg4459)) ^~ "zYzWQl8LMWXsgXag4QY2cWTA"),
                      {(wire4447 >> $signed(wire8)), (-$unsigned(wire8))}} ?
                  "HpX" : reg4461);
            end
        end
    end
  always
    @(posedge clk) begin
      reg4463 <= "RNYs";
    end
  always
    @(posedge clk) begin
      for (forvar4464 = (1'h0); (forvar4464 < (1'h1)); forvar4464 = (forvar4464 + (1'h1)))
        begin
          reg4465 <= wire4449;
          reg4466 <= ((-reg4465[(3'h5):(1'h0)]) ?
              reg4454 : (-(|$unsigned((wire6 ? (7'h4c) : forvar4458)))));
          reg4467 <= (reg4460[(3'h6):(1'h1)] ?
              {reg4465[(3'h4):(1'h0)]} : wire9);
        end
    end
  always
    @(posedge clk) begin
      reg4468 <= $signed($signed(((~^(reg4456 << (7'h44))) ^~ "Bd2hp5yGS5qI5u1Ru5Q")));
      for (forvar4469 = (1'h0); (forvar4469 < (3'h5)); forvar4469 = (forvar4469 + (1'h1)))
        begin
          reg4470 <= reg4461[(5'h10):(4'hc)];
          reg4471 = reg4459;
          reg4472 <= "";
          reg4473 <= wire4449;
          reg4474 <= "Xos9Yxr00dIyVq4CeQNVAXpH";
          reg4475 <= "52cFXnnM1Q9WUsx8";
        end
      reg4476 <= $signed($signed((~|(wire6[(2'h3):(2'h2)] ?
          (reg4456 ? (8'hae) : reg4459) : (wire6 << reg4465)))));
    end
  always
    @(posedge clk) begin
      reg4477 <= ("oTosRE8PR6oQNyIOJJw" ?
          {(+(8'hbf)), (~&("y0" ? $unsigned(reg4455) : reg4476))} : (8'ha6));
      reg4478 <= $signed((({reg4462,
          $unsigned(reg4456)} ^~ $unsigned("NemLvnQZOYOJLcDM0wPDzdc")) - ((&(forvar4464 >= reg4460)) && reg12)));
      reg4479 <= (-(8'hb7));
      for (forvar4480 = (1'h0); (forvar4480 < (3'h4)); forvar4480 = (forvar4480 + (1'h1)))
        begin
          reg4481 <= ((~^reg4475) <<< (({(wire6 ? reg4461 : reg4477),
              wire4453} <<< (-forvar4469)) != (reg16[(4'h8):(1'h0)] | reg4476)));
          reg4482 <= ((|($signed(reg4462) ?
                  "3wnKZ5WkR5" : reg4454[(4'hc):(3'h6)])) ?
              (reg4472 ~^ reg4468) : (8'ha3));
          reg4483 = $signed("Ec3U");
        end
      reg4484 <= ($signed(reg11[(4'h9):(3'h7)]) > forvar4457);
    end
  module3018 modinst4486 (.wire3023(reg4459), .wire3020(reg4479), .wire3019(wire4453), .y(wire4485), .wire3022(reg4454), .wire3021(forvar4457), .clk(clk));
  assign wire4487 = forvar4458[(5'h12):(4'hb)];
  always
    @(posedge clk) begin
      for (forvar4488 = (1'h0); (forvar4488 < (2'h2)); forvar4488 = (forvar4488 + (1'h1)))
        begin
          reg4489 <= {$signed(wire7[(1'h0):(1'h0)]), "2b3X"};
        end
      reg4490 = reg4482;
      reg4491 <= {reg4470,
          ({($signed(reg4479) | (reg4468 <= reg4455)), (&{reg4459})} ?
              reg4456 : $signed(({(8'haa)} || forvar4469[(1'h1):(1'h0)])))};
    end
  assign wire4492 = wire4487[(2'h2):(1'h1)];
  assign wire4493 = $unsigned(((~($signed(reg11) ?
                        (&wire4447) : (reg4476 ?
                            (7'h47) : reg4470))) || (wire9 ^~ ((&reg4461) ?
                        (forvar4457 | forvar4480) : reg4459[(4'ha):(4'ha)]))));
  assign wire4494 = ((reg4482 ?
                        reg13[(4'he):(3'h7)] : "Ez4rzLlqauiBPzE3sBeD84kdY") & (|(("3ZAJXyrOsJVHJS" * wire6) ?
                        (~&forvar4457) : $unsigned("XdOv754tIkemyVGs0A1Qx53Ed"))));
  always
    @(posedge clk) begin
      reg4495 <= reg4491[(1'h1):(1'h1)];
      reg4496 <= $unsigned(wire4447[(4'h9):(4'h9)]);
      reg4497 <= ($unsigned($unsigned(((wire4453 | wire4485) ?
          $signed(forvar4488) : "e4ZJN"))) >>> "uZ9W8cVWdHgh22Ms");
      reg4498 <= (wire10 != reg4478);
      reg4499 = {{forvar4488[(3'h6):(3'h6)]}};
      reg4500 = "wNxavzH";
    end
  always
    @(posedge clk) begin
      reg4501 <= $signed("SyXQRNG5JCimxIxZB5g5eH2n");
      for (forvar4502 = (1'h0); (forvar4502 < (1'h1)); forvar4502 = (forvar4502 + (1'h1)))
        begin
          for (forvar4503 = (1'h0); (forvar4503 < (1'h1)); forvar4503 = (forvar4503 + (1'h1)))
            begin
              for (forvar4504 = (1'h0); (forvar4504 < (2'h3)); forvar4504 = (forvar4504 + (1'h1)))
                begin
                  reg4505 <= $unsigned($signed(forvar4503));
                  reg4506 = $unsigned(((8'ha7) == $unsigned($signed($signed(reg4497)))));
                end
              for (forvar4507 = (1'h0); (forvar4507 < (2'h2)); forvar4507 = (forvar4507 + (1'h1)))
                begin
                  reg4508 <= (+$unsigned((+$unsigned(reg4475))));
                end
              for (forvar4509 = (1'h0); (forvar4509 < (3'h5)); forvar4509 = (forvar4509 + (1'h1)))
                begin
                  reg4510 = (((((reg4475 ?
                          wire4493 : reg4479) >>> reg4459) > (~&reg4466[(3'h4):(3'h4)])) ?
                      (7'h45) : (^~"B")) >= wire4493);
                  reg4511 <= (forvar4480 ?
                      $unsigned(reg4460[(3'h6):(1'h0)]) : reg15[(2'h2):(2'h2)]);
                  reg4512 <= $unsigned(wire7);
                end
              reg4513 = (+reg4471[(2'h2):(1'h1)]);
              reg4514 = ((!reg4491) ^ wire4449[(1'h0):(1'h0)]);
            end
          reg4515 <= reg4473;
          for (forvar4516 = (1'h0); (forvar4516 < (3'h5)); forvar4516 = (forvar4516 + (1'h1)))
            begin
              reg4517 <= (reg4496[(4'hd):(3'h7)] > "BzhJdxzMSc");
              for (forvar4518 = (1'h0); (forvar4518 < (3'h4)); forvar4518 = (forvar4518 + (1'h1)))
                begin
                  reg4519 <= (^{"vby2Th", reg4495});
                  reg4520 <= (reg4456 ?
                      $signed((~|"cGpT")) : $unsigned(wire4451[(3'h5):(3'h5)]));
                  reg4521 = reg4482;
                end
              reg4522 = ((forvar4480[(4'h8):(2'h2)] ?
                  $unsigned(((wire4449 ? reg4479 : wire9) ?
                      (wire4447 ?
                          forvar4480 : reg4491) : $signed(reg4499))) : (~wire4493)) << reg4497);
              reg4523 <= ($unsigned("") ?
                  reg4496[(3'h5):(1'h0)] : ($unsigned((+$signed(wire4494))) * (~|wire4494[(3'h5):(3'h5)])));
              for (forvar4524 = (1'h0); (forvar4524 < (3'h4)); forvar4524 = (forvar4524 + (1'h1)))
                begin
                  reg4525 <= "H1gKknkPaB7RyQ68C9fZUDXp";
                  reg4526 <= (reg4471 ~^ $unsigned($signed("BdbeZUvuBbaubBgJ9emnyiyT")));
                end
              reg4527 <= $unsigned(("oDRlCkzFIzqO8zWBCLgZPsXpS" <<< $signed(((forvar4480 ?
                  wire4494 : wire4453) - (forvar4509 + forvar4507)))));
            end
          for (forvar4528 = (1'h0); (forvar4528 < (2'h2)); forvar4528 = (forvar4528 + (1'h1)))
            begin
              reg4529 = (wire7 ?
                  $signed($unsigned(reg4514)) : reg4489[(5'h10):(2'h2)]);
              reg4530 = "ImtO7RZkpnG9S5OQRrRgnzf08";
              reg4531 <= $signed($unsigned((~&$signed("NGfB4CmgWqO8fic"))));
              reg4532 <= $signed($signed("tv5BKMOsTMQVgdzEOrqQQRzbq"));
              reg4533 <= ((($unsigned($signed(forvar4507)) > reg4517) ?
                  $signed(reg4482) : (reg4505 <= ($unsigned(wire4485) >> $unsigned(wire4494)))) >> ("aZ3m" ?
                  $unsigned(forvar4507[(5'h17):(5'h13)]) : wire7[(4'ha):(3'h4)]));
              reg4534 <= (((~(forvar4504[(4'hf):(3'h5)] ^ "XX26ZF")) ?
                  "kCnTfGWqf22" : reg4505[(4'h9):(4'h9)]) ^ ({(+"1lb"),
                      (-"t946vT5z8tGc43d90F7vZI")} ?
                  $unsigned((^~$signed(forvar4528))) : (reg4474[(2'h2):(1'h0)] - $unsigned(reg4514[(5'h12):(4'hd)]))));
            end
        end
      reg4535 <= $signed($signed({$signed(reg4483)}));
      reg4536 <= "CBGJgq5";
      reg4537 <= reg4484[(5'h13):(4'h8)];
    end
  always
    @(posedge clk) begin
      reg4538 = reg4522[(5'h16):(1'h0)];
      reg4539 <= $signed(($signed($signed((reg4514 <<< wire4485))) ?
          forvar4469[(1'h1):(1'h0)] : $unsigned(("yPvTA" ?
              $unsigned(reg4491) : (reg4466 - wire9)))));
      reg4540 <= ((~&reg4496[(4'h9):(3'h4)]) ?
          {"fq9N9lQp69FiZoQBkX0F"} : "bZ5bUp");
      reg4541 <= $unsigned((8'hb5));
    end
  module93 modinst4543 (wire4542, clk, reg4526, reg4513, reg4490, reg4531);
  always
    @(posedge clk) begin
      reg4544 = "S13W6qoI0V0qEfQyl";
      reg4545 = "zTL";
      for (forvar4546 = (1'h0); (forvar4546 < (1'h0)); forvar4546 = (forvar4546 + (1'h1)))
        begin
          for (forvar4547 = (1'h0); (forvar4547 < (3'h4)); forvar4547 = (forvar4547 + (1'h1)))
            begin
              for (forvar4548 = (1'h0); (forvar4548 < (1'h1)); forvar4548 = (forvar4548 + (1'h1)))
                begin
                  reg4549 = (reg4496 ?
                      (((^reg13) ?
                              forvar4464[(3'h7):(1'h1)] : (reg4497[(3'h7):(3'h4)] ?
                                  $unsigned(wire4453) : (reg4455 + wire8))) ?
                          {reg4477} : reg4455) : ({$signed(reg4527[(1'h0):(1'h0)])} <<< ({(reg4473 >>> reg15)} >> $signed("yHNGm7bbFkske8NVG8s20RlDw"))));
                  reg4550 <= (wire4447 ? reg4476[(4'ha):(3'h7)] : reg4527);
                  reg4551 <= (~"c0nZZEI76C78DlmAq");
                end
              reg4552 <= $unsigned((($unsigned(reg4479) + reg4455[(2'h3):(1'h0)]) | "7W"));
            end
          reg4553 <= reg4462;
          reg4554 <= (!$unsigned((~(~&(reg4466 ? reg4500 : reg4527)))));
        end
      reg4555 = $unsigned($signed(((wire4487 | "d") ?
          $unsigned((^~forvar4502)) : $unsigned(reg4529))));
    end
  assign wire4556 = (((~&(!$signed(forvar4464))) - "ZINdgUf8D") ?
                        reg4476[(3'h5):(1'h1)] : reg4466);
  assign wire4557 = reg4535[(5'h17):(5'h13)];
  always
    @(posedge clk) begin
      for (forvar4558 = (1'h0); (forvar4558 < (3'h4)); forvar4558 = (forvar4558 + (1'h1)))
        begin
          reg4559 = $unsigned(({("4Wecz" >> (~&reg4512)),
                  (forvar4469 * (reg4467 | wire4493))} ?
              $unsigned((8'hae)) : reg4526[(5'h11):(2'h2)]));
          for (forvar4560 = (1'h0); (forvar4560 < (3'h5)); forvar4560 = (forvar4560 + (1'h1)))
            begin
              reg4561 = (8'hb4);
              reg4562 <= {($signed(reg4460[(1'h1):(1'h1)]) ?
                      (reg4466 ^~ (reg11 ?
                          "LnHRHhGNUnpeB4bHgifaB" : $unsigned(reg4455))) : ((~forvar4504[(1'h1):(1'h0)]) ?
                          {reg4481} : (reg4527[(1'h0):(1'h0)] || forvar4509[(1'h1):(1'h0)]))),
                  ("i" ? reg4539[(4'h8):(3'h4)] : wire4453)};
              reg4563 = $unsigned((-(reg4491[(1'h0):(1'h0)] ?
                  $unsigned($signed(reg4519)) : (+(reg4466 ?
                      wire4453 : reg4500)))));
            end
          reg4564 = "2OWELipKZaUplC";
        end
      for (forvar4565 = (1'h0); (forvar4565 < (1'h0)); forvar4565 = (forvar4565 + (1'h1)))
        begin
          reg4566 = (!reg4499[(3'h5):(1'h1)]);
          reg4567 <= $unsigned((8'hbf));
          reg4568 <= reg4489;
        end
    end
  assign wire4569 = $signed(((+reg4567) ?
                        reg4531[(4'he):(4'he)] : $signed($unsigned($unsigned((8'ha0))))));
  always
    @(posedge clk) begin
      reg4570 <= (~(reg4567 ?
          {reg13[(3'h5):(1'h0)],
              reg4545[(4'h9):(1'h0)]} : forvar4558[(5'h10):(3'h5)]));
      reg4571 <= ((((reg13 && reg4550) ?
              reg4495[(4'ha):(2'h2)] : (&forvar4560[(2'h3):(1'h0)])) && ((|$signed(reg4495)) ?
              reg4460 : $signed((~reg4521)))) ?
          {$signed(("9" << "3TQd0MCAD0evuqA77B5qz")),
              {{"HMiKsZ9Zs0ZBHf7o83pJzm5", $signed(reg4537)},
                  wire9}} : (reg4549 >>> $signed((~((8'haf) ?
              (8'ha8) : reg4521)))));
      reg4572 <= ((((7'h4a) ~^ ((8'ha4) ?
              $signed(reg4529) : $unsigned((8'ha1)))) ?
          reg4455[(5'h11):(4'h9)] : (((8'haf) ?
              $unsigned(reg4533) : "Ftw2nzFpqBwseCAFA") >>> reg4530[(5'h10):(3'h6)])) == ("f3eL3VTyKsxk4LJ72Pr" != $signed((7'h4b))));
      reg4573 <= (|"nlPP");
      reg4574 <= ((+$signed($signed(reg13[(1'h1):(1'h1)]))) ?
          ($unsigned($signed((wire4449 >> reg4501))) ?
              (8'hac) : $signed("0WewNaZd4upo2qN64wS5TKg")) : (($unsigned((^(8'hb0))) ?
                  "23MvJ" : $signed((reg4521 ? reg4483 : wire4487))) ?
              "bWEUJPO3bZOPghp5d" : ((&(forvar4464 != wire4487)) ?
                  wire4449[(1'h0):(1'h0)] : ((~&(8'had)) ?
                      (forvar4458 <= (8'ha0)) : reg4461[(5'h15):(4'hf)]))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module17
#( parameter param4445 = {(({{(7'h49), (7'h42)}, (~|(7'h46))} >>> (((7'h4c) ^~ (8'hb1)) | {(8'hbd), (7'h40)})) ? (!(((8'hae) ? (8'ha1) : (7'h42)) | {(7'h46), (8'hb6)})) : ({(7'h49)} ~^ (~^((8'hba) ? (8'hb8) : (7'h41)))))}
, parameter param4446 = param4445 )
(y, clk, wire22, wire21, wire20, wire19, wire18);
  output wire [(32'h3fc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire22;
  input wire signed [(5'h18):(1'h0)] wire21;
  input wire signed [(4'h9):(1'h0)] wire20;
  input wire signed [(5'h18):(1'h0)] wire19;
  input wire signed [(5'h1a):(1'h0)] wire18;
  reg signed [(2'h2):(1'h0)] reg4444 = (1'h0);
  reg [(5'h17):(1'h0)] reg4443 = (1'h0);
  reg [(5'h12):(1'h0)] reg4442 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4441 = (1'h0);
  wire [(5'h14):(1'h0)] wire4439;
  wire [(5'h12):(1'h0)] wire4426;
  reg signed [(5'h12):(1'h0)] reg4425 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg4424 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4423 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg4422 = (1'h0);
  reg [(5'h11):(1'h0)] reg4421 = (1'h0);
  wire signed [(5'h16):(1'h0)] wire4420;
  wire [(5'h18):(1'h0)] wire4418;
  reg signed [(5'h11):(1'h0)] reg4417 = (1'h0);
  reg [(5'h15):(1'h0)] reg4416 = (1'h0);
  reg [(4'hc):(1'h0)] reg4415 = (1'h0);
  reg [(3'h7):(1'h0)] reg4414 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4413 = (1'h0);
  wire [(5'h12):(1'h0)] wire4404;
  reg signed [(4'hc):(1'h0)] reg52 = (1'h0);
  reg [(4'he):(1'h0)] reg51 = (1'h0);
  reg [(5'h1a):(1'h0)] reg50 = (1'h0);
  reg [(5'h1a):(1'h0)] reg49 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar48 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg47 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg46 = (1'h0);
  reg [(4'ha):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar44 = (1'h0);
  reg [(5'h13):(1'h0)] reg43 = (1'h0);
  reg [(5'h10):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg41 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar40 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg39 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg38 = (1'h0);
  reg [(3'h5):(1'h0)] reg37 = (1'h0);
  reg signed [(4'he):(1'h0)] reg36 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg35 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg34 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg33 = (1'h0);
  reg [(5'h18):(1'h0)] forvar32 = (1'h0);
  reg [(5'h17):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg29 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg28 = (1'h0);
  reg [(5'h19):(1'h0)] reg27 = (1'h0);
  reg [(5'h17):(1'h0)] reg26 = (1'h0);
  reg [(5'h18):(1'h0)] reg25 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar24 = (1'h0);
  wire [(5'h12):(1'h0)] wire23;
  wire [(3'h5):(1'h0)] wire4406;
  wire [(5'h19):(1'h0)] wire4408;
  reg [(4'h8):(1'h0)] reg4410 = (1'h0);
  wire [(5'h18):(1'h0)] wire4411;
  reg signed [(5'h14):(1'h0)] reg4428 = (1'h0);
  reg [(5'h14):(1'h0)] reg4429 = (1'h0);
  reg [(5'h19):(1'h0)] forvar4430 = (1'h0);
  reg [(5'h12):(1'h0)] reg4431 = (1'h0);
  reg [(4'hf):(1'h0)] reg4432 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg4433 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4434 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire4435;
  wire [(5'h11):(1'h0)] wire4437;
  assign y = {reg4444,
                 reg4443,
                 reg4442,
                 reg4441,
                 wire4439,
                 wire4426,
                 reg4425,
                 reg4424,
                 forvar4423,
                 reg4422,
                 reg4421,
                 wire4420,
                 wire4418,
                 reg4417,
                 reg4416,
                 reg4415,
                 reg4414,
                 reg4413,
                 wire4404,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 forvar48,
                 reg47,
                 reg46,
                 reg45,
                 forvar44,
                 reg43,
                 reg42,
                 reg41,
                 forvar40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 forvar32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 forvar24,
                 wire23,
                 wire4406,
                 wire4408,
                 reg4410,
                 wire4411,
                 reg4428,
                 reg4429,
                 forvar4430,
                 reg4431,
                 reg4432,
                 reg4433,
                 reg4434,
                 wire4435,
                 wire4437,
                 (1'h0)};
  assign wire23 = (8'h9e);
  always
    @(posedge clk) begin
      for (forvar24 = (1'h0); (forvar24 < (1'h1)); forvar24 = (forvar24 + (1'h1)))
        begin
          reg25 = wire22;
          reg26 = "p4iEH60dyUfo9HYfS";
        end
      reg27 <= (wire23[(2'h2):(1'h1)] ?
          {({$signed(wire22), $unsigned(wire19)} ?
                  $signed((+wire20)) : $signed((^~forvar24)))} : $signed(($unsigned(((8'ha4) ?
                  wire19 : wire23)) ?
              $unsigned($unsigned(wire20)) : (^wire18))));
      reg28 <= wire23[(4'h8):(1'h1)];
      reg29 <= (!reg28[(1'h1):(1'h0)]);
      reg30 <= "ZQTRBgZL";
    end
  always
    @(posedge clk) begin
      reg31 <= ((7'h4d) ? (8'hb7) : reg30);
      for (forvar32 = (1'h0); (forvar32 < (3'h5)); forvar32 = (forvar32 + (1'h1)))
        begin
          if (forvar32[(3'h7):(1'h1)])
            begin
              reg33 <= $unsigned((8'hb1));
            end
          else
            begin
              reg33 = $unsigned("SpSCuYkezcLzN");
              reg34 = {(reg25[(1'h1):(1'h1)] ? wire18 : $signed(reg33))};
              reg35 <= $unsigned(("dMWUY1lJ6paB" ?
                  (({reg31} | (wire18 ? reg27 : forvar32)) ?
                      reg27[(3'h5):(1'h0)] : ({reg25} || $unsigned(wire19))) : forvar32[(3'h7):(3'h6)]));
              reg36 = $signed(($unsigned(reg34[(1'h0):(1'h0)]) | $unsigned(((reg27 ?
                      wire19 : reg33) ?
                  $unsigned(reg33) : (^~wire21)))));
              reg37 <= (($unsigned($signed($unsigned(wire19))) <= "T") >>> $signed(((((7'h4e) + reg25) ?
                      wire18 : wire18[(3'h5):(2'h2)]) ?
                  (reg31 | forvar32[(3'h5):(2'h3)]) : reg36[(3'h6):(3'h4)])));
              reg38 = ($unsigned({"Vq"}) | wire18[(2'h3):(1'h0)]);
            end
          reg39 <= "uP5rh9w";
          for (forvar40 = (1'h0); (forvar40 < (2'h2)); forvar40 = (forvar40 + (1'h1)))
            begin
              reg41 <= ($signed((~&reg38[(1'h0):(1'h0)])) > reg37[(1'h0):(1'h0)]);
              reg42 <= (~|reg26);
              reg43 = $unsigned((8'ha6));
            end
          for (forvar44 = (1'h0); (forvar44 < (1'h1)); forvar44 = (forvar44 + (1'h1)))
            begin
              reg45 <= "8FcXVl8hbbhtud";
              reg46 <= (~|wire21[(4'hc):(3'h7)]);
              reg47 <= (~&{(~&$unsigned((~|reg30))), (~"lzU83XkzsT")});
              for (forvar48 = (1'h0); (forvar48 < (1'h1)); forvar48 = (forvar48 + (1'h1)))
                begin
                  reg49 <= (~((~{(&reg34)}) ?
                      (~((|reg46) ^ {wire23,
                          reg36})) : $signed($signed(reg45))));
                  reg50 <= (-(reg30 ?
                      (wire20 >= "PHdg2KkmqRlMKcoNW") : (7'h44)));
                  reg51 = reg34;
                end
              reg52 <= $signed($signed(("SGbT" >= $signed((reg46 ?
                  wire20 : wire18)))));
            end
        end
    end
  module53 modinst4405 (wire4404, clk, reg49, wire19, reg31, reg30, reg28);
  module2781 modinst4407 (.y(wire4406), .wire2782(forvar44), .wire2783(reg25), .wire2785(forvar32), .clk(clk), .wire2784(reg49));
  module4117 modinst4409 (.wire4121(reg45), .clk(clk), .wire4119(reg43), .wire4118(reg27), .wire4120(wire21), .y(wire4408));
  always
    @(posedge clk) begin
      reg4410 <= "";
    end
  module2282 modinst4412 (wire4411, clk, reg46, wire22, reg33, reg36, reg34);
  always
    @(posedge clk) begin
      reg4413 <= (&wire4411);
      reg4414 <= wire4406[(2'h3):(2'h2)];
      reg4415 = (reg47[(3'h7):(3'h5)] ?
          (~&(~&({reg35} && ((7'h48) ?
              reg49 : (8'hbc))))) : reg36[(1'h1):(1'h0)]);
      reg4416 <= {{$unsigned($unsigned((~|(8'ha4)))),
              (((^(7'h47)) ? (wire23 ^ (8'ha8)) : reg25[(2'h3):(1'h1)]) ?
                  reg36[(4'hc):(2'h2)] : (^~(reg39 ? reg27 : forvar48)))},
          reg41};
      reg4417 = ($signed(reg45[(1'h1):(1'h1)]) ? "" : forvar44);
    end
  module219 modinst4419 (.clk(clk), .wire221(reg30), .wire223(reg41), .wire222(wire19), .y(wire4418), .wire220(reg42));
  assign wire4420 = $signed((&((((8'hbd) ? reg4416 : reg4413) << (~&reg34)) ?
                        reg30 : (~&forvar24))));
  always
    @(posedge clk) begin
      reg4421 <= ((|reg26[(3'h7):(1'h1)]) ?
          reg4414[(3'h6):(2'h2)] : "ELRJ5i8qk06RpHvR2kP");
      reg4422 <= ($unsigned(((+reg4413[(2'h3):(1'h1)]) ?
          ((&reg25) ? "ECuw" : $signed(reg4410)) : {reg27[(4'h9):(1'h1)],
              (reg4415 ?
                  reg52 : reg41)})) | ($signed(($unsigned(wire4420) * (~&reg31))) | reg50));
      for (forvar4423 = (1'h0); (forvar4423 < (2'h2)); forvar4423 = (forvar4423 + (1'h1)))
        begin
          reg4424 = (($unsigned((~(reg51 ?
                  (8'hbc) : (8'ha9)))) >> ((8'ha9) << (~^wire21[(4'ha):(3'h5)]))) ?
              reg33 : $signed((forvar48 ? reg31 : "1E78pvDYJ5RGFoXPGJpd")));
        end
      reg4425 <= ($signed($unsigned(wire4420)) >> "d");
    end
  module3696 modinst4427 (wire4426, clk, reg26, reg50, reg27, wire18, reg39);
  always
    @(posedge clk) begin
      reg4428 <= reg41;
      reg4429 <= (7'h45);
      for (forvar4430 = (1'h0); (forvar4430 < (1'h0)); forvar4430 = (forvar4430 + (1'h1)))
        begin
          reg4431 <= $signed($unsigned(({(~^reg28), wire21[(4'hc):(1'h1)]} ?
              reg36[(4'hc):(3'h7)] : wire20)));
          reg4432 <= $signed(wire4418);
        end
      reg4433 = $unsigned(({{$signed(reg33), $signed(wire22)}} ?
          (reg31[(5'h13):(4'hd)] == {$unsigned(forvar32),
              $unsigned((7'h41))}) : $unsigned({$signed(reg4429)})));
      reg4434 <= "1I4yZcmZTLV0x0XMWUsHdU";
    end
  module1013 modinst4436 (wire4435, clk, reg4425, reg4424, reg4416, forvar32);
  module2841 modinst4438 (wire4437, clk, wire4420, reg4410, reg29, reg50, reg4417);
  module3981 modinst4440 (wire4439, clk, wire22, reg45, reg4431, reg49);
  always
    @(posedge clk) begin
      reg4441 = (reg30[(5'h15):(4'hc)] ?
          reg52[(4'h8):(3'h6)] : ("F2ZPIbzlWhvlWOS4" || (((forvar44 ?
              wire4408 : reg51) != ((7'h4e) ? reg4421 : reg47)) != (((8'ha5) ?
                  reg41 : reg4410) ?
              (reg35 | (8'ha2)) : reg46[(2'h3):(2'h3)]))));
      reg4442 <= $unsigned($signed({forvar4423[(1'h0):(1'h0)]}));
      reg4443 <= reg4414;
      reg4444 <= ((~^reg4433) ?
          {(+wire4426)} : (reg26[(4'hc):(2'h2)] ?
              "pp" : ({(wire4411 << forvar40), (wire23 ? wire4418 : reg27)} ?
                  {forvar4430[(2'h3):(1'h1)],
                      wire4411} : reg35[(3'h4):(1'h1)])));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module53
#( parameter param4403 = (({(((8'ha6) ^~ (7'h45)) + ((8'hb9) ? (8'ha0) : (7'h4e)))} == (({(7'h4b)} ? (8'hb4) : (8'ha9)) ? (((7'h45) << (8'h9e)) & ((8'hb2) || (8'ha8))) : ((8'hae) ? {(7'h4e), (8'hbd)} : ((7'h41) ? (8'hbc) : (8'hb6))))) ? ((^(7'h48)) ? (({(8'ha8), (7'h44)} >= ((8'ha4) >> (8'ha3))) ? ({(7'h4d)} || {(7'h45)}) : (-(8'h9c))) : (!(~((8'hac) | (8'h9f))))) : {(7'h41)}) )
(y, clk, wire54, wire55, wire56, wire57, wire58);
  output wire [(32'h6c3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h1a):(1'h0)] wire54;
  input wire signed [(5'h18):(1'h0)] wire55;
  input wire signed [(5'h17):(1'h0)] wire56;
  input wire signed [(5'h16):(1'h0)] wire57;
  input wire [(5'h1a):(1'h0)] wire58;
  wire [(3'h5):(1'h0)] wire4402;
  wire signed [(5'h13):(1'h0)] wire4401;
  reg [(5'h15):(1'h0)] reg4400 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4399 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg4398 = (1'h0);
  reg [(2'h3):(1'h0)] reg4397 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4396 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg4395 = (1'h0);
  reg [(4'hf):(1'h0)] reg4394 = (1'h0);
  reg [(5'h14):(1'h0)] reg4393 = (1'h0);
  reg [(5'h11):(1'h0)] forvar4392 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4391 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4390 = (1'h0);
  reg [(5'h18):(1'h0)] reg4389 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4388 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4387 = (1'h0);
  reg [(4'h9):(1'h0)] reg4386 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4385 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg4384 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire4383;
  reg [(3'h7):(1'h0)] reg4382 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4376 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4375 = (1'h0);
  reg [(4'h8):(1'h0)] reg4374 = (1'h0);
  reg [(5'h16):(1'h0)] reg4381 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4380 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4379 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4378 = (1'h0);
  reg [(3'h6):(1'h0)] reg4377 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar4376 = (1'h0);
  reg [(3'h7):(1'h0)] reg4375 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4374 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4373 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg4372 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4371 = (1'h0);
  reg [(5'h10):(1'h0)] reg4370 = (1'h0);
  wire [(5'h13):(1'h0)] wire4368;
  wire [(5'h18):(1'h0)] wire4366;
  wire signed [(4'h8):(1'h0)] wire4357;
  reg [(3'h4):(1'h0)] reg4356 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg4355 = (1'h0);
  reg [(4'h8):(1'h0)] reg4354 = (1'h0);
  reg [(5'h1a):(1'h0)] reg4353 = (1'h0);
  reg [(4'ha):(1'h0)] reg4352 = (1'h0);
  reg [(5'h18):(1'h0)] reg4351 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4350 = (1'h0);
  reg [(5'h13):(1'h0)] reg4349 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg4348 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4347 = (1'h0);
  reg [(4'h9):(1'h0)] reg4346 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar4345 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg4344 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar4343 = (1'h0);
  reg [(5'h11):(1'h0)] reg4342 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4341 = (1'h0);
  reg [(5'h10):(1'h0)] reg4340 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4339 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4338 = (1'h0);
  reg [(4'he):(1'h0)] forvar4337 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg4336 = (1'h0);
  reg [(5'h13):(1'h0)] reg4335 = (1'h0);
  reg [(3'h4):(1'h0)] reg4334 = (1'h0);
  reg [(5'h18):(1'h0)] reg4333 = (1'h0);
  reg [(5'h1a):(1'h0)] reg4332 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4331 = (1'h0);
  reg [(5'h11):(1'h0)] reg4330 = (1'h0);
  reg [(5'h18):(1'h0)] reg4329 = (1'h0);
  reg [(5'h15):(1'h0)] reg4328 = (1'h0);
  reg [(5'h19):(1'h0)] reg4327 = (1'h0);
  reg [(3'h6):(1'h0)] reg4326 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4325 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4324 = (1'h0);
  reg [(4'h9):(1'h0)] reg4323 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4322 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4321 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4320 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg4319 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4318 = (1'h0);
  wire [(4'h8):(1'h0)] wire4317;
  wire signed [(4'hd):(1'h0)] wire4316;
  wire signed [(5'h10):(1'h0)] wire4315;
  reg signed [(5'h15):(1'h0)] reg4314 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg4313 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg4312 = (1'h0);
  reg [(5'h11):(1'h0)] reg4311 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4310 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4309 = (1'h0);
  wire [(5'h19):(1'h0)] wire4308;
  reg signed [(5'h1a):(1'h0)] reg4307 = (1'h0);
  reg [(5'h12):(1'h0)] forvar4306 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4305 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar4304 = (1'h0);
  reg [(4'h9):(1'h0)] reg4303 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4302 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4301 = (1'h0);
  reg [(4'he):(1'h0)] forvar4300 = (1'h0);
  reg [(3'h7):(1'h0)] reg4299 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4298 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar4297 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar4296 = (1'h0);
  reg [(5'h11):(1'h0)] reg4295 = (1'h0);
  reg [(3'h5):(1'h0)] reg4294 = (1'h0);
  reg [(4'hc):(1'h0)] reg59 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar60 = (1'h0);
  reg signed [(4'he):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg62 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg63 = (1'h0);
  reg [(5'h16):(1'h0)] reg64 = (1'h0);
  reg [(5'h19):(1'h0)] reg65 = (1'h0);
  reg [(5'h13):(1'h0)] reg66 = (1'h0);
  reg [(4'h8):(1'h0)] reg67 = (1'h0);
  reg [(5'h11):(1'h0)] reg68 = (1'h0);
  reg [(4'hc):(1'h0)] reg69 = (1'h0);
  wire [(2'h2):(1'h0)] wire4292;
  reg signed [(5'h12):(1'h0)] reg4359 = (1'h0);
  reg [(4'h8):(1'h0)] reg4360 = (1'h0);
  reg [(5'h17):(1'h0)] reg4361 = (1'h0);
  reg [(4'ha):(1'h0)] reg4362 = (1'h0);
  reg [(5'h12):(1'h0)] reg4363 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire4364;
  assign y = {wire4402,
                 wire4401,
                 reg4400,
                 reg4399,
                 reg4398,
                 reg4397,
                 reg4396,
                 reg4395,
                 reg4394,
                 reg4393,
                 forvar4392,
                 reg4391,
                 forvar4390,
                 reg4389,
                 forvar4388,
                 reg4387,
                 reg4386,
                 forvar4385,
                 reg4384,
                 wire4383,
                 reg4382,
                 reg4376,
                 forvar4375,
                 reg4374,
                 reg4381,
                 reg4380,
                 reg4379,
                 reg4378,
                 reg4377,
                 forvar4376,
                 reg4375,
                 forvar4374,
                 reg4373,
                 reg4372,
                 forvar4371,
                 reg4370,
                 wire4368,
                 wire4366,
                 wire4357,
                 reg4356,
                 reg4355,
                 reg4354,
                 reg4353,
                 reg4352,
                 reg4351,
                 forvar4350,
                 reg4349,
                 reg4348,
                 reg4347,
                 reg4346,
                 forvar4345,
                 reg4344,
                 forvar4343,
                 reg4342,
                 reg4341,
                 reg4340,
                 reg4339,
                 reg4338,
                 forvar4337,
                 reg4336,
                 reg4335,
                 reg4334,
                 reg4333,
                 reg4332,
                 forvar4331,
                 reg4330,
                 reg4329,
                 reg4328,
                 reg4327,
                 reg4326,
                 reg4325,
                 forvar4324,
                 reg4323,
                 forvar4322,
                 reg4321,
                 reg4320,
                 reg4319,
                 forvar4318,
                 wire4317,
                 wire4316,
                 wire4315,
                 reg4314,
                 reg4313,
                 reg4312,
                 reg4311,
                 reg4310,
                 reg4309,
                 wire4308,
                 reg4307,
                 forvar4306,
                 reg4305,
                 forvar4304,
                 reg4303,
                 reg4302,
                 reg4301,
                 forvar4300,
                 reg4299,
                 reg4298,
                 forvar4297,
                 forvar4296,
                 reg4295,
                 reg4294,
                 reg59,
                 forvar60,
                 reg61,
                 reg62,
                 reg63,
                 reg64,
                 reg65,
                 reg66,
                 reg67,
                 reg68,
                 reg69,
                 wire4292,
                 reg4359,
                 reg4360,
                 reg4361,
                 reg4362,
                 reg4363,
                 wire4364,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg59 <= (|(($unsigned($signed(wire58)) ^~ $signed((wire56 ?
              wire58 : wire54))) ?
          "w0gXXf8SUwZz3vdD5Bdp" : (&wire56[(5'h12):(4'hb)])));
      for (forvar60 = (1'h0); (forvar60 < (2'h2)); forvar60 = (forvar60 + (1'h1)))
        begin
          reg61 = forvar60[(2'h2):(2'h2)];
          reg62 <= wire54;
          reg63 <= "3aDxZ3";
          reg64 <= {$signed("nT8oiAfuSUFbfHALL"), wire56[(5'h11):(3'h6)]};
        end
    end
  always
    @(posedge clk) begin
      reg65 <= (^$unsigned((~((reg63 <= (8'hb5)) << $unsigned(wire57)))));
      reg66 <= {"TuHnUP", "gNLWQZdNh5mkcCwrd3"};
      reg67 <= ((({(wire54 & reg65), "mYB2"} ?
          (forvar60 >= (reg64 ? wire56 : reg59)) : reg63) ~^ "") == reg64);
    end
  always
    @(posedge clk) begin
      reg68 <= (!($unsigned((^~reg61)) <= "8tYhpW7BCks4yW5WXzTv2"));
      reg69 <= $unsigned(($signed($signed((~&wire58))) ?
          reg67 : reg62[(4'ha):(3'h5)]));
    end
  module70 modinst4293 (.wire74(wire58), .clk(clk), .wire73(wire54), .wire75(reg64), .wire72(wire55), .wire71(reg67), .y(wire4292));
  always
    @(posedge clk) begin
      reg4294 <= reg69[(3'h5):(3'h5)];
      reg4295 <= (8'ha1);
      for (forvar4296 = (1'h0); (forvar4296 < (1'h1)); forvar4296 = (forvar4296 + (1'h1)))
        begin
          for (forvar4297 = (1'h0); (forvar4297 < (3'h5)); forvar4297 = (forvar4297 + (1'h1)))
            begin
              reg4298 = $unsigned($signed(($signed((forvar4296 >> reg68)) ?
                  (~|wire55) : reg4295[(3'h6):(2'h3)])));
              reg4299 = wire55[(4'h8):(3'h4)];
            end
          for (forvar4300 = (1'h0); (forvar4300 < (3'h4)); forvar4300 = (forvar4300 + (1'h1)))
            begin
              reg4301 <= (forvar60 ?
                  ({$signed($signed(reg4299))} ?
                      wire4292 : (~&(reg63 ?
                          reg63[(1'h0):(1'h0)] : (~^reg4294)))) : $unsigned(($unsigned((wire55 <<< forvar4296)) ^ (~^$unsigned((8'hb0))))));
            end
          reg4302 <= (("mKkysfHLJ6flVb" != $signed("Z95rcGZQL")) > wire57[(3'h4):(2'h2)]);
          reg4303 <= "gvzqT82OU";
        end
      for (forvar4304 = (1'h0); (forvar4304 < (3'h5)); forvar4304 = (forvar4304 + (1'h1)))
        begin
          reg4305 <= "w2KGHI7MP";
        end
      for (forvar4306 = (1'h0); (forvar4306 < (2'h3)); forvar4306 = (forvar4306 + (1'h1)))
        begin
          reg4307 <= {reg69[(2'h3):(1'h0)], forvar4306[(1'h0):(1'h0)]};
        end
    end
  assign wire4308 = wire57[(3'h4):(1'h0)];
  always
    @(posedge clk) begin
      reg4309 <= (^$unsigned((reg4301 ?
          reg67[(1'h0):(1'h0)] : (-$unsigned((8'haf))))));
      reg4310 = (reg67[(1'h0):(1'h0)] ? forvar4306 : "C");
      reg4311 <= $unsigned(reg63[(1'h1):(1'h1)]);
      reg4312 <= $unsigned((^$unsigned(reg4299[(3'h7):(3'h7)])));
      reg4313 <= reg4311;
      reg4314 <= {$signed((wire55[(5'h11):(3'h6)] >= $unsigned($signed(reg69)))),
          ("MGbmW3mi8vP" >= ($signed((reg4294 ? reg64 : reg4294)) ?
              {(forvar4304 <<< reg4295)} : reg65))};
    end
  assign wire4315 = "mk8piRSpvBwJ7kE8PqKxv";
  assign wire4316 = (("kxNwrbDhQ4oJiYSUWS1a2Q" ?
                        forvar4304[(5'h12):(5'h10)] : $unsigned(reg69)) >= reg65);
  assign wire4317 = (8'hb3);
  always
    @(posedge clk) begin
      for (forvar4318 = (1'h0); (forvar4318 < (3'h5)); forvar4318 = (forvar4318 + (1'h1)))
        begin
          reg4319 <= wire57;
          reg4320 <= wire54[(4'hd):(4'hb)];
          reg4321 = $unsigned("lVutu0IqlP8CtyYVxZQ");
          for (forvar4322 = (1'h0); (forvar4322 < (1'h0)); forvar4322 = (forvar4322 + (1'h1)))
            begin
              reg4323 <= ($signed(({$unsigned(reg4313),
                      (reg4321 >= forvar4318)} && $unsigned($signed(wire4317)))) ?
                  $unsigned(forvar4306) : (reg4311[(4'hc):(3'h5)] ?
                      $unsigned($signed(wire4317)) : (((reg4314 ^~ (7'h4e)) ?
                          (reg4301 ? forvar4304 : reg4313) : (reg61 ?
                              (8'ha2) : wire55)) != reg68)));
              for (forvar4324 = (1'h0); (forvar4324 < (1'h1)); forvar4324 = (forvar4324 + (1'h1)))
                begin
                  reg4325 = $unsigned($signed($signed(wire58)));
                  reg4326 <= "h8I1GGJYktUd";
                  reg4327 = $unsigned($signed("vyuR9E9Nd0tPO4WbRDu"));
                  reg4328 <= (!"W6VCSKPcLbMLLdLT");
                  reg4329 <= "Q";
                end
              reg4330 <= reg4302;
              for (forvar4331 = (1'h0); (forvar4331 < (1'h0)); forvar4331 = (forvar4331 + (1'h1)))
                begin
                  reg4332 <= $unsigned(forvar4300[(4'h8):(3'h6)]);
                  reg4333 <= (reg4328[(5'h15):(4'he)] ?
                      (~^(&((reg69 ? forvar4300 : reg4326) ?
                          "lRotBGfsEsCht7IccFgB" : $signed(reg4320)))) : reg4303);
                  reg4334 <= (~reg4320[(3'h4):(1'h0)]);
                  reg4335 = reg69[(4'h8):(2'h3)];
                  reg4336 = reg4334;
                end
              for (forvar4337 = (1'h0); (forvar4337 < (3'h5)); forvar4337 = (forvar4337 + (1'h1)))
                begin
                  reg4338 <= $unsigned(($unsigned("oicLHGqMShmGcfHlffNeF") ?
                      (|"DcgXhqCuZPgk") : $unsigned(({reg4334, wire54} ?
                          (forvar4297 <<< reg4327) : (^reg4299)))));
                  reg4339 <= ("teYWFV" ?
                      $signed($unsigned($signed($signed(reg4334)))) : (~$signed((~^(reg64 || reg4319)))));
                  reg4340 = (&forvar4296);
                  reg4341 = "UpBfBBYESW16Dz0um2kwc";
                end
              reg4342 <= $unsigned($signed((reg4338[(4'hc):(2'h3)] & (wire58 ?
                  (wire58 ? wire56 : wire4315) : (reg4305 ?
                      forvar4318 : wire55)))));
            end
        end
      for (forvar4343 = (1'h0); (forvar4343 < (3'h5)); forvar4343 = (forvar4343 + (1'h1)))
        begin
          reg4344 <= forvar4318[(1'h0):(1'h0)];
          for (forvar4345 = (1'h0); (forvar4345 < (2'h2)); forvar4345 = (forvar4345 + (1'h1)))
            begin
              reg4346 <= reg4321;
              reg4347 = ("nBtCXO" ?
                  ((|"C8PbcHNR6veB") ?
                      (~^$signed($signed(reg4321))) : ($signed((+reg4299)) ?
                          ($signed((8'hb3)) ~^ {(7'h40)}) : (~|((7'h4c) >> (8'hb6))))) : (|{reg4333}));
              reg4348 <= forvar4331;
              reg4349 = $signed($unsigned($signed(forvar4296)));
            end
          for (forvar4350 = (1'h0); (forvar4350 < (3'h4)); forvar4350 = (forvar4350 + (1'h1)))
            begin
              reg4351 = forvar4324;
              reg4352 <= $signed(($unsigned("J") ?
                  (reg4309 != wire4308[(5'h10):(4'he)]) : reg4320));
              reg4353 <= reg4352;
            end
        end
      reg4354 <= ((("8TLesoff6v79EQ7Hn73MIb" ?
              (reg4310[(1'h1):(1'h1)] >= (~^forvar4345)) : (8'hb0)) ?
          forvar4324 : $signed($unsigned($signed(forvar4345)))) | reg64);
      reg4355 <= (~^$unsigned($unsigned(({(8'hb3)} ?
          ((8'hae) ? wire56 : reg4330) : reg4351))));
      reg4356 = ($unsigned(({{reg4354}} & $unsigned($signed(reg4349)))) ?
          $signed(reg4320[(3'h7):(3'h6)]) : {"8WMos"});
    end
  module79 modinst4358 (wire4357, clk, reg4353, forvar4343, reg4348, forvar4306, forvar4296);
  always
    @(posedge clk) begin
      reg4359 <= wire55[(4'hd):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg4360 <= (^~$unsigned($signed("F1B4VOc")));
      reg4361 <= (~((~^reg4294) ?
          "fTwZdTQyEW" : ({$signed(reg4355), {(8'haf)}} ?
              $unsigned("Pag3HNDkki6wiBAvB9x4RpkC9") : reg4321[(3'h5):(3'h5)])));
      reg4362 = {(8'ha5)};
      reg4363 <= reg4347[(1'h1):(1'h1)];
    end
  module2841 modinst4365 (wire4364, clk, reg4321, reg4329, wire57, reg4332, reg4314);
  module1250 modinst4367 (wire4366, clk, reg4311, reg65, forvar4322, reg4362);
  module1250 modinst4369 (.clk(clk), .wire1251(reg4353), .wire1252(reg62), .y(wire4368), .wire1253(reg66), .wire1254(wire4315));
  always
    @(posedge clk) begin
      reg4370 <= ("CCg" * reg4362[(4'h8):(3'h5)]);
      for (forvar4371 = (1'h0); (forvar4371 < (1'h1)); forvar4371 = (forvar4371 + (1'h1)))
        begin
          reg4372 <= ("PUQHPvK3" ? reg67[(3'h7):(3'h7)] : "RWzcNwio");
        end
      reg4373 = reg4332;
    end
  always
    @(posedge clk) begin
      if ($signed((((((8'hbd) ? (7'h4a) : reg4349) < (reg4349 * reg4320)) ?
              ($unsigned((8'hac)) < reg4344[(2'h3):(1'h0)]) : $unsigned($signed(reg4310))) ?
          (&$unsigned((reg4314 ?
              wire55 : (8'ha2)))) : $unsigned($signed((reg4328 ^~ (8'hb1)))))))
        begin
          for (forvar4374 = (1'h0); (forvar4374 < (3'h5)); forvar4374 = (forvar4374 + (1'h1)))
            begin
              reg4375 <= (&$signed($signed(forvar4322[(3'h5):(1'h0)])));
            end
          for (forvar4376 = (1'h0); (forvar4376 < (1'h1)); forvar4376 = (forvar4376 + (1'h1)))
            begin
              reg4377 <= ((~|(({wire4317, reg64} ~^ {reg4319, reg4360}) ?
                      (^"Qqq0V") : $unsigned((forvar60 & (8'h9c))))) ?
                  $signed(wire55) : {"2NZ0XlfwZl1Pxe5a9JC0"});
              reg4378 = forvar4306;
              reg4379 <= (~|$signed(("k1cWX" >> $unsigned((reg66 >> reg4320)))));
            end
          reg4380 <= reg4328;
          reg4381 <= "JQCUi6cgL0r918ZxNMgJD";
        end
      else
        begin
          reg4374 <= (~|wire54[(5'h13):(3'h5)]);
          for (forvar4375 = (1'h0); (forvar4375 < (1'h0)); forvar4375 = (forvar4375 + (1'h1)))
            begin
              reg4376 <= (forvar4296 != "ozl6xfDNn6T2gtd1L3nFT");
              reg4377 <= "iEqK2zD7QtOsMUCiy";
              reg4378 <= wire4357;
              reg4379 <= "83R4CVbiScdOGRBmPm33";
            end
          reg4380 <= (reg4319[(5'h13):(1'h0)] ?
              "lgrOz4W8g2ce5HN" : ("eyoZLXH0TFPIQYkh080yVH" ?
                  (7'h43) : ((8'h9e) ?
                      $unsigned($signed(wire57)) : (~&"yKKpfHGrSPh"))));
          reg4381 <= {$unsigned((&"Zi8"))};
        end
      reg4382 <= (reg4333 <= $unsigned("TqvLUtOSSGrm12epvJGThnQ"));
    end
  assign wire4383 = (forvar4345 ? $unsigned(reg4326[(3'h5):(1'h0)]) : "F8f");
  always
    @(posedge clk) begin
      reg4384 <= $signed((7'h4e));
      for (forvar4385 = (1'h0); (forvar4385 < (2'h3)); forvar4385 = (forvar4385 + (1'h1)))
        begin
          reg4386 <= $unsigned((~|$signed((&$unsigned(reg65)))));
          reg4387 <= (~((reg4325 ?
              $unsigned(reg4348) : ({forvar60} ?
                  ((7'h45) ? (8'ha1) : (8'ha2)) : (forvar4304 ?
                      wire4357 : wire4366))) >>> $signed("kui3M3VuMVEUDG1M")));
          for (forvar4388 = (1'h0); (forvar4388 < (3'h4)); forvar4388 = (forvar4388 + (1'h1)))
            begin
              reg4389 <= {(&$unsigned({(reg4348 ? reg4336 : reg4320),
                      (8'had)})),
                  ($signed($unsigned($unsigned(reg4356))) ?
                      "TPWoMw98mLLNGNiISYs51LA" : $unsigned("Yf544JVcui4zBVdb2CvgYZlt4"))};
              for (forvar4390 = (1'h0); (forvar4390 < (1'h0)); forvar4390 = (forvar4390 + (1'h1)))
                begin
                  reg4391 = ((-$unsigned((forvar4375 ?
                          (forvar4318 ? reg4338 : forvar4306) : (8'ha8)))) ?
                      reg4342 : "Mi0o5PWA1bEcbHYZTZ4BbK");
                end
            end
          for (forvar4392 = (1'h0); (forvar4392 < (1'h0)); forvar4392 = (forvar4392 + (1'h1)))
            begin
              reg4393 <= (~|reg4311[(5'h10):(4'he)]);
              reg4394 <= (reg4314 ?
                  (({{reg4335}} <<< ($signed(reg4323) > (reg4329 ?
                          (7'h4a) : (7'h49)))) ?
                      $signed(($signed(wire4357) ~^ (reg4339 ~^ (8'h9d)))) : ({forvar60,
                          $unsigned(reg4389)} > ((reg59 < reg4321) ?
                          reg4320 : (reg4342 ?
                              (8'ha4) : reg4312)))) : (~|$unsigned(($unsigned(reg4328) ?
                      (reg4320 ?
                          forvar4385 : forvar4296) : ((8'ha2) <= forvar4392)))));
            end
          reg4395 <= forvar4388;
          reg4396 <= (forvar4297 - $signed($signed($unsigned((~^reg4329)))));
        end
      reg4397 <= ((reg4384[(4'hb):(4'h8)] ?
          {(+$unsigned((8'hb9))), $signed((~|(8'hb5)))} : (reg4311 ?
              $unsigned(forvar4350) : $unsigned((reg63 ?
                  reg4327 : forvar4385)))) < {forvar4343, "zDvYHCgZRswE"});
      reg4398 <= (8'ha2);
      reg4399 <= (~wire54[(4'ha):(4'h9)]);
      reg4400 <= (($signed("Kx5YN") & (8'hbe)) <<< (((|reg4394[(3'h7):(2'h3)]) >> {(~^wire4317),
              (reg4309 ? reg4299 : forvar4343)}) ?
          (~&$signed((~forvar4331))) : reg4382));
    end
  assign wire4401 = {wire56[(5'h15):(3'h7)],
                        (($signed("JZPOmNIxSnqGO2qZuzGT") > ({forvar4371} ?
                                $signed(forvar4392) : reg4381[(4'hd):(4'hd)])) ?
                            ({reg4348,
                                {forvar4350,
                                    reg4314}} | $signed($unsigned(reg4319))) : "SZXHUs")};
  assign wire4402 = reg63[(2'h2):(1'h1)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module70
#( parameter param4291 = ((&((((8'ha7) && (8'hbc)) < ((8'ha6) ? (7'h4c) : (8'hb8))) | {((8'ha7) ? (8'ha1) : (8'hab))})) ? {(8'ha1)} : ((7'h4c) ? ((8'hba) + {((8'hb3) < (8'hb8))}) : ((((7'h4d) ? (8'hb1) : (8'hb9)) + (~^(7'h4d))) * (8'ha7)))) )
(y, clk, wire71, wire72, wire73, wire74, wire75);
  output wire [(32'h55c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire71;
  input wire [(5'h18):(1'h0)] wire72;
  input wire [(5'h1a):(1'h0)] wire73;
  input wire [(5'h1a):(1'h0)] wire74;
  input wire [(5'h16):(1'h0)] wire75;
  reg signed [(3'h6):(1'h0)] reg4280 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg4290 = (1'h0);
  reg [(5'h18):(1'h0)] reg4289 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4288 = (1'h0);
  reg [(3'h5):(1'h0)] reg4287 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4286 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4285 = (1'h0);
  reg [(4'hd):(1'h0)] reg4284 = (1'h0);
  reg [(4'h8):(1'h0)] reg4283 = (1'h0);
  reg [(4'hb):(1'h0)] reg4282 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4281 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4280 = (1'h0);
  reg [(4'hd):(1'h0)] reg4279 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4278 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4277 = (1'h0);
  wire signed [(5'h16):(1'h0)] wire4275;
  wire signed [(5'h18):(1'h0)] wire4273;
  wire [(4'he):(1'h0)] wire4271;
  wire signed [(3'h7):(1'h0)] wire4270;
  reg [(5'h16):(1'h0)] reg4269 = (1'h0);
  reg [(5'h19):(1'h0)] reg4268 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4267 = (1'h0);
  reg [(3'h6):(1'h0)] reg4266 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4265 = (1'h0);
  reg [(3'h7):(1'h0)] reg4264 = (1'h0);
  reg [(5'h12):(1'h0)] forvar4263 = (1'h0);
  reg [(3'h6):(1'h0)] reg4262 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire4261;
  reg signed [(5'h17):(1'h0)] reg4260 = (1'h0);
  wire [(3'h4):(1'h0)] wire4258;
  reg signed [(5'h18):(1'h0)] reg4257 = (1'h0);
  reg [(2'h2):(1'h0)] reg4256 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4255 = (1'h0);
  reg [(5'h18):(1'h0)] forvar4254 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4253 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4252 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4251 = (1'h0);
  reg [(5'h11):(1'h0)] reg4250 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4249 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4248 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar4247 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg4246 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4245 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4244 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4243 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar4242 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4241 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4240 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4239 = (1'h0);
  reg [(4'hd):(1'h0)] reg4238 = (1'h0);
  wire [(5'h1a):(1'h0)] wire4229;
  reg signed [(5'h16):(1'h0)] reg4228 = (1'h0);
  reg [(4'ha):(1'h0)] reg4227 = (1'h0);
  reg [(5'h1a):(1'h0)] reg4226 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4225 = (1'h0);
  reg [(5'h16):(1'h0)] reg4224 = (1'h0);
  wire [(5'h10):(1'h0)] wire4223;
  wire signed [(4'he):(1'h0)] wire4222;
  wire signed [(3'h4):(1'h0)] wire4221;
  reg signed [(5'h17):(1'h0)] reg4220 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4219 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire4218;
  reg signed [(5'h13):(1'h0)] reg4217 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4216 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4215 = (1'h0);
  reg [(4'hf):(1'h0)] reg4214 = (1'h0);
  reg [(4'hd):(1'h0)] reg4213 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg4212 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4211 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg4210 = (1'h0);
  reg [(5'h1a):(1'h0)] reg4209 = (1'h0);
  reg [(4'h9):(1'h0)] reg4208 = (1'h0);
  wire [(2'h2):(1'h0)] wire4206;
  reg signed [(3'h7):(1'h0)] reg4205 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg4204 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4203 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg4202 = (1'h0);
  reg [(5'h14):(1'h0)] reg4201 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4200 = (1'h0);
  reg [(5'h19):(1'h0)] forvar4199 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4198 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg4197 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg4196 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg77 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg78 = (1'h0);
  wire [(3'h4):(1'h0)] wire4194;
  reg [(4'hf):(1'h0)] reg4231 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire4232;
  wire [(5'h13):(1'h0)] wire4233;
  wire [(5'h14):(1'h0)] wire4234;
  wire [(5'h14):(1'h0)] wire4236;
  assign y = {reg4280,
                 reg4290,
                 reg4289,
                 reg4288,
                 reg4287,
                 reg4286,
                 forvar4285,
                 reg4284,
                 reg4283,
                 reg4282,
                 reg4281,
                 forvar4280,
                 reg4279,
                 reg4278,
                 reg4277,
                 wire4275,
                 wire4273,
                 wire4271,
                 wire4270,
                 reg4269,
                 reg4268,
                 reg4267,
                 reg4266,
                 reg4265,
                 reg4264,
                 forvar4263,
                 reg4262,
                 wire4261,
                 reg4260,
                 wire4258,
                 reg4257,
                 reg4256,
                 reg4255,
                 forvar4254,
                 reg4253,
                 reg4252,
                 reg4251,
                 reg4250,
                 reg4249,
                 reg4248,
                 forvar4247,
                 reg4246,
                 reg4245,
                 reg4244,
                 reg4243,
                 forvar4242,
                 reg4241,
                 forvar4240,
                 forvar4239,
                 reg4238,
                 wire4229,
                 reg4228,
                 reg4227,
                 reg4226,
                 reg4225,
                 reg4224,
                 wire4223,
                 wire4222,
                 wire4221,
                 reg4220,
                 forvar4219,
                 wire4218,
                 reg4217,
                 reg4216,
                 reg4215,
                 reg4214,
                 reg4213,
                 reg4212,
                 reg4211,
                 reg4210,
                 reg4209,
                 reg4208,
                 wire4206,
                 reg4205,
                 reg4204,
                 reg4203,
                 reg4202,
                 reg4201,
                 reg4200,
                 forvar4199,
                 reg4198,
                 reg4197,
                 reg4196,
                 reg76,
                 reg77,
                 reg78,
                 wire4194,
                 reg4231,
                 wire4232,
                 wire4233,
                 wire4234,
                 wire4236,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg76 <= (wire75[(5'h13):(2'h3)] ?
          $unsigned({wire75[(3'h6):(2'h2)],
              $unsigned("3aXBgoYW0fhTF1giqFv5xA1")}) : $signed("lodt9NDYVl8WxGap7QY"));
      reg77 <= (($unsigned($unsigned(wire73)) ?
          {wire73[(2'h3):(2'h3)]} : (({wire71} + wire73) >> reg76[(2'h3):(2'h2)])) == "TJ9W4V6tU");
      reg78 <= {"o4Q8V", wire74[(3'h4):(1'h0)]};
    end
  module79 modinst4195 (.wire80(reg76), .clk(clk), .wire81(reg78), .wire82(wire73), .y(wire4194), .wire84(reg77), .wire83(wire74));
  always
    @(posedge clk) begin
      reg4196 = "oLA6ASeXHkWY92";
      reg4197 <= $signed(((wire4194 ?
          wire4194[(3'h4):(3'h4)] : wire73) + wire75));
      reg4198 <= $unsigned(reg77[(3'h4):(1'h1)]);
      for (forvar4199 = (1'h0); (forvar4199 < (3'h4)); forvar4199 = (forvar4199 + (1'h1)))
        begin
          reg4200 <= forvar4199;
          reg4201 <= wire75[(4'h9):(3'h4)];
          reg4202 <= reg77;
          reg4203 <= $unsigned({reg4198});
        end
      reg4204 <= $unsigned(reg77);
      reg4205 <= reg78;
    end
  module779 modinst4207 (.y(wire4206), .wire783(reg78), .wire781(reg4197), .wire780(wire74), .wire782(reg4198), .clk(clk));
  always
    @(posedge clk) begin
      reg4208 <= (wire73 != ("anhY49EwDc7hWL5qyGUAvnPi" != (8'hb5)));
      reg4209 <= (&reg4204[(5'h19):(5'h11)]);
      reg4210 <= $signed((8'hb8));
      reg4211 <= "";
      reg4212 <= {($signed((-"4cwM3utNQrwy9giHEHfgd3riM")) < ($signed((forvar4199 - reg77)) <= $signed(reg4209[(1'h1):(1'h1)])))};
      reg4213 <= $signed((~(($signed(reg4201) ? $signed(reg4208) : (&(8'hbd))) ?
          (-(~|reg4202)) : reg77)));
    end
  always
    @(posedge clk) begin
      reg4214 = reg4213;
      reg4215 = wire4194[(2'h3):(1'h0)];
      reg4216 <= $signed((8'h9f));
      reg4217 = $unsigned(("ci" ?
          ($unsigned({wire4206}) != ({reg4212, wire73} ?
              (~&reg4198) : $signed(reg4209))) : wire72));
    end
  assign wire4218 = reg4205;
  always
    @(posedge clk) begin
      for (forvar4219 = (1'h0); (forvar4219 < (2'h2)); forvar4219 = (forvar4219 + (1'h1)))
        begin
          reg4220 <= (($unsigned((reg4197 ?
                  reg4213[(1'h0):(1'h0)] : $signed(reg4209))) ?
              (&"Fr9vxTuyu3U8s8mJzB3B7YiZ") : (^($signed(reg4214) | (reg4198 ?
                  (8'hab) : reg76)))) <<< "GX");
        end
    end
  assign wire4221 = ($signed(($unsigned((^~(8'ha8))) | "LGsuDd")) ^~ reg4217);
  assign wire4222 = $signed($unsigned({wire4218[(1'h0):(1'h0)]}));
  assign wire4223 = $signed(wire72);
  always
    @(posedge clk) begin
      reg4224 <= $unsigned((-$signed($unsigned($signed(reg76)))));
      reg4225 <= "g";
      reg4226 <= $unsigned((reg4225[(4'hf):(4'he)] && $signed(reg4213[(2'h3):(1'h1)])));
      reg4227 <= wire4222[(2'h2):(1'h0)];
      reg4228 <= $signed("Z2piZ40");
    end
  module1872 modinst4230 (wire4229, clk, reg4213, reg76, reg4204, forvar4199, reg4224);
  always
    @(posedge clk) begin
      reg4231 = wire4229[(4'h9):(1'h1)];
    end
  assign wire4232 = $signed((reg4224[(4'hd):(4'hc)] >> reg76[(3'h7):(3'h5)]));
  assign wire4233 = reg77[(2'h3):(2'h3)];
  module1210 modinst4235 (wire4234, clk, reg4228, wire74, reg4227, reg4201);
  module3450 modinst4237 (.clk(clk), .wire3455(reg4215), .wire3454(wire74), .wire3452(wire4229), .wire3453(reg4231), .wire3451(reg4198), .y(wire4236));
  always
    @(posedge clk) begin
      reg4238 <= "MphtK2iF";
      for (forvar4239 = (1'h0); (forvar4239 < (1'h1)); forvar4239 = (forvar4239 + (1'h1)))
        begin
          for (forvar4240 = (1'h0); (forvar4240 < (1'h0)); forvar4240 = (forvar4240 + (1'h1)))
            begin
              reg4241 <= wire4223;
              for (forvar4242 = (1'h0); (forvar4242 < (2'h2)); forvar4242 = (forvar4242 + (1'h1)))
                begin
                  reg4243 <= $signed(wire73);
                  reg4244 = $unsigned($unsigned(reg4198));
                  reg4245 = ("cMo7u15" ?
                      reg76[(5'h14):(1'h0)] : "xAE1f1W2B2OxvrCvTKtfOs");
                end
              reg4246 <= "GVhRRYfB6aW";
            end
          for (forvar4247 = (1'h0); (forvar4247 < (3'h4)); forvar4247 = (forvar4247 + (1'h1)))
            begin
              reg4248 <= reg4245;
              reg4249 <= "pDZ8YT2QEwdlwWkc8rOpFy";
              reg4250 <= (reg76[(3'h5):(2'h2)] ?
                  reg4203 : {$signed(reg4224[(2'h2):(1'h0)])});
            end
          reg4251 <= ($signed("4qcp0Vn8T57kUd") ? $unsigned(reg4250) : reg4210);
          reg4252 <= "ZrtM";
          reg4253 <= $unsigned(wire4206);
          for (forvar4254 = (1'h0); (forvar4254 < (1'h0)); forvar4254 = (forvar4254 + (1'h1)))
            begin
              reg4255 <= ($signed("stBLGQi") >> "shwy9kM");
              reg4256 <= reg4201[(3'h4):(2'h3)];
              reg4257 <= $unsigned("UzBPzmG3IwYnIB6Ym2");
            end
        end
    end
  module2696 modinst4259 (wire4258, clk, reg4213, forvar4219, reg4196, reg4246);
  always
    @(posedge clk) begin
      reg4260 <= (("FKJgiJ0InROxra" <= ((~(reg4253 ? wire4232 : reg4225)) ?
              $signed((~^reg4213)) : $unsigned($signed((7'h4a))))) ?
          $unsigned((~|(reg4196[(5'h12):(3'h5)] ?
              (^~wire4233) : {reg4220}))) : "gE0O4");
    end
  assign wire4261 = $unsigned($unsigned((((~^reg4201) << {reg77}) >>> (~^$signed(reg4226)))));
  always
    @(posedge clk) begin
      reg4262 = ($signed("9oBnYfrhVkynn1x2VS") ^ $unsigned($unsigned("vOqDnsHiYAvZsl91")));
      for (forvar4263 = (1'h0); (forvar4263 < (3'h4)); forvar4263 = (forvar4263 + (1'h1)))
        begin
          reg4264 <= ({(|"Nks2BKNk"),
              ({$unsigned(reg4243), "AkVPbugHW"} ?
                  $unsigned(reg4205[(3'h7):(3'h4)]) : $signed($unsigned((8'ha7))))} ~^ ($unsigned(reg4253) - "egZkBNzaCchdA6QK7h"));
          reg4265 <= forvar4254[(5'h10):(4'h8)];
          reg4266 <= "3ZLyYaXnTR";
          reg4267 <= (wire4233 == (~&$unsigned(($unsigned(reg4244) ?
              $unsigned(reg4216) : (7'h4a)))));
          reg4268 <= wire4194;
          reg4269 = reg4231;
        end
    end
  assign wire4270 = {reg4267[(1'h0):(1'h0)]};
  module1250 modinst4272 (.wire1254(reg4215), .clk(clk), .wire1252(reg4231), .wire1251(reg4200), .y(wire4271), .wire1253(reg4210));
  module3068 modinst4274 (.wire3072(wire4223), .clk(clk), .y(wire4273), .wire3069(reg4257), .wire3070(reg4212), .wire3071(reg4269));
  module1914 modinst4276 (wire4275, clk, reg4220, reg4264, reg4226, reg4209);
  always
    @(posedge clk) begin
      reg4277 <= ($signed((^~wire4261[(4'hb):(2'h3)])) ?
          (reg4251 == ("ntdhghgwzhhgvhWKqbYuHqiz" ?
              ({reg4244, forvar4219} ?
                  $unsigned(wire4271) : reg4268[(4'hb):(4'hb)]) : (|$signed((8'ha9))))) : wire4218[(4'h8):(3'h6)]);
      reg4278 = forvar4219[(4'h9):(3'h7)];
      if ((8'h9c))
        begin
          reg4279 <= "0ERqIr";
          for (forvar4280 = (1'h0); (forvar4280 < (2'h2)); forvar4280 = (forvar4280 + (1'h1)))
            begin
              reg4281 <= (+"4DllzlSaNFks04ODQu");
              reg4282 <= ("mgIbzHRBfO" ^~ reg4197[(5'h12):(4'he)]);
              reg4283 <= reg4212[(4'hd):(2'h2)];
              reg4284 <= (~&(~^wire75[(5'h16):(5'h15)]));
              for (forvar4285 = (1'h0); (forvar4285 < (2'h2)); forvar4285 = (forvar4285 + (1'h1)))
                begin
                  reg4286 <= {$unsigned($unsigned({$unsigned(reg4284),
                          $signed(reg4253)})),
                      $unsigned($signed($signed((^(8'h9d)))))};
                  reg4287 <= (({$signed(reg4284[(4'h9):(2'h2)])} > ($signed(reg4286) ~^ reg4282[(3'h6):(3'h4)])) ?
                      ((reg4266[(3'h6):(1'h0)] ?
                              "6" : (+wire74[(5'h15):(5'h12)])) ?
                          "7ViTkaL" : $unsigned(wire4270)) : ($signed($unsigned("mQGGCkU7mWyE6xKeyYAphrB")) ?
                          wire4273[(4'h8):(2'h2)] : $signed($unsigned((forvar4219 != (8'ha7))))));
                  reg4288 <= $signed(wire4233);
                end
            end
          reg4289 = $signed(reg4217);
          reg4290 = (~&"JWqmkiohat1XQJPLRka85gTo");
        end
      else
        begin
          reg4279 <= reg4197[(3'h6):(2'h3)];
          reg4280 <= wire4236;
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module79  (y, clk, wire84, wire83, wire82, wire81, wire80);
  output wire [(32'hef):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h1a):(1'h0)] wire84;
  input wire [(5'h1a):(1'h0)] wire83;
  input wire [(5'h1a):(1'h0)] wire82;
  input wire signed [(5'h12):(1'h0)] wire81;
  input wire [(5'h18):(1'h0)] wire80;
  wire signed [(4'h9):(1'h0)] wire4193;
  wire [(5'h18):(1'h0)] wire2679;
  reg [(5'h18):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg85 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire2681;
  wire [(4'hd):(1'h0)] wire2682;
  wire [(3'h4):(1'h0)] wire2683;
  wire signed [(2'h2):(1'h0)] wire2684;
  wire [(5'h17):(1'h0)] wire2685;
  reg signed [(4'ha):(1'h0)] reg2686 = (1'h0);
  reg [(5'h13):(1'h0)] reg2687 = (1'h0);
  reg [(5'h13):(1'h0)] reg2688 = (1'h0);
  wire [(5'h19):(1'h0)] wire2689;
  wire [(5'h19):(1'h0)] wire4191;
  assign y = {wire4193,
                 wire2679,
                 reg86,
                 reg85,
                 wire2681,
                 wire2682,
                 wire2683,
                 wire2684,
                 wire2685,
                 reg2686,
                 reg2687,
                 reg2688,
                 wire2689,
                 wire4191,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg85 <= wire84;
      reg86 <= {(("QWdDQRkMWbM0zp5W7YG" ?
                  $unsigned(reg85[(4'hb):(4'ha)]) : wire84) ?
              "QTgfPkbp4SsROhL2TeNnBSl9" : $signed(($unsigned(wire84) ?
                  $signed(wire84) : $signed(wire82)))),
          $unsigned(wire81)};
    end
  module87 modinst2680 (wire2679, clk, wire81, reg85, wire82, wire80, reg86);
  assign wire2681 = ("3dGpRw" ? (~^"AbK9JxIqbYhs2AMGaarYy4XS") : (7'h40));
  assign wire2682 = (&wire80);
  assign wire2683 = ($unsigned(reg85) ?
                        ((($signed(wire82) ?
                            (+wire82) : $unsigned(wire84)) << reg86) < (&((wire84 ?
                                (8'ha4) : wire82) ?
                            (wire80 ? wire83 : wire81) : {reg85,
                                reg85}))) : wire83);
  assign wire2684 = (+$unsigned("vXiIuxAB"));
  assign wire2685 = "0yUufZsCDPeu";
  always
    @(posedge clk) begin
      reg2686 = (8'hb1);
      reg2687 <= ((((~|(wire2684 && wire81)) - ($unsigned(wire82) ?
                  wire2679 : {wire2684, wire80})) ?
              $signed(reg2686) : $unsigned(wire2685[(4'h9):(4'h9)])) ?
          $unsigned(wire2682) : $signed("z"));
      reg2688 <= reg2686;
    end
  assign wire2689 = ((!($signed(reg2686) ?
                        ({wire2685} ?
                            "MDlnASuvfSe" : $signed((8'hb8))) : (reg2688 >> (8'h9f)))) * (((((7'h4b) - reg85) ^~ "T") ?
                        $signed(wire2684[(1'h0):(1'h0)]) : $unsigned($unsigned((8'ha9)))) && "mMuLWpg8xET"));
  module2690 modinst4192 (.wire2693(wire2685), .wire2692(wire2689), .clk(clk), .wire2691(reg2687), .y(wire4191), .wire2695(wire83), .wire2694(reg85));
  assign wire4193 = wire81[(3'h7):(1'h1)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2690
#( parameter param4190 = {((-(((8'ha5) << (8'hbe)) ? ((7'h43) ? (8'h9e) : (8'haa)) : ((7'h4b) && (8'ha2)))) ? (!(((7'h4a) ? (8'ha2) : (8'ha8)) ? ((7'h46) ^~ (8'h9c)) : (~&(8'hbf)))) : (7'h49))} )
(y, clk, wire2695, wire2694, wire2693, wire2692, wire2691);
  output wire [(32'h575):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h1a):(1'h0)] wire2695;
  input wire signed [(5'h1a):(1'h0)] wire2694;
  input wire [(5'h17):(1'h0)] wire2693;
  input wire signed [(5'h15):(1'h0)] wire2692;
  input wire signed [(5'h13):(1'h0)] wire2691;
  wire [(4'hf):(1'h0)] wire4188;
  wire signed [(5'h17):(1'h0)] wire4116;
  wire [(4'h8):(1'h0)] wire3977;
  wire [(5'h18):(1'h0)] wire3636;
  wire signed [(4'hf):(1'h0)] wire3447;
  wire [(2'h2):(1'h0)] wire3399;
  wire [(4'h8):(1'h0)] wire3202;
  wire signed [(5'h19):(1'h0)] wire2982;
  wire signed [(5'h13):(1'h0)] wire2839;
  reg [(5'h1a):(1'h0)] reg2780 = (1'h0);
  reg [(4'he):(1'h0)] reg2779 = (1'h0);
  reg [(5'h18):(1'h0)] reg2778 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2777 = (1'h0);
  reg [(3'h6):(1'h0)] reg2776 = (1'h0);
  reg [(5'h18):(1'h0)] reg2775 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2774 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2773 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2772 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2771 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2770 = (1'h0);
  reg [(5'h16):(1'h0)] reg2769 = (1'h0);
  wire [(5'h15):(1'h0)] wire2767;
  reg signed [(5'h1a):(1'h0)] reg2984 = (1'h0);
  reg [(4'hb):(1'h0)] reg2985 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar2986 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2987 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2988 = (1'h0);
  reg [(5'h17):(1'h0)] reg2989 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2990 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2991 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2992 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2993 = (1'h0);
  reg [(5'h11):(1'h0)] reg2994 = (1'h0);
  reg [(4'hb):(1'h0)] reg2995 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2996 = (1'h0);
  reg [(5'h19):(1'h0)] reg2997 = (1'h0);
  reg [(2'h2):(1'h0)] reg2998 = (1'h0);
  reg [(5'h19):(1'h0)] reg2999 = (1'h0);
  reg [(5'h15):(1'h0)] forvar3000 = (1'h0);
  reg [(4'he):(1'h0)] reg3001 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar3002 = (1'h0);
  reg [(5'h17):(1'h0)] reg3003 = (1'h0);
  reg [(5'h12):(1'h0)] reg3004 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar3005 = (1'h0);
  reg [(5'h11):(1'h0)] reg3006 = (1'h0);
  reg [(5'h12):(1'h0)] reg3007 = (1'h0);
  reg [(5'h13):(1'h0)] reg3008 = (1'h0);
  reg [(5'h13):(1'h0)] reg3009 = (1'h0);
  reg [(5'h17):(1'h0)] reg3010 = (1'h0);
  reg [(5'h12):(1'h0)] reg3011 = (1'h0);
  reg [(5'h12):(1'h0)] reg3012 = (1'h0);
  reg [(5'h14):(1'h0)] reg3013 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar3014 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3015 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3016 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3017 = (1'h0);
  wire [(4'ha):(1'h0)] wire3066;
  wire [(5'h14):(1'h0)] wire3449;
  wire signed [(5'h10):(1'h0)] wire3566;
  wire [(2'h3):(1'h0)] wire3694;
  reg signed [(5'h14):(1'h0)] reg3979 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3980 = (1'h0);
  wire [(5'h13):(1'h0)] wire4006;
  wire [(5'h14):(1'h0)] wire4008;
  reg signed [(5'h11):(1'h0)] reg4009 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4010 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg4011 = (1'h0);
  reg [(5'h19):(1'h0)] reg4012 = (1'h0);
  reg [(5'h11):(1'h0)] reg4013 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4014 = (1'h0);
  reg [(5'h11):(1'h0)] forvar4015 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4016 = (1'h0);
  reg [(5'h19):(1'h0)] reg4017 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4018 = (1'h0);
  reg [(2'h2):(1'h0)] reg4019 = (1'h0);
  reg [(5'h16):(1'h0)] reg4020 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4021 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg4022 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg4023 = (1'h0);
  wire [(5'h1a):(1'h0)] wire4114;
  assign y = {wire4188,
                 wire4116,
                 wire3977,
                 wire3636,
                 wire3447,
                 wire3399,
                 wire3202,
                 wire2982,
                 wire2839,
                 reg2780,
                 reg2779,
                 reg2778,
                 reg2777,
                 reg2776,
                 reg2775,
                 forvar2774,
                 forvar2773,
                 reg2772,
                 reg2771,
                 forvar2770,
                 reg2769,
                 wire2767,
                 reg2984,
                 reg2985,
                 forvar2986,
                 forvar2987,
                 forvar2988,
                 reg2989,
                 reg2990,
                 reg2991,
                 reg2992,
                 forvar2993,
                 reg2994,
                 reg2995,
                 reg2996,
                 reg2997,
                 reg2998,
                 reg2999,
                 forvar3000,
                 reg3001,
                 forvar3002,
                 reg3003,
                 reg3004,
                 forvar3005,
                 reg3006,
                 reg3007,
                 reg3008,
                 reg3009,
                 reg3010,
                 reg3011,
                 reg3012,
                 reg3013,
                 forvar3014,
                 reg3015,
                 reg3016,
                 reg3017,
                 wire3066,
                 wire3449,
                 wire3566,
                 wire3694,
                 reg3979,
                 reg3980,
                 wire4006,
                 wire4008,
                 reg4009,
                 forvar4010,
                 reg4011,
                 reg4012,
                 reg4013,
                 forvar4014,
                 forvar4015,
                 reg4016,
                 reg4017,
                 reg4018,
                 reg4019,
                 reg4020,
                 reg4021,
                 reg4022,
                 reg4023,
                 wire4114,
                 (1'h0)};
  module2696 modinst2768 (wire2767, clk, wire2693, wire2694, wire2695, wire2692);
  always
    @(posedge clk) begin
      reg2769 <= $signed(($unsigned((8'haa)) ?
          $signed($signed($signed(wire2691))) : wire2767[(3'h4):(1'h1)]));
      for (forvar2770 = (1'h0); (forvar2770 < (3'h4)); forvar2770 = (forvar2770 + (1'h1)))
        begin
          reg2771 <= $signed(wire2767);
          reg2772 <= wire2694;
          for (forvar2773 = (1'h0); (forvar2773 < (1'h0)); forvar2773 = (forvar2773 + (1'h1)))
            begin
              for (forvar2774 = (1'h0); (forvar2774 < (2'h3)); forvar2774 = (forvar2774 + (1'h1)))
                begin
                  reg2775 <= wire2694[(5'h1a):(4'hc)];
                  reg2776 <= forvar2770;
                  reg2777 <= {reg2769, "DorB6eaHQvzF7tIZI"};
                end
              reg2778 = $unsigned(((8'ha8) ?
                  "tL6yYcglaPEcmfYElv48Fv" : {{(wire2694 ^ wire2767)}}));
              reg2779 <= $unsigned($unsigned(({reg2772[(4'hc):(3'h5)]} & ((wire2694 - (8'ha5)) ~^ $unsigned(reg2777)))));
            end
        end
      reg2780 <= (~|$signed((~^(^~reg2779[(1'h1):(1'h1)]))));
    end
  module2781 modinst2840 (.wire2783(reg2775), .clk(clk), .wire2782(forvar2773), .wire2785(reg2777), .y(wire2839), .wire2784(wire2695));
  module2841 modinst2983 (wire2982, clk, forvar2770, reg2779, wire2693, reg2780, wire2767);
  always
    @(posedge clk) begin
      reg2984 <= $unsigned((^~((8'h9d) ?
          $unsigned("LhWPzPYvg") : wire2692[(4'hd):(4'h8)])));
      reg2985 <= "ur";
      for (forvar2986 = (1'h0); (forvar2986 < (2'h2)); forvar2986 = (forvar2986 + (1'h1)))
        begin
          for (forvar2987 = (1'h0); (forvar2987 < (2'h3)); forvar2987 = (forvar2987 + (1'h1)))
            begin
              for (forvar2988 = (1'h0); (forvar2988 < (3'h5)); forvar2988 = (forvar2988 + (1'h1)))
                begin
                  reg2989 <= {"NePFKPqtff7vZn0dw"};
                  reg2990 <= {"WQHMM8Dh"};
                  reg2991 <= (wire2691 ^ reg2989[(1'h1):(1'h0)]);
                end
            end
        end
      reg2992 <= ("5Upv8Y" ~^ reg2780[(5'h16):(2'h3)]);
    end
  always
    @(posedge clk) begin
      for (forvar2993 = (1'h0); (forvar2993 < (3'h4)); forvar2993 = (forvar2993 + (1'h1)))
        begin
          reg2994 <= reg2779;
          reg2995 <= wire2691;
          reg2996 <= (+$unsigned((|$unsigned($unsigned(reg2769)))));
          reg2997 <= reg2775[(5'h12):(1'h1)];
        end
      reg2998 = $unsigned((!(((~^wire2767) ?
              $unsigned(reg2984) : $unsigned(forvar2993)) ?
          {(forvar2773 ? reg2991 : forvar2993)} : (~^(forvar2770 ?
              reg2778 : reg2777)))));
      reg2999 = "DxyOAld7Lbd4E";
      for (forvar3000 = (1'h0); (forvar3000 < (3'h5)); forvar3000 = (forvar3000 + (1'h1)))
        begin
          reg3001 <= {reg2994[(4'hb):(4'hb)]};
          for (forvar3002 = (1'h0); (forvar3002 < (3'h5)); forvar3002 = (forvar3002 + (1'h1)))
            begin
              reg3003 <= wire2693[(5'h10):(3'h4)];
              reg3004 = "4lDJA4QigafmbmH3Rf4fz8l";
              for (forvar3005 = (1'h0); (forvar3005 < (1'h1)); forvar3005 = (forvar3005 + (1'h1)))
                begin
                  reg3006 <= reg2771;
                  reg3007 <= ($signed((((reg2989 & reg2985) ?
                          ((8'h9f) ?
                              forvar2774 : reg2996) : forvar2993) ^~ {reg3003[(5'h12):(4'hf)]})) ?
                      forvar3002[(2'h3):(1'h0)] : "xWsINhb5yTh3v");
                  reg3008 = "y";
                end
              reg3009 = ((reg2991 - reg2994[(3'h4):(1'h1)]) ?
                  {{"xTAzvDR9AacY3v"}} : $unsigned(forvar2988));
            end
          reg3010 <= forvar2773[(5'h10):(3'h6)];
          reg3011 <= reg2780[(3'h4):(3'h4)];
          reg3012 <= {reg2984};
          reg3013 <= "u0L2b6VERTdaR1IMfEGtHD";
        end
      for (forvar3014 = (1'h0); (forvar3014 < (1'h1)); forvar3014 = (forvar3014 + (1'h1)))
        begin
          reg3015 <= $signed(forvar3000);
          reg3016 <= (~^$unsigned("UvTesTpS4IUgfoDdMDKV79C3"));
        end
      reg3017 <= (!("WAJBt3mfSInwAv3PqiaE9xB0" ?
          $signed((|(reg2777 ?
              (8'ha2) : (8'hbd)))) : ((&(~^forvar3005)) >= reg2996[(1'h1):(1'h1)])));
    end
  module3018 modinst3067 (.y(wire3066), .wire3020(forvar3002), .wire3021(reg2989), .clk(clk), .wire3019(wire2839), .wire3022(reg2992), .wire3023(reg3006));
  module3068 modinst3203 (.clk(clk), .wire3072(reg2776), .wire3070(reg2991), .y(wire3202), .wire3069(reg3016), .wire3071(reg2769));
  module3204 modinst3400 (wire3399, clk, forvar3002, reg2992, wire3202, wire2982);
  module3401 modinst3448 (wire3447, clk, reg3010, wire2767, reg3008, reg2984, reg2992);
  assign wire3449 = $unsigned(($signed(((-reg2772) << (^~reg3015))) << "tdHkQE3RDcVXe6yI7Jyan5CQf"));
  module3450 modinst3567 (wire3566, clk, forvar3000, reg3009, reg3006, reg2997, reg2992);
  module3568 modinst3637 (wire3636, clk, forvar2987, forvar2993, reg3013, reg2992, reg2778);
  module3638 modinst3695 (.wire3642(forvar3014), .wire3643(forvar3000), .clk(clk), .wire3641(wire2693), .wire3640(reg2777), .y(wire3694), .wire3639(reg2991));
  module3696 modinst3978 (wire3977, clk, forvar2993, wire2693, reg2777, forvar3005, reg2779);
  always
    @(posedge clk) begin
      reg3979 <= {"S0gHaPRaMEiHpcKP", (+(|("rVRsZ1UTzgfUzbht" != wire2694)))};
      reg3980 <= ($signed({reg2996}) | wire2692);
    end
  module3981 modinst4007 (.wire3982(reg2984), .y(wire4006), .wire3984(forvar2986), .clk(clk), .wire3985(wire3449), .wire3983(reg3004));
  assign wire4008 = $signed(wire2982);
  always
    @(posedge clk) begin
      reg4009 <= $unsigned(((^~$unsigned($unsigned(reg2999))) == reg3004));
      for (forvar4010 = (1'h0); (forvar4010 < (3'h5)); forvar4010 = (forvar4010 + (1'h1)))
        begin
          reg4011 <= {$signed($unsigned($unsigned(reg3007)))};
        end
      reg4012 <= ((wire3399[(1'h0):(1'h0)] ?
          "wB1u8UIMll5Fcpq" : (8'hb7)) << wire3449[(5'h11):(3'h5)]);
      reg4013 <= {(&$unsigned(((reg3980 || reg2985) ?
              $signed(forvar4010) : $unsigned(wire2695))))};
      for (forvar4014 = (1'h0); (forvar4014 < (2'h2)); forvar4014 = (forvar4014 + (1'h1)))
        begin
          for (forvar4015 = (1'h0); (forvar4015 < (3'h4)); forvar4015 = (forvar4015 + (1'h1)))
            begin
              reg4016 <= (^~forvar2986[(3'h7):(3'h4)]);
              reg4017 <= ({reg2998[(1'h1):(1'h0)],
                      {(8'ha3),
                          ($unsigned(reg2992) > wire3566[(4'he):(4'h8)])}} ?
                  reg3006 : $unsigned((wire2695[(3'h4):(3'h4)] ?
                      (forvar4015[(4'h9):(4'h9)] ?
                          $unsigned(forvar3005) : (reg2996 << reg2994)) : wire3066[(4'ha):(4'ha)])));
              reg4018 <= $signed(({forvar3002, reg2772} ?
                  ("odiZaiAahxLhmi9" ?
                      reg3017[(4'hf):(4'hd)] : reg2994) : (!"MK8m4uCdr88CBC8KD9M")));
              reg4019 <= wire2767;
              reg4020 <= (wire3399[(1'h1):(1'h0)] ?
                  ((($unsigned(reg4018) ?
                          $unsigned(wire2694) : (forvar2993 * reg4016)) >> ((reg2777 ?
                              forvar2987 : (8'hac)) ?
                          $signed(reg3009) : $signed(wire3566))) ?
                      $unsigned({forvar3014[(2'h3):(2'h3)],
                          forvar3000[(2'h2):(1'h0)]}) : (&wire3694)) : reg2996);
            end
          reg4021 = $signed(($unsigned(($unsigned((7'h49)) ?
              reg3012[(2'h2):(1'h0)] : "WSX5QKbxYeUBChI")) << reg3980));
          reg4022 <= {(($unsigned(forvar2770[(2'h2):(1'h1)]) ?
                      $unsigned((-reg3006)) : ((reg3010 + reg3010) ?
                          (~|reg2998) : (forvar2993 > wire3636))) ?
                  "mrsVnBsNb" : $signed(reg2992)),
              (^(!$signed((reg4009 >= (8'h9c)))))};
          reg4023 <= $unsigned(wire4006[(4'hb):(4'ha)]);
        end
    end
  module4024 modinst4115 (wire4114, clk, reg3001, reg3012, wire4008, reg2772, wire3977);
  assign wire4116 = ((~^$signed($unsigned((^(8'hb9))))) > $unsigned({(wire2694[(3'h5):(3'h5)] * (reg2999 ?
                            reg4020 : reg2990)),
                        reg4019[(1'h1):(1'h0)]}));
  module4117 modinst4189 (wire4188, clk, wire3066, wire3636, forvar3002, forvar2986);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module87
#( parameter param2677 = (|((8'hb5) | ((((7'h49) ? (8'hbd) : (7'h45)) != ((8'haf) < (7'h4d))) ? ((~^(7'h45)) ? ((7'h45) <<< (8'ha2)) : ((8'hbb) ? (7'h4c) : (8'hb5))) : (((8'ha3) ? (8'hb2) : (8'haa)) >= {(8'hbe)}))))
, parameter param2678 = (~&(~&param2677)) )
(y, clk, wire88, wire89, wire90, wire91, wire92);
  output wire [(32'h9a2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire88;
  input wire [(4'ha):(1'h0)] wire89;
  input wire signed [(5'h11):(1'h0)] wire90;
  input wire [(3'h7):(1'h0)] wire91;
  input wire [(5'h18):(1'h0)] wire92;
  wire [(5'h1a):(1'h0)] wire2532;
  wire [(5'h16):(1'h0)] wire2281;
  wire signed [(4'hb):(1'h0)] wire1912;
  reg [(5'h18):(1'h0)] reg1871 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1870 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1869 = (1'h0);
  reg [(4'h8):(1'h0)] reg1868 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1867 = (1'h0);
  reg [(5'h10):(1'h0)] reg1866 = (1'h0);
  reg [(4'h9):(1'h0)] reg1865 = (1'h0);
  reg [(2'h3):(1'h0)] reg1864 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1863 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1862 = (1'h0);
  reg [(4'he):(1'h0)] forvar1861 = (1'h0);
  reg [(3'h7):(1'h0)] reg1860 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1859 = (1'h0);
  reg [(5'h19):(1'h0)] reg1858 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1857 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1856 = (1'h0);
  reg [(5'h11):(1'h0)] reg1855 = (1'h0);
  reg [(5'h13):(1'h0)] reg1854 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1853 = (1'h0);
  reg [(5'h19):(1'h0)] reg1852 = (1'h0);
  reg [(3'h4):(1'h0)] reg1851 = (1'h0);
  reg [(4'he):(1'h0)] forvar1850 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1849 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1848 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1847 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1846 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1845 = (1'h0);
  reg [(5'h15):(1'h0)] reg1844 = (1'h0);
  reg [(5'h10):(1'h0)] reg1843 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1842 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1841 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1840 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1839 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1838 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1837 = (1'h0);
  wire [(5'h16):(1'h0)] wire750;
  wire [(4'hd):(1'h0)] wire175;
  reg [(5'h1a):(1'h0)] forvar177 = (1'h0);
  reg [(5'h10):(1'h0)] forvar178 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar180 = (1'h0);
  reg [(5'h15):(1'h0)] reg181 = (1'h0);
  reg [(3'h7):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg183 = (1'h0);
  reg [(5'h13):(1'h0)] forvar184 = (1'h0);
  reg [(5'h19):(1'h0)] reg185 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg187 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg188 = (1'h0);
  reg [(4'hb):(1'h0)] reg189 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar190 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg191 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg192 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg193 = (1'h0);
  reg [(5'h13):(1'h0)] reg194 = (1'h0);
  reg [(5'h18):(1'h0)] forvar195 = (1'h0);
  reg [(4'hb):(1'h0)] forvar196 = (1'h0);
  reg [(5'h18):(1'h0)] reg197 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg200 = (1'h0);
  reg [(5'h16):(1'h0)] reg201 = (1'h0);
  reg [(3'h6):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg203 = (1'h0);
  reg [(5'h15):(1'h0)] reg204 = (1'h0);
  reg [(5'h16):(1'h0)] reg205 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg206 = (1'h0);
  reg [(5'h13):(1'h0)] forvar207 = (1'h0);
  reg [(4'hf):(1'h0)] forvar208 = (1'h0);
  reg [(4'he):(1'h0)] reg209 = (1'h0);
  reg [(5'h17):(1'h0)] reg210 = (1'h0);
  reg [(5'h18):(1'h0)] reg211 = (1'h0);
  reg [(5'h14):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg213 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg214 = (1'h0);
  reg [(4'h8):(1'h0)] forvar215 = (1'h0);
  reg [(4'hb):(1'h0)] reg216 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg217 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire218;
  wire [(3'h6):(1'h0)] wire446;
  reg [(3'h7):(1'h0)] reg448 = (1'h0);
  reg signed [(4'he):(1'h0)] reg449 = (1'h0);
  reg [(3'h6):(1'h0)] forvar450 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg451 = (1'h0);
  reg [(5'h15):(1'h0)] reg452 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar453 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg454 = (1'h0);
  reg [(5'h17):(1'h0)] reg455 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg456 = (1'h0);
  reg [(4'h8):(1'h0)] reg457 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg458 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire558;
  wire signed [(3'h5):(1'h0)] wire752;
  reg [(4'h8):(1'h0)] forvar753 = (1'h0);
  reg [(4'hf):(1'h0)] reg754 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg755 = (1'h0);
  reg [(3'h7):(1'h0)] forvar756 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg757 = (1'h0);
  reg [(4'h9):(1'h0)] reg758 = (1'h0);
  reg [(3'h5):(1'h0)] forvar759 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg760 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg761 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg762 = (1'h0);
  reg [(5'h17):(1'h0)] reg763 = (1'h0);
  reg [(5'h1a):(1'h0)] reg764 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg765 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg766 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar767 = (1'h0);
  reg [(4'h8):(1'h0)] reg768 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg769 = (1'h0);
  reg [(4'he):(1'h0)] reg770 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg771 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg772 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg773 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg774 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg775 = (1'h0);
  reg [(5'h19):(1'h0)] reg776 = (1'h0);
  reg [(5'h11):(1'h0)] reg777 = (1'h0);
  wire [(5'h15):(1'h0)] wire778;
  wire [(5'h17):(1'h0)] wire982;
  wire [(5'h14):(1'h0)] wire1011;
  wire [(5'h17):(1'h0)] wire1208;
  wire [(5'h10):(1'h0)] wire1248;
  wire [(5'h18):(1'h0)] wire1481;
  wire signed [(4'h9):(1'h0)] wire1672;
  wire signed [(4'hd):(1'h0)] wire1835;
  wire signed [(4'he):(1'h0)] wire2068;
  reg signed [(5'h11):(1'h0)] reg2070 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2071 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2072 = (1'h0);
  reg [(5'h17):(1'h0)] reg2073 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2074 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2075 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2074 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2075 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2076 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2077 = (1'h0);
  reg [(5'h13):(1'h0)] reg2078 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2079 = (1'h0);
  reg [(3'h4):(1'h0)] reg2080 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2081 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2082 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2083 = (1'h0);
  reg [(5'h18):(1'h0)] reg2084 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2085 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2086 = (1'h0);
  reg [(5'h15):(1'h0)] reg2087 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2088 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2089 = (1'h0);
  wire [(4'h9):(1'h0)] wire2279;
  wire [(3'h6):(1'h0)] wire2675;
  assign y = {wire2532,
                 wire2281,
                 wire1912,
                 reg1871,
                 reg1870,
                 reg1869,
                 reg1868,
                 reg1867,
                 reg1866,
                 reg1865,
                 reg1864,
                 reg1863,
                 forvar1862,
                 forvar1861,
                 reg1860,
                 forvar1859,
                 reg1858,
                 reg1857,
                 reg1856,
                 reg1855,
                 reg1854,
                 reg1853,
                 reg1852,
                 reg1851,
                 forvar1850,
                 reg1849,
                 forvar1848,
                 reg1847,
                 reg1846,
                 reg1845,
                 reg1844,
                 reg1843,
                 reg1842,
                 reg1841,
                 forvar1840,
                 reg1839,
                 forvar1838,
                 forvar1837,
                 wire750,
                 wire175,
                 forvar177,
                 forvar178,
                 reg179,
                 forvar180,
                 reg181,
                 reg182,
                 reg183,
                 forvar184,
                 reg185,
                 reg186,
                 reg187,
                 reg188,
                 reg189,
                 forvar190,
                 reg191,
                 reg192,
                 reg193,
                 reg194,
                 forvar195,
                 forvar196,
                 reg197,
                 reg198,
                 reg199,
                 reg200,
                 reg201,
                 reg202,
                 reg203,
                 reg204,
                 reg205,
                 reg206,
                 forvar207,
                 forvar208,
                 reg209,
                 reg210,
                 reg211,
                 reg212,
                 reg213,
                 reg214,
                 forvar215,
                 reg216,
                 reg217,
                 wire218,
                 wire446,
                 reg448,
                 reg449,
                 forvar450,
                 reg451,
                 reg452,
                 forvar453,
                 reg454,
                 reg455,
                 reg456,
                 reg457,
                 reg458,
                 wire558,
                 wire752,
                 forvar753,
                 reg754,
                 reg755,
                 forvar756,
                 reg757,
                 reg758,
                 forvar759,
                 reg760,
                 reg761,
                 reg762,
                 reg763,
                 reg764,
                 reg765,
                 reg766,
                 forvar767,
                 reg768,
                 reg769,
                 reg770,
                 reg771,
                 reg772,
                 reg773,
                 reg774,
                 reg775,
                 reg776,
                 reg777,
                 wire778,
                 wire982,
                 wire1011,
                 wire1208,
                 wire1248,
                 wire1481,
                 wire1672,
                 wire1835,
                 wire2068,
                 reg2070,
                 reg2071,
                 reg2072,
                 reg2073,
                 reg2074,
                 reg2075,
                 forvar2074,
                 forvar2075,
                 reg2076,
                 reg2077,
                 reg2078,
                 reg2079,
                 reg2080,
                 reg2081,
                 reg2082,
                 forvar2083,
                 reg2084,
                 reg2085,
                 reg2086,
                 reg2087,
                 reg2088,
                 reg2089,
                 wire2279,
                 wire2675,
                 (1'h0)};
  module93 modinst176 (.y(wire175), .wire94(wire90), .wire95(wire88), .wire96(wire89), .wire97(wire92), .clk(clk));
  always
    @(posedge clk) begin
      for (forvar177 = (1'h0); (forvar177 < (3'h4)); forvar177 = (forvar177 + (1'h1)))
        begin
          for (forvar178 = (1'h0); (forvar178 < (1'h0)); forvar178 = (forvar178 + (1'h1)))
            begin
              reg179 <= wire92;
              for (forvar180 = (1'h0); (forvar180 < (1'h0)); forvar180 = (forvar180 + (1'h1)))
                begin
                  reg181 <= ($signed($signed({$signed(forvar180),
                      wire88[(4'he):(3'h4)]})) ^~ wire89);
                  reg182 <= wire90[(3'h5):(1'h0)];
                end
              reg183 <= (((((reg181 >>> wire92) ?
                              "qgEgqnfOUIMn" : {forvar180}) ?
                          wire91[(2'h2):(1'h0)] : (forvar180[(3'h5):(1'h1)] ?
                              (wire88 ? forvar178 : wire91) : (~&reg182))) ?
                      (($signed(forvar177) == (|(8'ha8))) || $unsigned("OysANuhZxrvgWP9iiAyrPna")) : $unsigned((&wire89[(4'h9):(1'h1)]))) ?
                  wire92 : ({wire92} ?
                      $unsigned($unsigned({(8'ha4)})) : $signed((~(wire90 ^ wire90)))));
              for (forvar184 = (1'h0); (forvar184 < (3'h4)); forvar184 = (forvar184 + (1'h1)))
                begin
                  reg185 <= ((~^forvar180[(1'h0):(1'h0)]) ? reg179 : reg182);
                  reg186 <= $signed((^(8'hab)));
                  reg187 = "DV9VAu3QpkrlReemxtUF";
                  reg188 <= ({"RFEzR46FL9ZZnuL8FTCAp"} && wire89[(3'h5):(2'h2)]);
                  reg189 <= (((({forvar184, forvar177} ?
                      "mZ" : $unsigned(forvar184)) >> (+wire91[(2'h3):(2'h2)])) ^~ wire91) | (($signed((^wire89)) >>> (wire89 * (wire90 ?
                          forvar184 : reg183))) ?
                      (-$signed((&wire89))) : "pPTzlbpIYRN"));
                end
            end
          for (forvar190 = (1'h0); (forvar190 < (2'h2)); forvar190 = (forvar190 + (1'h1)))
            begin
              if ((forvar184[(2'h2):(2'h2)] >= $unsigned(wire91)))
                begin
                  reg191 = $signed($signed($signed(((~|forvar180) & (^wire88)))));
                  reg192 <= "WfN7hrBslDSATarS6zV";
                  reg193 = wire90;
                  reg194 <= (reg185[(1'h1):(1'h1)] ?
                      "kVIOwVWyaYXBSpz9AnZe" : reg183);
                end
              else
                begin
                  reg191 <= reg194[(4'hd):(2'h3)];
                  reg192 <= $signed($signed($signed(wire89[(3'h7):(3'h4)])));
                  reg193 <= $signed(forvar178[(4'h9):(3'h4)]);
                  reg194 <= $signed({reg182[(3'h5):(2'h2)]});
                end
            end
          for (forvar195 = (1'h0); (forvar195 < (1'h1)); forvar195 = (forvar195 + (1'h1)))
            begin
              for (forvar196 = (1'h0); (forvar196 < (2'h3)); forvar196 = (forvar196 + (1'h1)))
                begin
                  reg197 <= (("HGa5ilJ4Y7o" ?
                          $unsigned("e5mP") : $signed((wire92 >> wire89))) ?
                      forvar190 : $unsigned({(wire92 & ((8'hb2) ?
                              wire89 : wire175)),
                          wire88}));
                  reg198 <= $signed(forvar195[(1'h0):(1'h0)]);
                  reg199 = ($unsigned((forvar190[(3'h6):(1'h1)] ?
                      ((~reg179) >> $signed(reg181)) : {$unsigned(forvar180),
                          (forvar184 >>> wire89)})) >> (~|forvar196));
                  reg200 = $signed(((((^~wire91) ? {forvar177} : "9") ?
                      ((-(7'h4e)) == reg193) : reg199[(2'h3):(2'h3)]) == ({reg182[(3'h4):(2'h3)],
                      (reg179 & (7'h49))} || ($signed(reg185) ?
                      "ckZB" : (forvar177 ? reg194 : reg194)))));
                  reg201 <= $signed((forvar184[(4'h8):(3'h5)] ?
                      (&(!reg200[(5'h11):(3'h7)])) : forvar196[(4'ha):(3'h7)]));
                end
              reg202 <= (forvar178[(4'hf):(4'hb)] < reg194);
              reg203 = ((^$unsigned(((reg188 <<< reg200) ^ $unsigned(reg183)))) ?
                  $signed(reg191) : (|"m"));
              reg204 <= reg200[(5'h13):(4'hf)];
              reg205 <= {reg191,
                  (~|($unsigned($unsigned(forvar178)) ?
                      (7'h49) : $unsigned((~^forvar195))))};
              reg206 = reg204[(4'ha):(4'h8)];
            end
          for (forvar207 = (1'h0); (forvar207 < (2'h2)); forvar207 = (forvar207 + (1'h1)))
            begin
              for (forvar208 = (1'h0); (forvar208 < (1'h0)); forvar208 = (forvar208 + (1'h1)))
                begin
                  reg209 <= "aGyBkL";
                  reg210 <= "G";
                end
              reg211 <= $unsigned(reg183[(5'h12):(5'h10)]);
              reg212 <= (+reg210);
              reg213 <= reg205[(5'h15):(3'h5)];
              reg214 <= (((!"zb7ibgxAsQ0BXc73X7thRVpA") ?
                  $unsigned(forvar190) : $unsigned($unsigned({(8'hb8),
                      reg185}))) != reg199);
            end
          for (forvar215 = (1'h0); (forvar215 < (3'h4)); forvar215 = (forvar215 + (1'h1)))
            begin
              reg216 = reg194;
            end
        end
      reg217 <= $unsigned($signed($unsigned(reg205)));
    end
  assign wire218 = (8'hbb);
  module219 modinst447 (.clk(clk), .y(wire446), .wire220(reg191), .wire221(reg197), .wire222(reg213), .wire223(reg182));
  always
    @(posedge clk) begin
      reg448 <= "Ir";
      reg449 <= $signed((|$unsigned(wire92[(5'h11):(4'ha)])));
      for (forvar450 = (1'h0); (forvar450 < (2'h2)); forvar450 = (forvar450 + (1'h1)))
        begin
          reg451 <= $signed(forvar208[(3'h6):(1'h0)]);
          reg452 <= ((|reg179[(1'h0):(1'h0)]) ?
              ($signed("Kdsf28xL4U3C") ^~ $signed((^~$unsigned(wire92)))) : reg201[(4'hb):(1'h1)]);
          for (forvar453 = (1'h0); (forvar453 < (1'h0)); forvar453 = (forvar453 + (1'h1)))
            begin
              reg454 <= (+$signed((~reg199)));
            end
          reg455 <= reg454;
        end
      reg456 = reg185;
      reg457 <= wire175;
      reg458 <= "O0aAXuN9I0XM";
    end
  module459 modinst559 (wire558, clk, reg452, wire92, reg181, reg213, forvar190);
  module560 modinst751 (.wire562(reg202), .wire565(reg188), .y(wire750), .wire561(wire92), .wire563(forvar177), .wire564(reg185), .clk(clk));
  assign wire752 = {$unsigned($unsigned(reg191))};
  always
    @(posedge clk) begin
      for (forvar753 = (1'h0); (forvar753 < (2'h3)); forvar753 = (forvar753 + (1'h1)))
        begin
          reg754 <= ($signed(reg187) >> ($signed((!reg458[(4'hc):(4'h9)])) ~^ ($unsigned((&reg188)) >> {(!reg197),
              $signed(reg200)})));
          reg755 <= "";
          for (forvar756 = (1'h0); (forvar756 < (2'h3)); forvar756 = (forvar756 + (1'h1)))
            begin
              reg757 <= "O7CsPPy1UaOfGk2bT5";
              reg758 <= forvar195[(4'h8):(3'h4)];
              for (forvar759 = (1'h0); (forvar759 < (2'h3)); forvar759 = (forvar759 + (1'h1)))
                begin
                  reg760 <= "k4AYTWqmyBi8Hy10UIQ";
                  reg761 <= $unsigned($unsigned($signed($signed(reg193[(1'h0):(1'h0)]))));
                  reg762 = $signed((^~"grdvNAtWYSi5NtbvY"));
                  reg763 <= $signed(((~|(^~"E2XLxSQ2PpgamP")) ^ "1HoRqxJcD"));
                  reg764 <= $unsigned($unsigned(reg456[(1'h0):(1'h0)]));
                end
              reg765 <= reg457;
              reg766 <= $signed(($unsigned(reg185[(4'h9):(1'h1)]) == reg181));
              for (forvar767 = (1'h0); (forvar767 < (2'h2)); forvar767 = (forvar767 + (1'h1)))
                begin
                  reg768 <= ((8'h9d) ?
                      $signed(reg198[(5'h16):(2'h3)]) : forvar453[(2'h3):(1'h1)]);
                  reg769 <= reg213[(2'h2):(1'h0)];
                  reg770 = "ECvJW3";
                  reg771 <= $unsigned($signed(((|wire750[(4'ha):(4'h8)]) ?
                      (reg769 ^~ (wire89 ? reg205 : reg755)) : "xz")));
                  reg772 <= ((-{($unsigned(reg186) ?
                          (|wire89) : {forvar215})}) != "OKU4xcaQ3YA");
                  reg773 <= $unsigned($signed(reg452[(4'ha):(3'h6)]));
                end
            end
          reg774 <= forvar756[(2'h2):(1'h0)];
        end
      reg775 <= {$unsigned($unsigned(""))};
      reg776 <= $signed(reg189[(3'h4):(1'h0)]);
      reg777 <= ("7Q47ddbGlYRb0lTUCe2gfxgp" ^~ ($signed((^$signed(forvar450))) ?
          ((7'h40) + ((forvar450 ? (8'hb7) : forvar215) & (forvar184 ?
              reg457 : wire446))) : reg769));
    end
  assign wire778 = "sExxb3g8xe7YIqx";
  module779 modinst983 (.clk(clk), .wire781(reg213), .y(wire982), .wire782(reg183), .wire783(reg451), .wire780(reg764));
  module984 modinst1012 (wire1011, clk, reg204, reg197, reg761, forvar195);
  module1013 modinst1209 (.clk(clk), .y(wire1208), .wire1017(forvar180), .wire1014(reg454), .wire1015(reg203), .wire1016(reg199));
  module1210 modinst1249 (wire1248, clk, reg197, reg199, reg193, reg765);
  module1250 modinst1482 (.wire1253(reg203), .wire1254(wire558), .wire1251(forvar195), .wire1252(reg191), .clk(clk), .y(wire1481));
  module1483 modinst1673 (wire1672, clk, reg192, wire778, reg773, wire90);
  module1674 modinst1836 (wire1835, clk, reg774, forvar207, wire750, wire446, reg191);
  always
    @(posedge clk) begin
      for (forvar1837 = (1'h0); (forvar1837 < (1'h1)); forvar1837 = (forvar1837 + (1'h1)))
        begin
          for (forvar1838 = (1'h0); (forvar1838 < (3'h5)); forvar1838 = (forvar1838 + (1'h1)))
            begin
              reg1839 <= reg771;
              for (forvar1840 = (1'h0); (forvar1840 < (3'h5)); forvar1840 = (forvar1840 + (1'h1)))
                begin
                  reg1841 <= reg763;
                  reg1842 = reg754;
                  reg1843 = $signed({(^(reg182 >= $signed(reg194)))});
                  reg1844 <= $unsigned(reg217[(5'h14):(5'h11)]);
                  reg1845 <= $unsigned($unsigned((~&((reg765 * (8'h9c)) ?
                      $signed(forvar1838) : {reg200}))));
                end
            end
        end
      reg1846 <= reg451;
      reg1847 = ({wire218[(3'h5):(1'h1)],
          ($unsigned((reg186 ? wire175 : reg449)) ?
              ((8'ha9) ?
                  reg199 : (~&(8'had))) : ("uDoKXimaeIoM8" | reg179[(1'h0):(1'h0)]))} * $unsigned((8'hab)));
      for (forvar1848 = (1'h0); (forvar1848 < (3'h4)); forvar1848 = (forvar1848 + (1'h1)))
        begin
          reg1849 <= "GI";
          for (forvar1850 = (1'h0); (forvar1850 < (1'h1)); forvar1850 = (forvar1850 + (1'h1)))
            begin
              reg1851 = $unsigned((reg769 + "6HTdri1sek4GCa"));
              reg1852 <= reg766;
              reg1853 <= ($signed({(forvar453[(3'h4):(3'h4)] <= {(8'hb4)}),
                  (^{wire1835})}) <<< reg193);
              reg1854 = (($unsigned(("kPg0EHFCA" <= $unsigned(reg209))) ?
                  "3P9hOY6" : reg204) < (!$unsigned("cfBEiwM6JDOguYvh")));
            end
          reg1855 <= "pRZHrC144I";
          reg1856 <= ((+$signed($signed((^(8'ha1))))) ?
              (($signed("JVzQhRs") ?
                      $signed($unsigned(reg210)) : $signed((-(8'ha2)))) ?
                  ({(~|reg1845), wire218} == ($unsigned(forvar177) ?
                      (wire218 ?
                          reg185 : wire1481) : "otJiKgd8ktTOpZ2KlH1M")) : ($unsigned((reg760 ?
                      forvar184 : forvar1838)) != ((wire982 ? reg209 : reg768) ?
                      (reg1847 ^ forvar450) : reg186[(3'h6):(3'h5)]))) : $unsigned($signed(reg766[(3'h6):(2'h2)])));
          reg1857 <= (~&($unsigned((!(reg761 ?
              reg772 : reg197))) | ((reg458[(4'hf):(4'hf)] <<< $signed(reg772)) ?
              ((wire750 >>> (8'ha7)) || $signed(forvar450)) : forvar1848)));
          reg1858 <= ($unsigned((($unsigned(reg768) != {(8'h9f)}) | ((reg451 ?
                  forvar184 : wire446) ?
              ((8'hba) ?
                  wire1248 : reg213) : (forvar190 >= forvar196)))) <<< "UZDP2oPdnz2gQuWBgq7Eb");
        end
      for (forvar1859 = (1'h0); (forvar1859 < (1'h1)); forvar1859 = (forvar1859 + (1'h1)))
        begin
          reg1860 = ("kSJh1JbBD13neWU" <<< (wire750 ?
              {reg213} : $signed(reg760)));
          for (forvar1861 = (1'h0); (forvar1861 < (1'h0)); forvar1861 = (forvar1861 + (1'h1)))
            begin
              for (forvar1862 = (1'h0); (forvar1862 < (3'h5)); forvar1862 = (forvar1862 + (1'h1)))
                begin
                  reg1863 <= reg760;
                  reg1864 <= wire778;
                  reg1865 <= (~|(~|$unsigned($unsigned($unsigned(reg213)))));
                  reg1866 <= forvar1840[(1'h0):(1'h0)];
                  reg1867 <= "It2YyhICFeStJ4wgbYwwUh";
                  reg1868 = {(!(^reg1856)),
                      (((~|{wire1208, reg187}) * wire92[(5'h11):(3'h6)]) ?
                          reg179[(1'h1):(1'h1)] : "ZzK7ssPe")};
                end
              reg1869 <= (8'hbb);
              reg1870 <= (+($unsigned(((^~(7'h42)) << $signed(forvar1862))) << (&reg185)));
            end
        end
      reg1871 <= ({(|(8'ha6))} ?
          (&(!$signed($signed(reg214)))) : (-(~^{reg1854[(1'h1):(1'h0)]})));
    end
  module1872 modinst1913 (.wire1877(reg456), .y(wire1912), .wire1873(reg201), .wire1874(forvar190), .clk(clk), .wire1875(forvar1837), .wire1876(wire1481));
  module1914 modinst2069 (.wire1917(forvar1838), .y(wire2068), .clk(clk), .wire1916(reg1849), .wire1915(reg179), .wire1918(reg455));
  always
    @(posedge clk) begin
      reg2070 <= $unsigned(reg1871[(1'h1):(1'h0)]);
      if (((reg1871[(2'h3):(2'h2)] ~^ reg769[(5'h16):(4'h9)]) ?
          (((~(-(8'hb7))) >= "cM") ?
              reg1851 : forvar450[(1'h1):(1'h0)]) : ((&((reg197 <<< reg1845) ?
              $unsigned(reg763) : wire1481[(4'h8):(1'h1)])) < $unsigned(($signed(reg774) >= (~&reg191))))))
        begin
          reg2071 = ((~^{"DEJX2WPb0Gw32P6",
              ($signed(reg1852) << (forvar208 ?
                  (8'hb4) : reg1839))}) != ({(7'h45)} ?
              $unsigned($unsigned(wire982)) : "td53xZ2Oe"));
          reg2072 <= $signed((+(|({wire1208} ? $signed(forvar1861) : reg179))));
          reg2073 <= reg199[(5'h11):(5'h10)];
          reg2074 <= (~|(!{(reg1858 < "1nLaBEubgo5vMUYnReW")}));
          reg2075 <= $signed(reg768[(4'h8):(2'h2)]);
        end
      else
        begin
          reg2071 <= $signed(reg217[(5'h11):(5'h11)]);
          reg2072 <= ((~&({(&reg761), reg457} ?
              "D2a06sP2kmbDrE4w7okdO6" : reg448[(2'h2):(1'h0)])) * "GwGrCDLToUL99ECQekoht6");
          reg2073 <= (&$unsigned($signed((forvar756[(2'h2):(1'h0)] <= "ZNMKJ1xtkPuKrKR9MhzYYCu"))));
          for (forvar2074 = (1'h0); (forvar2074 < (3'h4)); forvar2074 = (forvar2074 + (1'h1)))
            begin
              for (forvar2075 = (1'h0); (forvar2075 < (1'h0)); forvar2075 = (forvar2075 + (1'h1)))
                begin
                  reg2076 <= {$signed($signed($unsigned((-(8'hab)))))};
                  reg2077 <= ({reg181[(4'hf):(1'h0)]} >= $signed((($unsigned(reg1847) ?
                          $unsigned(reg216) : $unsigned(reg185)) ?
                      ({forvar196,
                          forvar180} ^~ $signed(reg2071)) : wire1835)));
                  reg2078 <= $unsigned(wire91);
                  reg2079 <= ($signed((^~reg198)) >>> $unsigned({("vazifaUk5tebG" | reg771[(5'h12):(4'hf)]),
                      $signed($unsigned(wire2068))}));
                end
              reg2080 <= "gwthg9e";
              reg2081 <= "7oz9wBQw9XnrUkASroXBz";
              reg2082 <= reg2074;
            end
          for (forvar2083 = (1'h0); (forvar2083 < (2'h2)); forvar2083 = (forvar2083 + (1'h1)))
            begin
              reg2084 <= (!("NGCJP6r6rzxf" + ($unsigned((reg183 ?
                  (8'ha4) : (8'ha9))) << reg212[(4'hf):(3'h6)])));
              reg2085 <= "6FbURCu2";
              reg2086 <= {$unsigned((~^$unsigned({(8'hb9), reg197})))};
            end
        end
      reg2087 <= ((-(8'hb6)) <<< reg2084);
    end
  always
    @(posedge clk) begin
      reg2088 <= (~^(+reg206[(3'h4):(2'h2)]));
      reg2089 <= (($signed(forvar2083) ?
              (-($unsigned(wire89) ~^ (reg769 < reg187))) : reg1854[(4'hc):(4'ha)]) ?
          wire982[(4'hf):(4'hf)] : (~$unsigned(wire558)));
    end
  module2090 modinst2280 (.wire2094(reg1858), .wire2091(reg211), .y(wire2279), .wire2092(reg2088), .wire2095(reg203), .clk(clk), .wire2093(reg179));
  assign wire2281 = (^~(|$signed(forvar195[(3'h5):(2'h3)])));
  module2282 modinst2533 (.wire2286(reg205), .wire2284(reg1857), .wire2287(wire1835), .y(wire2532), .wire2285(reg213), .wire2283(reg1855), .clk(clk));
  module2534 modinst2676 (.wire2535(reg210), .wire2536(reg1860), .clk(clk), .wire2538(forvar178), .wire2537(wire175), .y(wire2675), .wire2539(forvar177));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2534
#( parameter param2673 = ((((~&((7'h4d) ? (8'hb7) : (7'h45))) ? (+((7'h4d) ? (8'haa) : (8'hb9))) : (~(~^(7'h4c)))) ? (~|(((8'hab) ? (7'h4e) : (8'ha3)) < ((8'h9e) ? (8'hae) : (8'haa)))) : (~{((8'hb7) ? (7'h4a) : (7'h42))})) ? (((^~((7'h4e) ? (7'h4d) : (8'h9c))) == (((7'h47) | (8'ha8)) ^ (~^(7'h43)))) ? (~&(((8'hab) ^~ (7'h42)) > (+(8'h9d)))) : ((((8'ha3) >> (8'hb6)) ^~ ((7'h4e) >> (7'h40))) >>> (((8'hb7) ? (8'hab) : (8'hb2)) ? ((8'hb4) <<< (8'ha0)) : {(8'ha3)}))) : ((|(((7'h42) ? (8'hb6) : (7'h47)) ? {(8'ha7), (7'h43)} : ((8'hb1) ? (8'hb2) : (8'hbc)))) - ((((7'h49) ? (8'h9c) : (7'h47)) >= {(7'h4c)}) > (((8'haf) ? (7'h4c) : (8'ha2)) <= {(8'hb9), (8'hb8)}))))
, parameter param2674 = ((8'hb8) == (8'hb7)) )
(y, clk, wire2539, wire2538, wire2537, wire2536, wire2535);
  output wire [(32'h78e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h16):(1'h0)] wire2539;
  input wire [(4'h8):(1'h0)] wire2538;
  input wire signed [(4'hc):(1'h0)] wire2537;
  input wire signed [(3'h7):(1'h0)] wire2536;
  input wire [(5'h17):(1'h0)] wire2535;
  reg signed [(3'h6):(1'h0)] reg2672 = (1'h0);
  reg [(4'he):(1'h0)] reg2671 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2670 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2669 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar2668 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2667 = (1'h0);
  wire [(5'h11):(1'h0)] wire2666;
  wire [(5'h1a):(1'h0)] wire2665;
  reg signed [(3'h7):(1'h0)] reg2664 = (1'h0);
  reg [(5'h15):(1'h0)] reg2663 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2662 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2661 = (1'h0);
  reg [(4'h9):(1'h0)] reg2660 = (1'h0);
  reg [(5'h15):(1'h0)] reg2659 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2658 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2657 = (1'h0);
  reg [(3'h7):(1'h0)] reg2656 = (1'h0);
  reg [(4'he):(1'h0)] forvar2655 = (1'h0);
  reg [(2'h3):(1'h0)] reg2654 = (1'h0);
  wire signed [(5'h18):(1'h0)] wire2653;
  wire [(5'h16):(1'h0)] wire2652;
  reg [(5'h11):(1'h0)] reg2651 = (1'h0);
  wire signed [(5'h19):(1'h0)] wire2650;
  reg signed [(3'h4):(1'h0)] reg2649 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2648 = (1'h0);
  reg [(4'h9):(1'h0)] reg2647 = (1'h0);
  reg [(4'hc):(1'h0)] reg2646 = (1'h0);
  reg [(4'he):(1'h0)] reg2645 = (1'h0);
  reg [(5'h11):(1'h0)] reg2644 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2643 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2642 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar2641 = (1'h0);
  reg [(5'h15):(1'h0)] reg2640 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2639 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2638 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2637 = (1'h0);
  reg [(4'ha):(1'h0)] reg2636 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2635 = (1'h0);
  reg [(5'h14):(1'h0)] reg2634 = (1'h0);
  reg [(5'h14):(1'h0)] reg2633 = (1'h0);
  reg [(3'h7):(1'h0)] reg2632 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2631 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2630 = (1'h0);
  reg [(2'h2):(1'h0)] reg2629 = (1'h0);
  reg [(5'h10):(1'h0)] reg2628 = (1'h0);
  reg [(3'h4):(1'h0)] reg2627 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2626 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2625 = (1'h0);
  reg [(4'hc):(1'h0)] reg2624 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2623 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2622 = (1'h0);
  reg [(5'h12):(1'h0)] forvar2621 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2620 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2619 = (1'h0);
  reg [(5'h14):(1'h0)] reg2618 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2617 = (1'h0);
  reg [(4'he):(1'h0)] reg2616 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2615 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2614 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2613 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2612 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2611 = (1'h0);
  reg [(5'h19):(1'h0)] reg2610 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire2609;
  reg [(4'h8):(1'h0)] reg2608 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2607 = (1'h0);
  reg [(5'h16):(1'h0)] reg2606 = (1'h0);
  reg [(2'h2):(1'h0)] reg2605 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2604 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2603 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2602 = (1'h0);
  reg [(4'hb):(1'h0)] reg2601 = (1'h0);
  reg [(2'h3):(1'h0)] reg2600 = (1'h0);
  reg [(3'h6):(1'h0)] reg2597 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2595 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2599 = (1'h0);
  reg [(5'h11):(1'h0)] reg2598 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2597 = (1'h0);
  reg [(4'he):(1'h0)] reg2596 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2595 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2594 = (1'h0);
  reg [(5'h12):(1'h0)] reg2593 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2592 = (1'h0);
  reg [(4'ha):(1'h0)] reg2591 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2590 = (1'h0);
  reg [(4'ha):(1'h0)] reg2589 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2588 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2587 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2586 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2585 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2584 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2583 = (1'h0);
  reg [(5'h17):(1'h0)] reg2582 = (1'h0);
  reg [(3'h7):(1'h0)] reg2581 = (1'h0);
  reg [(5'h12):(1'h0)] reg2580 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2579 = (1'h0);
  reg [(5'h13):(1'h0)] reg2578 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2577 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2576 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2575 = (1'h0);
  reg [(4'ha):(1'h0)] reg2574 = (1'h0);
  reg [(3'h7):(1'h0)] reg2573 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire2572;
  reg [(5'h16):(1'h0)] reg2571 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2570 = (1'h0);
  reg [(4'h8):(1'h0)] reg2569 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2568 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2567 = (1'h0);
  reg [(5'h12):(1'h0)] reg2566 = (1'h0);
  reg [(5'h13):(1'h0)] reg2565 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2564 = (1'h0);
  reg [(5'h11):(1'h0)] reg2563 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2562 = (1'h0);
  reg [(3'h6):(1'h0)] reg2561 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2559 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2556 = (1'h0);
  reg [(3'h7):(1'h0)] reg2560 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2559 = (1'h0);
  reg [(4'h9):(1'h0)] reg2553 = (1'h0);
  reg [(5'h13):(1'h0)] reg2558 = (1'h0);
  reg [(5'h13):(1'h0)] reg2557 = (1'h0);
  reg [(2'h3):(1'h0)] reg2556 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2555 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2554 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2553 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2552 = (1'h0);
  reg [(5'h13):(1'h0)] reg2551 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2550 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2549 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2548 = (1'h0);
  reg [(3'h5):(1'h0)] reg2547 = (1'h0);
  reg [(5'h15):(1'h0)] reg2546 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2545 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2544 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2543 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2542 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2541 = (1'h0);
  reg [(4'ha):(1'h0)] reg2540 = (1'h0);
  assign y = {reg2672,
                 reg2671,
                 reg2670,
                 reg2669,
                 forvar2668,
                 reg2667,
                 wire2666,
                 wire2665,
                 reg2664,
                 reg2663,
                 reg2662,
                 reg2661,
                 reg2660,
                 reg2659,
                 reg2658,
                 forvar2657,
                 reg2656,
                 forvar2655,
                 reg2654,
                 wire2653,
                 wire2652,
                 reg2651,
                 wire2650,
                 reg2649,
                 reg2648,
                 reg2647,
                 reg2646,
                 reg2645,
                 reg2644,
                 reg2643,
                 reg2642,
                 forvar2641,
                 reg2640,
                 forvar2639,
                 reg2638,
                 reg2637,
                 reg2636,
                 forvar2635,
                 reg2634,
                 reg2633,
                 reg2632,
                 reg2631,
                 reg2630,
                 reg2629,
                 reg2628,
                 reg2627,
                 reg2626,
                 reg2625,
                 reg2624,
                 reg2623,
                 forvar2622,
                 forvar2621,
                 reg2620,
                 reg2619,
                 reg2618,
                 reg2617,
                 reg2616,
                 reg2615,
                 reg2614,
                 reg2613,
                 reg2612,
                 reg2611,
                 reg2610,
                 wire2609,
                 reg2608,
                 reg2607,
                 reg2606,
                 reg2605,
                 reg2604,
                 reg2603,
                 reg2602,
                 reg2601,
                 reg2600,
                 reg2597,
                 forvar2595,
                 reg2599,
                 reg2598,
                 forvar2597,
                 reg2596,
                 reg2595,
                 reg2594,
                 reg2593,
                 reg2592,
                 reg2591,
                 forvar2590,
                 reg2589,
                 forvar2588,
                 forvar2587,
                 reg2586,
                 reg2585,
                 reg2584,
                 reg2583,
                 reg2582,
                 reg2581,
                 reg2580,
                 reg2579,
                 reg2578,
                 forvar2577,
                 reg2576,
                 forvar2575,
                 reg2574,
                 reg2573,
                 wire2572,
                 reg2571,
                 reg2570,
                 reg2569,
                 reg2568,
                 reg2567,
                 reg2566,
                 reg2565,
                 reg2564,
                 reg2563,
                 forvar2562,
                 reg2561,
                 reg2559,
                 forvar2556,
                 reg2560,
                 forvar2559,
                 reg2553,
                 reg2558,
                 reg2557,
                 reg2556,
                 reg2555,
                 reg2554,
                 forvar2553,
                 reg2552,
                 reg2551,
                 reg2550,
                 reg2549,
                 reg2548,
                 reg2547,
                 reg2546,
                 reg2545,
                 reg2544,
                 reg2543,
                 reg2542,
                 reg2541,
                 reg2540,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg2540 <= (&"B3K82cOHm");
      reg2541 = "4hmZnF9zRZSD9Yi";
      reg2542 <= (^wire2535[(4'h8):(4'h8)]);
      reg2543 <= (~^$signed((~|($signed(reg2540) ?
          $unsigned(wire2538) : $signed((8'hb9))))));
      reg2544 <= ("AsGWYSVC1O" ?
          ($unsigned($unsigned($signed((8'hb5)))) < $signed("Szhz3uUg")) : wire2538);
      reg2545 <= $signed(reg2543);
    end
  always
    @(posedge clk) begin
      reg2546 <= reg2540;
      reg2547 <= reg2546;
    end
  always
    @(posedge clk) begin
      reg2548 <= (~^reg2547[(1'h1):(1'h0)]);
      reg2549 <= "xp29ZvQz";
      if (wire2536[(3'h7):(2'h3)])
        begin
          if ("mJVOiA")
            begin
              reg2550 = reg2543[(4'ha):(3'h7)];
              reg2551 <= (~^{reg2545[(2'h2):(1'h0)]});
              reg2552 <= $signed(({(reg2540 ?
                      "owO5V4" : $signed(wire2538))} & $unsigned($signed((reg2540 <= reg2540)))));
              for (forvar2553 = (1'h0); (forvar2553 < (1'h0)); forvar2553 = (forvar2553 + (1'h1)))
                begin
                  reg2554 <= ("4ddg2R2WSJhAItsKxCGdbB3Cd" ?
                      ((reg2544 ?
                          reg2544 : $signed((reg2540 >= reg2549))) <= wire2536[(2'h2):(1'h1)]) : forvar2553[(5'h15):(4'he)]);
                  reg2555 <= ($unsigned((&(|"hRfp8msMsOiKCUDhYq3MvZKe"))) ?
                      $signed($signed(({reg2545} ?
                          {reg2552, forvar2553} : (wire2538 ?
                              reg2547 : (8'hba))))) : (~&$unsigned(((^~reg2548) ?
                          $unsigned(reg2545) : $signed(reg2551)))));
                  reg2556 <= $unsigned($signed($unsigned((^forvar2553))));
                  reg2557 <= $unsigned("Pz18Ox7");
                  reg2558 <= $signed(("R5iCSZO19WR" ?
                      forvar2553[(4'h8):(3'h4)] : $unsigned(((7'h48) ?
                          ((8'ha8) ? reg2540 : reg2547) : (!reg2556)))));
                end
            end
          else
            begin
              reg2550 = (-$unsigned($unsigned($unsigned($unsigned(reg2542)))));
              reg2551 <= ("4A1HS0KXaL4zKG2xf5GJt" >> $signed(reg2555[(5'h10):(3'h5)]));
              reg2552 = {wire2535[(4'h9):(2'h3)], reg2546};
              reg2553 = ((~|(~$signed((reg2540 & wire2538)))) ?
                  (+($unsigned((-reg2552)) ?
                      $signed((reg2546 ^ wire2537)) : $signed(reg2541[(2'h2):(1'h1)]))) : ((reg2556 >> ("74gY3AMk81GpDiWT1YRH" ?
                          "qTC" : $signed(wire2536))) ?
                      $signed(reg2543[(4'he):(2'h3)]) : $unsigned($unsigned((-(7'h4a))))));
            end
          for (forvar2559 = (1'h0); (forvar2559 < (2'h3)); forvar2559 = (forvar2559 + (1'h1)))
            begin
              reg2560 = $unsigned($unsigned((^reg2541[(3'h5):(3'h4)])));
            end
        end
      else
        begin
          reg2550 <= (~|({forvar2559[(2'h2):(1'h1)], reg2546} ?
              $unsigned((~&"dFSefAlSn")) : $unsigned($signed("7NTT41niLpILKT1P4X"))));
          reg2551 <= $unsigned(($unsigned(reg2555) <<< (^~$signed(reg2543[(4'ha):(1'h0)]))));
          reg2552 = $signed("0I5Guhf1M");
          for (forvar2553 = (1'h0); (forvar2553 < (2'h2)); forvar2553 = (forvar2553 + (1'h1)))
            begin
              reg2554 <= reg2546;
              reg2555 <= ($signed(forvar2559) <= {$unsigned($unsigned((reg2544 ~^ wire2535))),
                  (reg2558 ?
                      reg2560[(3'h5):(2'h3)] : $unsigned((|forvar2559)))});
              for (forvar2556 = (1'h0); (forvar2556 < (1'h0)); forvar2556 = (forvar2556 + (1'h1)))
                begin
                  reg2557 <= ($signed(wire2539[(5'h13):(3'h4)]) & (~$signed("faiMZPmkXnYCRFUklH1KHYOn")));
                  reg2558 <= forvar2553[(4'hf):(4'h9)];
                  reg2559 <= $signed(reg2548);
                  reg2560 <= wire2539[(4'hf):(4'hb)];
                end
              reg2561 <= $signed((&(wire2536[(1'h0):(1'h0)] <<< ((forvar2553 ?
                      reg2551 : (8'hbd)) ?
                  reg2540[(4'h8):(3'h4)] : $unsigned((7'h4d))))));
              for (forvar2562 = (1'h0); (forvar2562 < (3'h5)); forvar2562 = (forvar2562 + (1'h1)))
                begin
                  reg2563 <= "G62L57KlTxc";
                  reg2564 <= ((reg2556 ?
                      reg2561[(3'h4):(1'h0)] : (((reg2556 | wire2535) <<< reg2543) && reg2563)) && ({reg2545[(1'h1):(1'h1)],
                          reg2542[(4'he):(1'h1)]} ?
                      (((reg2560 != reg2545) ?
                          (reg2542 * (7'h4e)) : reg2546) * ("qSilRe3O15N9pO" ?
                          (~^reg2549) : (~&reg2541))) : ($unsigned($signed(reg2556)) << ($signed(forvar2559) > $signed(reg2559)))));
                end
              reg2565 = reg2549;
            end
        end
      reg2566 <= $unsigned(((^~((wire2537 ? forvar2559 : reg2553) ?
          reg2561 : (reg2552 ^ wire2535))) | $signed({reg2554})));
      reg2567 <= reg2558[(3'h4):(1'h0)];
      reg2568 <= $signed((~^($unsigned("cyE3Gf2YTPobvTVvW5Obn") ?
          "HX8MagvnF" : forvar2562[(3'h5):(3'h4)])));
    end
  always
    @(posedge clk) begin
      reg2569 = "73bUvDWITS99zSlPx";
      reg2570 <= {reg2543[(4'h9):(4'h9)]};
      reg2571 <= reg2558;
    end
  assign wire2572 = reg2542[(4'hc):(3'h4)];
  always
    @(posedge clk) begin
      reg2573 = "WGu9Vdop";
      reg2574 <= ($unsigned($unsigned(((&reg2569) >>> "WHpV7wGQ3ryZY21qsaMi66"))) ?
          $unsigned((8'hab)) : "Cdq86u4eUwSUNT0lYdq");
    end
  always
    @(posedge clk) begin
      for (forvar2575 = (1'h0); (forvar2575 < (2'h2)); forvar2575 = (forvar2575 + (1'h1)))
        begin
          reg2576 <= "aKgv5x1DXKqRJax4GIp0d";
          for (forvar2577 = (1'h0); (forvar2577 < (3'h4)); forvar2577 = (forvar2577 + (1'h1)))
            begin
              reg2578 <= $signed(reg2571);
              reg2579 <= $unsigned((($unsigned($signed(reg2566)) > $unsigned($signed(reg2573))) ?
                  "kHbOs4xOix624ExNOdz" : (reg2573[(3'h7):(3'h6)] ?
                      "MSxvV4XfZCLFFiafJybC" : $signed($signed(reg2571)))));
              reg2580 <= "vTI3k";
              reg2581 <= $signed((((wire2538 != $signed((8'haf))) ?
                      $unsigned({reg2560}) : $unsigned(reg2551)) ?
                  (+"oEGno2C39lV") : (8'ha2)));
            end
          reg2582 <= $unsigned(forvar2559[(3'h4):(1'h0)]);
          reg2583 = "UUelCEv1n";
          reg2584 <= "p66TRll7cOC9QsIh0lR5Uq0Ym";
          reg2585 <= $signed($unsigned((reg2574 != "zUdRe")));
        end
      reg2586 = (({(reg2543 ? forvar2559 : forvar2562)} ?
              reg2552 : $signed(((reg2579 ?
                  (8'hb9) : reg2549) >> "Nem7LrkEEaf"))) ?
          (!reg2560[(1'h0):(1'h0)]) : (reg2555 >> (|$unsigned((reg2578 != reg2582)))));
      for (forvar2587 = (1'h0); (forvar2587 < (3'h4)); forvar2587 = (forvar2587 + (1'h1)))
        begin
          for (forvar2588 = (1'h0); (forvar2588 < (2'h3)); forvar2588 = (forvar2588 + (1'h1)))
            begin
              reg2589 <= ($unsigned(reg2582[(4'hd):(4'hb)]) ?
                  (7'h48) : (8'hb6));
            end
          for (forvar2590 = (1'h0); (forvar2590 < (2'h2)); forvar2590 = (forvar2590 + (1'h1)))
            begin
              reg2591 <= reg2568[(3'h5):(2'h2)];
              reg2592 <= (^~"w62UL0JLSh9nLHbICb5");
              reg2593 <= $signed($unsigned({({wire2538,
                      reg2555} ~^ forvar2562[(3'h5):(3'h5)])}));
            end
          reg2594 <= (forvar2588 ?
              $unsigned("F6") : (+$signed("Kl31xV40TyNA9KDqei")));
          if (reg2559)
            begin
              reg2595 = (7'h48);
              reg2596 <= reg2545[(3'h4):(1'h0)];
              for (forvar2597 = (1'h0); (forvar2597 < (1'h1)); forvar2597 = (forvar2597 + (1'h1)))
                begin
                  reg2598 <= ({(|$unsigned((reg2553 ?
                          (8'h9c) : reg2594)))} == (($unsigned(reg2591[(3'h5):(2'h2)]) ?
                          reg2548[(3'h4):(1'h0)] : "47eOr1DJUXTO7WNuM") ?
                      $signed(reg2557[(3'h5):(2'h3)]) : (-wire2537)));
                  reg2599 <= ($signed($signed((8'had))) ?
                      ({wire2572[(3'h5):(2'h3)]} + $signed(($signed(reg2557) ?
                          wire2538 : $signed(forvar2575)))) : (~^{$unsigned(reg2583)}));
                end
            end
          else
            begin
              for (forvar2595 = (1'h0); (forvar2595 < (2'h2)); forvar2595 = (forvar2595 + (1'h1)))
                begin
                  reg2596 <= $signed((((~|(&reg2552)) ?
                          reg2580 : reg2563[(4'hd):(3'h7)]) ?
                      $signed($unsigned((reg2593 ?
                          reg2593 : reg2579))) : $signed(reg2569[(3'h5):(2'h2)])));
                  reg2597 = $unsigned("ZtgSOwqVpnG6vLqIP5c");
                  reg2598 = ("qc1y" - reg2586[(1'h1):(1'h0)]);
                  reg2599 = "IRPgyE6TTtOsKAwlbuZe";
                  reg2600 <= ($unsigned(("kw" ?
                          "Qal3miS0bAnmxnrU" : (-{reg2550}))) ?
                      forvar2553 : forvar2595[(4'hc):(4'hb)]);
                  reg2601 <= "m0HWLTBYbiVNqJv";
                end
              reg2602 <= {reg2582[(5'h15):(5'h11)],
                  $unsigned($unsigned(({wire2572} ~^ (reg2542 ?
                      (8'hbf) : forvar2553))))};
              reg2603 = ({{reg2581[(2'h3):(1'h1)],
                      ($signed(reg2563) ?
                          $unsigned(reg2585) : ((8'ha6) >= (8'hb6)))},
                  $unsigned(reg2553)} << ((!$signed({reg2579,
                  reg2578})) == ((|"kGGq1QhRGMno6") ?
                  {wire2538[(3'h7):(3'h6)]} : "Yo2UdPk5c")));
              reg2604 <= ("dfv" ? (~"P") : reg2546);
              reg2605 = "uuAdzbAy";
            end
          reg2606 = $unsigned(forvar2553[(3'h7):(3'h6)]);
          reg2607 <= "N";
        end
      reg2608 <= (!($signed(reg2571) ?
          (^~$signed((reg2571 ?
              forvar2597 : reg2605))) : $unsigned(("VF4Zq7OJofNmXcc1E" ?
              "" : "4RTkaxhD3TO8YD2b11"))));
    end
  assign wire2609 = reg2583[(3'h4):(1'h0)];
  always
    @(posedge clk) begin
      reg2610 <= {$signed("exAO9FfHk2pCWPmH8iO"), reg2573};
      reg2611 <= (8'hba);
      reg2612 <= reg2596;
      reg2613 <= (^~(+(-$signed(reg2545[(2'h2):(2'h2)]))));
      reg2614 <= forvar2556[(3'h6):(3'h6)];
    end
  always
    @(posedge clk) begin
      reg2615 <= (^{(((7'h48) ?
              (forvar2577 ?
                  reg2606 : reg2578) : reg2555[(3'h7):(1'h1)]) >>> $unsigned(reg2561[(3'h6):(2'h3)]))});
      reg2616 <= reg2603[(4'hd):(4'ha)];
    end
  always
    @(posedge clk) begin
      reg2617 <= "vKFaMYJRSDmGGFCsofAB";
      reg2618 <= reg2549;
      reg2619 <= reg2556;
      reg2620 <= (~^forvar2559);
      for (forvar2621 = (1'h0); (forvar2621 < (3'h5)); forvar2621 = (forvar2621 + (1'h1)))
        begin
          for (forvar2622 = (1'h0); (forvar2622 < (1'h1)); forvar2622 = (forvar2622 + (1'h1)))
            begin
              reg2623 <= $unsigned("ZxkeKVAv7hiHoqf4u1gvs");
              reg2624 = reg2563[(4'h9):(3'h7)];
              reg2625 <= $unsigned(reg2612);
              reg2626 <= "t8xoCw";
              reg2627 <= "ZgYw0Io";
              reg2628 = $signed((((8'hb4) < $signed($unsigned((8'hb1)))) - (reg2571 * "F26MtObDKpcUuq0")));
            end
          reg2629 = (|(wire2539 == $signed($unsigned({wire2539, (8'hb8)}))));
          reg2630 <= $signed("tz");
        end
      reg2631 <= (~&forvar2590[(1'h1):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg2632 <= ($unsigned("n3KfksJkh1CWuSFHHbizSqF5t") ?
          ((^~$signed((reg2548 >= (7'h46)))) >>> "f1zw7Ia73fr9mJqWI") : ($signed(reg2554[(5'h10):(4'hd)]) ?
              ($unsigned((reg2556 & reg2543)) == reg2614) : reg2544));
      reg2633 <= {$signed(((-"2VFLxIzb68Ef2ycszw0Bpmg") >>> $unsigned((reg2602 ?
              reg2591 : reg2547)))),
          $unsigned(reg2556[(1'h0):(1'h0)])};
      reg2634 <= wire2538[(3'h5):(1'h1)];
      for (forvar2635 = (1'h0); (forvar2635 < (3'h4)); forvar2635 = (forvar2635 + (1'h1)))
        begin
          reg2636 <= forvar2597;
          reg2637 = $signed(($signed(reg2613) && reg2585));
        end
      reg2638 <= (8'ha0);
      for (forvar2639 = (1'h0); (forvar2639 < (2'h3)); forvar2639 = (forvar2639 + (1'h1)))
        begin
          reg2640 = ((({{reg2566}, $unsigned(reg2542)} ?
                  $signed((&(8'h9e))) : ($signed(reg2617) ?
                      "mb1XNQlb" : "ne0oQOkRo6ZbNOnSaBRpf")) || {("1boXXOoKbwt3" >> $unsigned((8'h9d)))}) ?
              $signed((reg2554 && (^((8'ha4) ?
                  forvar2621 : (8'had))))) : reg2581[(3'h4):(1'h0)]);
          for (forvar2641 = (1'h0); (forvar2641 < (2'h2)); forvar2641 = (forvar2641 + (1'h1)))
            begin
              reg2642 <= (|"CztF4K7OBGEpHbOiLiOz");
            end
          reg2643 <= $signed({(|(^(reg2551 ? reg2634 : reg2633)))});
          reg2644 = reg2546[(3'h5):(2'h2)];
          reg2645 <= (reg2599 ?
              reg2558[(4'ha):(4'ha)] : (forvar2556[(5'h11):(4'hc)] ?
                  reg2545 : $unsigned(((wire2536 ? (8'hb8) : reg2579) ?
                      (~|reg2617) : forvar2641[(4'ha):(2'h3)]))));
        end
    end
  always
    @(posedge clk) begin
      reg2646 = reg2564[(1'h0):(1'h0)];
      reg2647 = "KOl6RkGalrO";
      reg2648 <= {$signed(reg2619)};
      reg2649 <= reg2582;
    end
  assign wire2650 = reg2580;
  always
    @(posedge clk) begin
      reg2651 <= ((8'ha7) ?
          ({(reg2544[(3'h6):(3'h6)] ?
                      $signed(forvar2635) : reg2599[(1'h0):(1'h0)]),
                  wire2538} ?
              $signed($unsigned(reg2592)) : "W7") : reg2579);
    end
  assign wire2652 = (reg2571[(4'hd):(4'h9)] - $signed(reg2585));
  assign wire2653 = $signed($unsigned("Z8Kq8H5"));
  always
    @(posedge clk) begin
      reg2654 = ($unsigned($signed(("JP" ?
              "xqalZpL02E" : $unsigned((8'ha0))))) ?
          $signed(reg2628[(5'h10):(3'h4)]) : $signed((+(reg2580 ?
              $signed((8'ha2)) : reg2636))));
      for (forvar2655 = (1'h0); (forvar2655 < (3'h4)); forvar2655 = (forvar2655 + (1'h1)))
        begin
          reg2656 <= (reg2589 ? (7'h45) : $unsigned((|reg2549[(3'h4):(2'h3)])));
          for (forvar2657 = (1'h0); (forvar2657 < (2'h2)); forvar2657 = (forvar2657 + (1'h1)))
            begin
              reg2658 = (~"vrSF9JRu15MEOF70ET0");
              reg2659 = $signed($unsigned(reg2555[(4'he):(4'ha)]));
              reg2660 = forvar2559;
              reg2661 <= "zpntw6Q9LUspPf8VYh003KWL";
            end
          reg2662 <= {(^~wire2538)};
        end
    end
  always
    @(posedge clk) begin
      reg2663 <= ((+reg2625[(4'hc):(2'h3)]) >>> forvar2556);
      reg2664 <= reg2596;
    end
  assign wire2665 = $signed("c3UBNgYVpqUQuXvIRF");
  assign wire2666 = ((("gyts2bY35XhTr3qFgwCIoN" ^~ wire2572[(3'h7):(1'h1)]) | ({((8'hae) ?
                                reg2586 : wire2665),
                            $signed(forvar2577)} ?
                        reg2603[(1'h1):(1'h1)] : "E1SO")) ~^ reg2560);
  always
    @(posedge clk) begin
      reg2667 <= ($unsigned(wire2572[(3'h7):(3'h5)]) ^ $signed(reg2589));
      for (forvar2668 = (1'h0); (forvar2668 < (1'h0)); forvar2668 = (forvar2668 + (1'h1)))
        begin
          reg2669 = ($signed(reg2578) || {{("gi2msWElk7I4Pzk" <= (reg2606 ?
                      reg2548 : reg2597)),
                  $unsigned((reg2540 ? reg2651 : reg2605))},
              reg2625[(2'h3):(1'h1)]});
          reg2670 <= (^{(&$signed((reg2567 ? reg2544 : reg2566)))});
          reg2671 = $unsigned("bwNPM0leLCBGBF7K");
        end
      reg2672 <= {"hEq67C3wKFtMvwt3xDt"};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2282
#(parameter param2531 = (+(8'ha4)))
(y, clk, wire2287, wire2286, wire2285, wire2284, wire2283);
  output wire [(32'hdeb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire2287;
  input wire signed [(5'h14):(1'h0)] wire2286;
  input wire [(2'h3):(1'h0)] wire2285;
  input wire [(4'he):(1'h0)] wire2284;
  input wire signed [(5'h11):(1'h0)] wire2283;
  wire signed [(4'hf):(1'h0)] wire2530;
  reg signed [(5'h13):(1'h0)] reg2529 = (1'h0);
  reg [(3'h5):(1'h0)] reg2528 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2527 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2526 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2525 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2524 = (1'h0);
  reg [(5'h13):(1'h0)] reg2523 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2522 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2521 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2520 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2519 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2518 = (1'h0);
  reg [(5'h10):(1'h0)] reg2517 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2516 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2515 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2514 = (1'h0);
  reg [(4'h9):(1'h0)] reg2513 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2512 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2511 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2510 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2509 = (1'h0);
  reg [(3'h4):(1'h0)] reg2508 = (1'h0);
  reg [(4'hd):(1'h0)] reg2507 = (1'h0);
  reg [(4'he):(1'h0)] reg2506 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2505 = (1'h0);
  reg [(5'h16):(1'h0)] forvar2504 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2503 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2502 = (1'h0);
  reg [(4'h8):(1'h0)] reg2501 = (1'h0);
  reg [(5'h17):(1'h0)] reg2500 = (1'h0);
  reg [(5'h17):(1'h0)] reg2499 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2498 = (1'h0);
  reg [(4'hb):(1'h0)] reg2497 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2496 = (1'h0);
  reg [(5'h12):(1'h0)] forvar2495 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2494 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2493 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2492 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2481 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2480 = (1'h0);
  reg [(4'ha):(1'h0)] reg2491 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2490 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2489 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2488 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2487 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2486 = (1'h0);
  reg [(4'hd):(1'h0)] reg2485 = (1'h0);
  reg [(5'h19):(1'h0)] reg2484 = (1'h0);
  reg [(4'h8):(1'h0)] reg2483 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2482 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2481 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2480 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2479 = (1'h0);
  reg [(2'h3):(1'h0)] reg2478 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2477 = (1'h0);
  reg [(4'h9):(1'h0)] reg2476 = (1'h0);
  reg [(3'h5):(1'h0)] reg2475 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2474 = (1'h0);
  reg [(5'h10):(1'h0)] reg2473 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2472 = (1'h0);
  reg [(5'h10):(1'h0)] reg2471 = (1'h0);
  reg [(5'h16):(1'h0)] reg2470 = (1'h0);
  reg [(5'h15):(1'h0)] reg2469 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2468 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2467 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2466 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2465 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2464 = (1'h0);
  reg [(3'h7):(1'h0)] reg2463 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2462 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2461 = (1'h0);
  reg [(5'h16):(1'h0)] reg2460 = (1'h0);
  reg [(5'h17):(1'h0)] reg2459 = (1'h0);
  reg [(4'ha):(1'h0)] reg2458 = (1'h0);
  reg [(3'h6):(1'h0)] reg2457 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2456 = (1'h0);
  reg [(5'h16):(1'h0)] reg2455 = (1'h0);
  reg [(3'h4):(1'h0)] reg2454 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2453 = (1'h0);
  reg [(2'h3):(1'h0)] reg2452 = (1'h0);
  reg [(4'hc):(1'h0)] reg2451 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2450 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2449 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2448 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2447 = (1'h0);
  reg [(2'h2):(1'h0)] reg2446 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2445 = (1'h0);
  wire [(4'h8):(1'h0)] wire2444;
  wire [(4'he):(1'h0)] wire2443;
  reg [(4'h8):(1'h0)] reg2442 = (1'h0);
  reg [(5'h11):(1'h0)] reg2441 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2440 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2439 = (1'h0);
  reg [(5'h10):(1'h0)] reg2438 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2437 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2436 = (1'h0);
  reg [(2'h3):(1'h0)] reg2435 = (1'h0);
  reg [(5'h19):(1'h0)] reg2434 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2433 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2432 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2431 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2430 = (1'h0);
  reg [(3'h5):(1'h0)] reg2429 = (1'h0);
  reg [(3'h5):(1'h0)] reg2428 = (1'h0);
  reg [(2'h2):(1'h0)] reg2427 = (1'h0);
  reg [(4'hf):(1'h0)] reg2426 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2425 = (1'h0);
  reg [(3'h5):(1'h0)] reg2424 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2423 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2422 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2421 = (1'h0);
  reg [(2'h3):(1'h0)] reg2420 = (1'h0);
  reg [(3'h5):(1'h0)] reg2419 = (1'h0);
  reg [(5'h19):(1'h0)] forvar2418 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar2417 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2416 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2415 = (1'h0);
  reg [(4'hb):(1'h0)] reg2414 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2413 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2412 = (1'h0);
  reg [(5'h13):(1'h0)] reg2411 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2410 = (1'h0);
  reg [(5'h18):(1'h0)] reg2409 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2408 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2407 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2406 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2405 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2404 = (1'h0);
  reg [(5'h19):(1'h0)] forvar2403 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2402 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2401 = (1'h0);
  reg [(5'h15):(1'h0)] reg2400 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2399 = (1'h0);
  reg [(5'h16):(1'h0)] reg2398 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2397 = (1'h0);
  reg [(4'hb):(1'h0)] reg2396 = (1'h0);
  reg [(5'h11):(1'h0)] reg2395 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2394 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2393 = (1'h0);
  reg [(3'h6):(1'h0)] reg2392 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2391 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2390 = (1'h0);
  reg [(5'h19):(1'h0)] reg2389 = (1'h0);
  reg [(3'h6):(1'h0)] reg2388 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2387 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2386 = (1'h0);
  reg [(3'h4):(1'h0)] reg2385 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2384 = (1'h0);
  reg [(4'hb):(1'h0)] reg2383 = (1'h0);
  reg [(5'h12):(1'h0)] reg2382 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2381 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2380 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2379 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2378 = (1'h0);
  reg [(5'h13):(1'h0)] reg2377 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2376 = (1'h0);
  reg [(4'ha):(1'h0)] reg2375 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2374 = (1'h0);
  reg [(2'h3):(1'h0)] reg2373 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2358 = (1'h0);
  reg [(3'h6):(1'h0)] reg2357 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2372 = (1'h0);
  reg [(5'h10):(1'h0)] reg2371 = (1'h0);
  reg [(3'h7):(1'h0)] reg2370 = (1'h0);
  reg [(5'h10):(1'h0)] reg2369 = (1'h0);
  reg [(5'h13):(1'h0)] reg2368 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2367 = (1'h0);
  reg [(4'hb):(1'h0)] reg2366 = (1'h0);
  reg [(4'ha):(1'h0)] reg2365 = (1'h0);
  reg [(5'h17):(1'h0)] reg2364 = (1'h0);
  reg [(4'h8):(1'h0)] reg2363 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2362 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2361 = (1'h0);
  reg [(3'h6):(1'h0)] reg2360 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2359 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2358 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2357 = (1'h0);
  reg [(4'ha):(1'h0)] reg2356 = (1'h0);
  reg [(3'h6):(1'h0)] reg2355 = (1'h0);
  reg [(3'h6):(1'h0)] reg2354 = (1'h0);
  reg [(5'h19):(1'h0)] reg2353 = (1'h0);
  reg [(4'h8):(1'h0)] reg2352 = (1'h0);
  wire [(5'h12):(1'h0)] wire2351;
  reg signed [(4'ha):(1'h0)] reg2350 = (1'h0);
  reg [(4'h8):(1'h0)] reg2339 = (1'h0);
  reg [(2'h3):(1'h0)] reg2349 = (1'h0);
  reg [(5'h16):(1'h0)] reg2348 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2347 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2346 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2345 = (1'h0);
  reg [(5'h18):(1'h0)] reg2344 = (1'h0);
  reg [(4'hb):(1'h0)] reg2343 = (1'h0);
  reg [(4'ha):(1'h0)] reg2342 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2341 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2340 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2339 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2338 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2337 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2336 = (1'h0);
  reg [(5'h11):(1'h0)] reg2335 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2334 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2333 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2332 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2331 = (1'h0);
  reg [(5'h19):(1'h0)] reg2330 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2329 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar2328 = (1'h0);
  reg [(4'hf):(1'h0)] reg2327 = (1'h0);
  reg [(4'hb):(1'h0)] reg2326 = (1'h0);
  reg [(5'h13):(1'h0)] reg2325 = (1'h0);
  reg [(5'h17):(1'h0)] reg2324 = (1'h0);
  reg [(5'h14):(1'h0)] reg2323 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar2322 = (1'h0);
  reg [(3'h7):(1'h0)] reg2321 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2320 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2319 = (1'h0);
  reg [(4'h8):(1'h0)] reg2318 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2317 = (1'h0);
  reg [(5'h10):(1'h0)] reg2316 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire2315;
  wire [(4'hf):(1'h0)] wire2314;
  reg signed [(5'h12):(1'h0)] reg2313 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2312 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2311 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2310 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2309 = (1'h0);
  reg [(5'h18):(1'h0)] forvar2308 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2307 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2306 = (1'h0);
  reg [(4'he):(1'h0)] reg2305 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2304 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2303 = (1'h0);
  reg [(4'h8):(1'h0)] reg2302 = (1'h0);
  reg [(5'h16):(1'h0)] reg2301 = (1'h0);
  reg [(3'h4):(1'h0)] reg2300 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2299 = (1'h0);
  reg [(4'h8):(1'h0)] reg2298 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2297 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2296 = (1'h0);
  reg [(3'h4):(1'h0)] reg2295 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2294 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2293 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2292 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2291 = (1'h0);
  reg [(5'h10):(1'h0)] reg2290 = (1'h0);
  reg [(5'h14):(1'h0)] reg2289 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2288 = (1'h0);
  assign y = {wire2530,
                 reg2529,
                 reg2528,
                 forvar2527,
                 reg2526,
                 reg2525,
                 reg2524,
                 reg2523,
                 reg2522,
                 reg2521,
                 reg2520,
                 forvar2519,
                 reg2518,
                 reg2517,
                 reg2516,
                 reg2515,
                 reg2514,
                 reg2513,
                 forvar2512,
                 forvar2511,
                 reg2510,
                 reg2509,
                 reg2508,
                 reg2507,
                 reg2506,
                 reg2505,
                 forvar2504,
                 reg2503,
                 reg2502,
                 reg2501,
                 reg2500,
                 reg2499,
                 reg2498,
                 reg2497,
                 reg2496,
                 forvar2495,
                 reg2494,
                 forvar2493,
                 reg2492,
                 reg2481,
                 forvar2480,
                 reg2491,
                 reg2490,
                 reg2489,
                 reg2488,
                 forvar2487,
                 reg2486,
                 reg2485,
                 reg2484,
                 reg2483,
                 reg2482,
                 forvar2481,
                 reg2480,
                 reg2479,
                 reg2478,
                 reg2477,
                 reg2476,
                 reg2475,
                 reg2474,
                 reg2473,
                 reg2472,
                 reg2471,
                 reg2470,
                 reg2469,
                 reg2468,
                 reg2467,
                 forvar2466,
                 forvar2465,
                 reg2464,
                 reg2463,
                 forvar2462,
                 reg2461,
                 reg2460,
                 reg2459,
                 reg2458,
                 reg2457,
                 reg2456,
                 reg2455,
                 reg2454,
                 forvar2453,
                 reg2452,
                 reg2451,
                 reg2450,
                 forvar2449,
                 forvar2448,
                 forvar2447,
                 reg2446,
                 forvar2445,
                 wire2444,
                 wire2443,
                 reg2442,
                 reg2441,
                 reg2440,
                 reg2439,
                 reg2438,
                 reg2437,
                 reg2436,
                 reg2435,
                 reg2434,
                 reg2433,
                 reg2432,
                 forvar2431,
                 reg2430,
                 reg2429,
                 reg2428,
                 reg2427,
                 reg2426,
                 forvar2425,
                 reg2424,
                 reg2423,
                 reg2422,
                 reg2421,
                 reg2420,
                 reg2419,
                 forvar2418,
                 forvar2417,
                 reg2416,
                 reg2415,
                 reg2414,
                 forvar2413,
                 reg2412,
                 reg2411,
                 reg2410,
                 reg2409,
                 reg2408,
                 forvar2407,
                 forvar2406,
                 reg2405,
                 reg2404,
                 forvar2403,
                 reg2402,
                 reg2401,
                 reg2400,
                 reg2399,
                 reg2398,
                 reg2397,
                 reg2396,
                 reg2395,
                 reg2394,
                 forvar2393,
                 reg2392,
                 reg2391,
                 reg2390,
                 reg2389,
                 reg2388,
                 reg2387,
                 forvar2386,
                 reg2385,
                 reg2384,
                 reg2383,
                 reg2382,
                 reg2381,
                 forvar2380,
                 reg2379,
                 forvar2378,
                 reg2377,
                 reg2376,
                 reg2375,
                 reg2374,
                 reg2373,
                 reg2358,
                 reg2357,
                 reg2372,
                 reg2371,
                 reg2370,
                 reg2369,
                 reg2368,
                 reg2367,
                 reg2366,
                 reg2365,
                 reg2364,
                 reg2363,
                 reg2362,
                 reg2361,
                 reg2360,
                 reg2359,
                 forvar2358,
                 forvar2357,
                 reg2356,
                 reg2355,
                 reg2354,
                 reg2353,
                 reg2352,
                 wire2351,
                 reg2350,
                 reg2339,
                 reg2349,
                 reg2348,
                 reg2347,
                 reg2346,
                 reg2345,
                 reg2344,
                 reg2343,
                 reg2342,
                 reg2341,
                 reg2340,
                 forvar2339,
                 reg2338,
                 reg2337,
                 reg2336,
                 reg2335,
                 reg2334,
                 reg2333,
                 forvar2332,
                 forvar2331,
                 reg2330,
                 reg2329,
                 forvar2328,
                 reg2327,
                 reg2326,
                 reg2325,
                 reg2324,
                 reg2323,
                 forvar2322,
                 reg2321,
                 forvar2320,
                 reg2319,
                 reg2318,
                 forvar2317,
                 reg2316,
                 wire2315,
                 wire2314,
                 reg2313,
                 reg2312,
                 forvar2311,
                 forvar2310,
                 reg2309,
                 forvar2308,
                 reg2307,
                 reg2306,
                 reg2305,
                 reg2304,
                 reg2303,
                 reg2302,
                 reg2301,
                 reg2300,
                 forvar2299,
                 reg2298,
                 reg2297,
                 forvar2296,
                 reg2295,
                 reg2294,
                 forvar2293,
                 reg2292,
                 reg2291,
                 reg2290,
                 reg2289,
                 forvar2288,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar2288 = (1'h0); (forvar2288 < (1'h0)); forvar2288 = (forvar2288 + (1'h1)))
        begin
          reg2289 <= wire2283;
          reg2290 = {((reg2289 ?
                      wire2287[(1'h1):(1'h0)] : "Vpeh0MP9mUDUnCxotvRFYAQ") ?
                  (!(~|(reg2289 & wire2285))) : "mHv77TyxR")};
          reg2291 <= $signed(((~&wire2284) >= ("gHTN" ?
              $signed((^~forvar2288)) : ((wire2287 >= wire2284) & "rc3911todarwI4QA3ih6"))));
        end
      reg2292 = {reg2289[(2'h3):(2'h3)],
          ("h0NWMH6HeqdKgCJ4vochh" ?
              wire2287 : $unsigned(($signed(reg2289) | "6D9q0MMGR2K7dgKN")))};
    end
  always
    @(posedge clk) begin
      for (forvar2293 = (1'h0); (forvar2293 < (1'h1)); forvar2293 = (forvar2293 + (1'h1)))
        begin
          reg2294 <= ((|$signed(reg2292)) ?
              ("h" >> "4wwiSfJL1lR1lt6gc38g9lR0A") : reg2290[(3'h5):(3'h4)]);
          reg2295 <= forvar2288;
          for (forvar2296 = (1'h0); (forvar2296 < (1'h0)); forvar2296 = (forvar2296 + (1'h1)))
            begin
              reg2297 <= $signed((wire2287 < ($signed(wire2284) ?
                  (~|(reg2291 * wire2283)) : "Z")));
            end
        end
      reg2298 <= $signed((~|((forvar2293[(1'h0):(1'h0)] ?
          forvar2293[(1'h0):(1'h0)] : wire2284) & {((8'hbf) ?
              forvar2288 : forvar2293)})));
      for (forvar2299 = (1'h0); (forvar2299 < (3'h5)); forvar2299 = (forvar2299 + (1'h1)))
        begin
          reg2300 <= ($unsigned(($signed((~|(8'hb4))) ^ $signed($unsigned(forvar2299)))) ?
              (((-wire2284[(4'hb):(3'h7)]) ?
                      ("u" << wire2285[(2'h2):(1'h1)]) : (~^$signed(forvar2288))) ?
                  wire2287 : $signed(wire2287[(1'h0):(1'h0)])) : wire2285[(2'h3):(2'h3)]);
        end
      reg2301 <= $signed(forvar2299);
      reg2302 <= ((|(^~$signed(reg2298[(2'h2):(2'h2)]))) && reg2298[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg2303 <= (|reg2298[(1'h1):(1'h0)]);
      reg2304 <= $signed("O0gIo");
      reg2305 <= $unsigned((&$unsigned($unsigned("t2dH"))));
      reg2306 = $unsigned(reg2289);
      reg2307 <= $signed(wire2285[(2'h2):(1'h0)]);
      for (forvar2308 = (1'h0); (forvar2308 < (2'h2)); forvar2308 = (forvar2308 + (1'h1)))
        begin
          reg2309 <= $signed(reg2290[(4'hd):(3'h5)]);
          for (forvar2310 = (1'h0); (forvar2310 < (1'h0)); forvar2310 = (forvar2310 + (1'h1)))
            begin
              for (forvar2311 = (1'h0); (forvar2311 < (1'h1)); forvar2311 = (forvar2311 + (1'h1)))
                begin
                  reg2312 <= {({forvar2310[(3'h5):(1'h1)],
                              $signed($signed(reg2303))} ?
                          (^forvar2288) : (((reg2292 <= wire2284) ?
                                  (forvar2299 ~^ wire2286) : (forvar2299 == reg2304)) ?
                              (reg2292[(5'h10):(2'h3)] ?
                                  (reg2292 > reg2304) : $unsigned((8'hba))) : ("" ?
                                  $signed(forvar2299) : $signed(reg2289))))};
                end
              reg2313 <= ((+forvar2311[(4'h8):(4'h8)]) ^ (^{(reg2312[(1'h0):(1'h0)] + $signed(wire2284))}));
            end
        end
    end
  assign wire2314 = $unsigned(reg2292);
  assign wire2315 = "55ABTXztgmMRqIr";
  always
    @(posedge clk) begin
      reg2316 = ($unsigned((^(^(reg2290 ? (8'hbc) : (8'ha5))))) ?
          (8'ha0) : $signed("xDxarIkmFhT5PTOhlRE0kH"));
    end
  always
    @(posedge clk) begin
      for (forvar2317 = (1'h0); (forvar2317 < (1'h0)); forvar2317 = (forvar2317 + (1'h1)))
        begin
          reg2318 <= reg2316;
          reg2319 <= forvar2317[(1'h1):(1'h1)];
          for (forvar2320 = (1'h0); (forvar2320 < (3'h4)); forvar2320 = (forvar2320 + (1'h1)))
            begin
              reg2321 <= ((-reg2294[(4'he):(4'he)]) * $signed(((reg2292 != (reg2309 ?
                  (8'ha2) : forvar2311)) ^~ $signed((forvar2320 <= (8'ha5))))));
            end
          for (forvar2322 = (1'h0); (forvar2322 < (1'h0)); forvar2322 = (forvar2322 + (1'h1)))
            begin
              reg2323 = ((!(reg2309 == {(forvar2299 ?
                          forvar2288 : forvar2310)})) ?
                  (~$signed((forvar2320[(3'h7):(3'h6)] ?
                      "ya" : (reg2297 ?
                          reg2298 : forvar2311)))) : ($unsigned($signed($unsigned(reg2290))) << forvar2299[(2'h3):(2'h3)]));
              reg2324 <= (8'hb2);
              reg2325 = $signed($signed((~^reg2309[(3'h5):(1'h0)])));
            end
          reg2326 <= $signed(("cJKVxXOR2IK8rJHlf" | reg2312));
        end
      reg2327 <= reg2324;
      for (forvar2328 = (1'h0); (forvar2328 < (3'h4)); forvar2328 = (forvar2328 + (1'h1)))
        begin
          reg2329 <= reg2325;
          reg2330 <= ({"uAdU3tU7GWnFePofb"} >>> reg2324[(5'h14):(5'h13)]);
        end
      for (forvar2331 = (1'h0); (forvar2331 < (2'h2)); forvar2331 = (forvar2331 + (1'h1)))
        begin
          if (forvar2331)
            begin
              for (forvar2332 = (1'h0); (forvar2332 < (3'h4)); forvar2332 = (forvar2332 + (1'h1)))
                begin
                  reg2333 <= ("M6" ?
                      $unsigned($signed((&reg2307))) : "RcO4SkQ9qRGpHXqEfKKzO0z");
                  reg2334 <= (reg2298[(4'h8):(3'h4)] && reg2300[(1'h1):(1'h0)]);
                  reg2335 <= (-"nEyszp8uAu");
                  reg2336 = ((7'h48) ?
                      (((reg2329[(5'h19):(5'h19)] & $unsigned(reg2302)) <<< (-{reg2290})) ^~ (8'hbe)) : $signed(reg2294));
                  reg2337 = ("RArLPyQqUlnxJoUvWAr" | "Md");
                  reg2338 <= (reg2319[(4'h9):(2'h2)] * "QJm1dshb3vdfOzA4qiHt");
                end
              for (forvar2339 = (1'h0); (forvar2339 < (3'h5)); forvar2339 = (forvar2339 + (1'h1)))
                begin
                  reg2340 <= (forvar2339 ?
                      {reg2323[(3'h4):(3'h4)]} : {(|reg2327[(3'h7):(1'h1)]),
                          $signed((reg2300 - forvar2288))});
                  reg2341 <= ("EVRQ9L" == {$signed(reg2298)});
                  reg2342 <= (8'ha2);
                  reg2343 = reg2302;
                  reg2344 = reg2289[(2'h3):(1'h0)];
                  reg2345 <= {$unsigned({"yT0o7RwAD"}),
                      (reg2300[(3'h4):(1'h0)] ~^ (($signed(reg2295) ?
                              reg2312 : $unsigned(reg2319)) ?
                          ((forvar2339 <= forvar2332) ?
                              $signed(reg2291) : "ngFJIRZr1wl8pcQRBt8") : ($unsigned(reg2342) ^ (reg2307 ?
                              reg2304 : forvar2331))))};
                end
              reg2346 <= (^~forvar2299[(2'h3):(2'h2)]);
              reg2347 <= {"Rc8GOXw1wIlTiAa"};
              reg2348 <= forvar2310;
              reg2349 <= {(({(!reg2292), (reg2337 - reg2289)} ?
                          (-(forvar2339 ?
                              forvar2296 : (8'had))) : ((^~(7'h41)) | (reg2343 >> wire2284))) ?
                      $signed($unsigned((!forvar2339))) : "cBJz1BGFX"),
                  $signed((("yzdJHODh" ?
                      $unsigned((8'hb4)) : {forvar2320,
                          reg2303}) <= (^(&reg2342))))};
            end
          else
            begin
              for (forvar2332 = (1'h0); (forvar2332 < (1'h0)); forvar2332 = (forvar2332 + (1'h1)))
                begin
                  reg2333 = reg2341[(1'h1):(1'h1)];
                  reg2334 <= reg2329;
                  reg2335 <= forvar2299[(3'h4):(1'h1)];
                  reg2336 <= (reg2307 <= $unsigned((8'haf)));
                end
              reg2337 <= {wire2315[(3'h4):(3'h4)], reg2316};
              reg2338 <= (forvar2310[(2'h3):(1'h0)] <= ({(reg2321 ?
                      (+reg2312) : (reg2334 + reg2321))} & $unsigned("h926h1cyw")));
              reg2339 <= ($signed({$signed((reg2291 + forvar2339))}) <= $unsigned($unsigned($signed(reg2334[(1'h0):(1'h0)]))));
            end
          reg2350 = (|$unsigned($signed($signed(reg2345))));
        end
    end
  assign wire2351 = (-"ye92");
  always
    @(posedge clk) begin
      reg2352 <= reg2337;
      reg2353 = "CdSLzLg6g6kSrcP7Rbc6";
      reg2354 <= $unsigned({{reg2305},
          ({(reg2289 ^~ reg2339)} || $signed(forvar2308[(4'ha):(3'h5)]))});
      reg2355 <= {({(|reg2349[(1'h0):(1'h0)]), $unsigned($signed((8'ha8)))} ?
              ("SROwrAXARD6IkMG8Q" > ((!forvar2331) ?
                  "" : "yqg9SvXDJGzpp3dTLIn1")) : ($unsigned(reg2321) ?
                  {((8'hbe) ? reg2353 : reg2323)} : $signed(wire2315)))};
      reg2356 <= (reg2292 ?
          ({$unsigned((~|reg2352)),
                  (((7'h41) ? forvar2322 : forvar2293) && (&reg2297))} ?
              $unsigned("G") : reg2303[(3'h4):(1'h0)]) : $unsigned(reg2297[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      if ((^~reg2309))
        begin
          for (forvar2357 = (1'h0); (forvar2357 < (1'h0)); forvar2357 = (forvar2357 + (1'h1)))
            begin
              for (forvar2358 = (1'h0); (forvar2358 < (1'h0)); forvar2358 = (forvar2358 + (1'h1)))
                begin
                  reg2359 <= $unsigned($signed($unsigned((~&(forvar2331 ?
                      wire2315 : reg2307)))));
                  reg2360 <= (reg2348[(5'h10):(4'hb)] ?
                      ($unsigned($unsigned(reg2341)) ?
                          (((-reg2291) ?
                              reg2354 : ((8'ha1) ?
                                  (8'h9f) : reg2346)) ~^ (~|reg2330[(1'h0):(1'h0)])) : (forvar2296[(5'h15):(4'hd)] ^ forvar2310)) : $unsigned(reg2335));
                end
              reg2361 <= reg2292[(4'h8):(4'h8)];
              reg2362 = ((("8eplaqMcnGQRL2" ?
                      $signed(reg2305[(4'h8):(1'h0)]) : $signed($unsigned(reg2305))) ?
                  "lNiph9J" : reg2318[(4'h8):(3'h6)]) && reg2335[(4'hf):(2'h3)]);
              if ({"8DryJPgOz7qQuxg", {($unsigned((~^reg2354)) ^ reg2303)}})
                begin
                  reg2363 = reg2306;
                  reg2364 <= ((~"7xQM39lgfkxDfGW9") <<< reg2337);
                  reg2365 = $unsigned(((8'h9c) ?
                      $signed(("WMvcoWsodOV9HsU1yB5Ct" - reg2294)) : $unsigned(((^wire2314) ?
                          reg2291 : $signed(reg2361)))));
                  reg2366 <= ($unsigned(reg2354) || reg2300[(1'h0):(1'h0)]);
                end
              else
                begin
                  reg2363 <= forvar2317;
                  reg2364 = wire2284[(4'ha):(4'h9)];
                  reg2365 <= $signed($signed($signed($unsigned(reg2333))));
                  reg2366 <= ("cSCkREob7F" >= (&(~^(~^wire2284))));
                  reg2367 = (|(reg2334[(1'h0):(1'h0)] ?
                      (reg2337[(3'h5):(1'h1)] ~^ "zHOIvIbEb7Pnf5D60A") : $unsigned(((reg2353 ?
                          reg2333 : wire2283) < (reg2305 ?
                          forvar2288 : reg2359)))));
                end
              if ($unsigned($signed((~reg2324))))
                begin
                  reg2368 <= ((^~(~^$signed($signed(reg2297)))) >= reg2309[(3'h5):(2'h3)]);
                  reg2369 = $unsigned(reg2346[(5'h13):(5'h12)]);
                  reg2370 <= (^"d6ryJxpYT63XaI9E7yQVlS1kJ");
                end
              else
                begin
                  reg2368 <= ($signed("w") ?
                      "7VfSm9SomwavBldWd7S" : forvar2328[(2'h3):(1'h1)]);
                  reg2369 = "tYa";
                end
              reg2371 <= "T8u69sI8zHuXDeLHLFVy";
            end
          reg2372 <= ((~|reg2295[(1'h1):(1'h1)]) - reg2326);
        end
      else
        begin
          reg2357 <= $signed(reg2344);
          reg2358 = reg2350[(3'h7):(1'h0)];
          reg2359 <= $signed($unsigned(reg2336[(1'h1):(1'h0)]));
        end
    end
  always
    @(posedge clk) begin
      reg2373 <= ((({"", reg2295} ?
                  ((-reg2350) ? reg2370 : (|forvar2339)) : (7'h40)) ?
              {reg2316,
                  "m1by0oCPDkwuzw0m"} : (reg2358 && $signed("Mw7JMSYUo"))) ?
          ("dWen00Zqfc3M0i7bsyh7FANY9" ?
              $unsigned(((reg2356 ? reg2302 : (7'h44)) ?
                  (forvar2311 & reg2370) : (reg2312 ?
                      (7'h4c) : reg2302))) : {((reg2354 ? reg2368 : (8'hbe)) ?
                      (7'h47) : (reg2371 <= reg2353)),
                  (&(reg2353 ?
                      reg2321 : (7'h42)))}) : "9ipntc9Ds4IYWAX6JH7I7lT5x");
      reg2374 = forvar2310;
      reg2375 <= ((^~$unsigned(($unsigned((7'h46)) ?
          reg2329[(4'hb):(3'h5)] : (wire2287 ?
              wire2315 : (7'h44))))) || wire2287[(3'h7):(3'h4)]);
      reg2376 <= $signed(((({forvar2293} ?
              "kxRlnTrlGmbfxdwmbhgdzN" : (reg2359 ?
                  (8'ha1) : reg2300)) << (7'h4c)) ?
          (reg2329 <<< (~&"HK")) : "KlSu"));
      reg2377 <= "UaMz";
      for (forvar2378 = (1'h0); (forvar2378 < (3'h4)); forvar2378 = (forvar2378 + (1'h1)))
        begin
          reg2379 <= ($signed("k4rHG") - {$unsigned(reg2377),
              $signed($unsigned({reg2313}))});
          for (forvar2380 = (1'h0); (forvar2380 < (1'h1)); forvar2380 = (forvar2380 + (1'h1)))
            begin
              reg2381 <= ((+($unsigned($unsigned(reg2313)) | $signed((reg2343 ?
                  reg2319 : reg2312)))) ^~ reg2304[(4'he):(2'h2)]);
              reg2382 <= $unsigned($signed(reg2292));
              reg2383 <= (^(reg2304[(1'h0):(1'h0)] ?
                  (^"oB7cbL9F5p9t0VdtUis") : ($signed({wire2314,
                      reg2350}) ^~ reg2289)));
              reg2384 = (reg2348[(4'h9):(3'h6)] ?
                  (~($signed($signed(reg2329)) * ((reg2339 <= (8'hb9)) || (reg2354 ?
                      reg2358 : reg2349)))) : ($unsigned($unsigned(reg2370)) > reg2291));
              reg2385 <= {($unsigned($unsigned($unsigned((8'ha6)))) ?
                      $unsigned(forvar2320) : $unsigned(reg2349))};
            end
          for (forvar2386 = (1'h0); (forvar2386 < (2'h3)); forvar2386 = (forvar2386 + (1'h1)))
            begin
              reg2387 <= "";
              reg2388 <= (&forvar2331[(1'h0):(1'h0)]);
            end
          reg2389 <= $signed(($signed((^(^~reg2372))) ?
              "iyrxv" : {$unsigned($signed(reg2325)),
                  "nkT66K7xnPHNhxdasQUkt72"}));
          reg2390 <= ({(8'hbc)} ?
              ("2vd6DU1uw9eMFv3az5HVV" ^ "W1xV0gHPmc0JHM2") : "6");
          reg2391 <= forvar2299;
        end
    end
  always
    @(posedge clk) begin
      reg2392 <= "z0t95T";
      for (forvar2393 = (1'h0); (forvar2393 < (3'h4)); forvar2393 = (forvar2393 + (1'h1)))
        begin
          reg2394 <= (~"TZ3tdDz9n");
          reg2395 <= ((((reg2313 ? reg2313 : $unsigned(forvar2331)) ?
                      $unsigned(reg2300) : reg2290[(3'h4):(2'h2)]) ?
                  (~^(&$unsigned(reg2347))) : wire2351) ?
              wire2283 : (forvar2380 > reg2392[(2'h2):(2'h2)]));
          reg2396 = reg2298;
          reg2397 = reg2366;
          reg2398 <= $signed($signed($unsigned($signed({reg2366, reg2396}))));
          reg2399 <= reg2298[(2'h3):(2'h2)];
        end
    end
  always
    @(posedge clk) begin
      reg2400 <= $unsigned((reg2348[(4'h8):(1'h0)] <= $signed(((reg2323 > reg2376) ?
          reg2379[(1'h0):(1'h0)] : (reg2361 || reg2373)))));
    end
  always
    @(posedge clk) begin
      reg2401 <= {{reg2330[(4'he):(4'hd)],
              $unsigned($signed($signed(reg2399)))},
          ((reg2365 ^ (7'h4a)) < $signed("lB0DGGz"))};
      reg2402 <= "Anxox4HuYv15kQiIJZ";
      for (forvar2403 = (1'h0); (forvar2403 < (1'h0)); forvar2403 = (forvar2403 + (1'h1)))
        begin
          reg2404 = ($signed(((8'hb2) + reg2291)) >> {reg2340[(5'h17):(2'h3)]});
          reg2405 <= $signed("wFWERqDtD6PFhGhVlcgc26Z");
        end
      for (forvar2406 = (1'h0); (forvar2406 < (3'h4)); forvar2406 = (forvar2406 + (1'h1)))
        begin
          for (forvar2407 = (1'h0); (forvar2407 < (2'h3)); forvar2407 = (forvar2407 + (1'h1)))
            begin
              reg2408 <= $signed(((~&reg2358) ^ forvar2407[(1'h0):(1'h0)]));
              reg2409 = $unsigned($signed(("s" <<< (reg2321 << "vZ"))));
              reg2410 <= reg2369;
            end
          reg2411 = "P1fuw1yXdlrRT";
        end
      reg2412 <= ($unsigned($signed(reg2397[(3'h6):(3'h6)])) && {"uPkaJ3Gk2nIp22JINf3yCcK",
          $signed(((reg2363 ? (8'had) : forvar2299) | ((7'h4c) ?
              reg2305 : wire2314)))});
      for (forvar2413 = (1'h0); (forvar2413 < (2'h2)); forvar2413 = (forvar2413 + (1'h1)))
        begin
          reg2414 <= reg2324[(4'ha):(3'h7)];
          reg2415 <= "XNKMH";
          reg2416 <= (|"4lwR0Mc");
          for (forvar2417 = (1'h0); (forvar2417 < (2'h3)); forvar2417 = (forvar2417 + (1'h1)))
            begin
              for (forvar2418 = (1'h0); (forvar2418 < (3'h4)); forvar2418 = (forvar2418 + (1'h1)))
                begin
                  reg2419 <= reg2297[(1'h0):(1'h0)];
                  reg2420 <= (&"PKmA");
                  reg2421 = wire2283;
                  reg2422 <= "dhbNsNN2";
                  reg2423 = (reg2400[(4'h9):(1'h1)] ? reg2371 : (~^""));
                  reg2424 <= {(reg2304[(4'hc):(3'h4)] ?
                          (~&$unsigned(((8'hbe) - reg2375))) : $unsigned((reg2373[(1'h1):(1'h0)] ?
                              "XQurxmTVKvOYIPlho75h0UB" : "ROPFnzEOvp1"))),
                      {(~^"X"), wire2283}};
                end
            end
          for (forvar2425 = (1'h0); (forvar2425 < (2'h3)); forvar2425 = (forvar2425 + (1'h1)))
            begin
              reg2426 <= (((^reg2301[(4'ha):(1'h0)]) >> (8'ha3)) - reg2369);
              reg2427 <= ($unsigned(reg2390) ?
                  ($signed($signed($signed(reg2401))) >> reg2362) : {forvar2328[(5'h12):(2'h3)]});
              reg2428 <= $signed((~"BfCMs9zau1sXN0RR"));
              reg2429 <= $unsigned("UfZBciRLkQGEtKa0siKHfY");
              reg2430 <= {$signed(((-$unsigned(wire2284)) ?
                      ((reg2423 * reg2345) <<< reg2390[(4'he):(1'h0)]) : $unsigned((^~reg2428)))),
                  "PZIzwxwnyE8w0"};
              for (forvar2431 = (1'h0); (forvar2431 < (1'h1)); forvar2431 = (forvar2431 + (1'h1)))
                begin
                  reg2432 = reg2356[(1'h1):(1'h0)];
                  reg2433 = (|$signed($signed(((^~(7'h40)) ?
                      wire2314 : "kDALrvgH7QoZoSs7ur02IpQF"))));
                  reg2434 <= reg2353;
                  reg2435 <= forvar2357[(3'h5):(2'h2)];
                end
            end
        end
    end
  always
    @(posedge clk) begin
      reg2436 <= wire2287[(2'h2):(1'h0)];
      reg2437 <= $signed(((+((forvar2407 | reg2358) ?
          (reg2326 ?
              reg2383 : reg2384) : reg2400[(3'h7):(1'h0)])) - $unsigned((8'hb6))));
      reg2438 <= $signed($unsigned($signed(wire2283)));
      reg2439 <= ($unsigned("EFH") != ($unsigned(reg2303[(2'h3):(2'h3)]) <= $signed($unsigned(((8'hbc) * reg2370)))));
      reg2440 <= $signed("WJrKAiN5eb1Qltxc8ir7e4");
      reg2441 = $unsigned((~"MPXw"));
    end
  always
    @(posedge clk) begin
      reg2442 <= (7'h40);
    end
  assign wire2443 = $unsigned(((~|($unsigned(reg2420) | ((7'h48) && reg2339))) << (7'h46)));
  assign wire2444 = ($signed(reg2402[(4'hf):(4'ha)]) ?
                        "EvAy32X" : (reg2294 ?
                            reg2295[(3'h4):(2'h3)] : $signed(reg2374)));
  always
    @(posedge clk) begin
      for (forvar2445 = (1'h0); (forvar2445 < (2'h2)); forvar2445 = (forvar2445 + (1'h1)))
        begin
          reg2446 <= $unsigned(forvar2311[(4'h8):(4'h8)]);
        end
      for (forvar2447 = (1'h0); (forvar2447 < (2'h3)); forvar2447 = (forvar2447 + (1'h1)))
        begin
          for (forvar2448 = (1'h0); (forvar2448 < (3'h5)); forvar2448 = (forvar2448 + (1'h1)))
            begin
              for (forvar2449 = (1'h0); (forvar2449 < (1'h1)); forvar2449 = (forvar2449 + (1'h1)))
                begin
                  reg2450 <= reg2303;
                end
              reg2451 <= $signed($unsigned({reg2424}));
              reg2452 <= ({(~$unsigned(forvar2308[(2'h3):(1'h1)]))} << $unsigned($signed((|(8'ha6)))));
              for (forvar2453 = (1'h0); (forvar2453 < (3'h5)); forvar2453 = (forvar2453 + (1'h1)))
                begin
                  reg2454 = (~&(-"InVsKonEKyRMt4dSX"));
                  reg2455 <= $signed(({reg2365[(1'h1):(1'h1)],
                      {$signed(wire2283)}} - ("fTbGv2PZtNDUdC" >>> (-$signed(reg2375)))));
                  reg2456 <= reg2404[(1'h0):(1'h0)];
                  reg2457 = (~$unsigned((8'ha7)));
                  reg2458 <= ($signed("OPTi2tZHIDWTsC8byDwX2BA") + (~&(8'hb8)));
                  reg2459 = "cQfpzIhCIdtV5eLMhdDUTPP";
                end
              reg2460 <= (((7'h4d) && ((~&reg2306[(2'h2):(1'h0)]) == $unsigned($unsigned(reg2375)))) || {{forvar2449[(3'h5):(3'h4)]},
                  reg2414[(4'h8):(3'h4)]});
            end
          reg2461 = $signed(((("tXrf8To81FIemHquL8b7hKDw" ?
                  $signed((8'hb4)) : reg2303) ?
              $unsigned((8'hbd)) : (!((8'hb1) ?
                  (8'hbd) : reg2391))) != ((&(reg2290 ?
              reg2361 : (8'ha2))) ^~ $unsigned("WkwVOUu"))));
          for (forvar2462 = (1'h0); (forvar2462 < (1'h1)); forvar2462 = (forvar2462 + (1'h1)))
            begin
              reg2463 <= $unsigned("M6szeDqkXuURyu");
              reg2464 = $unsigned(reg2304[(3'h7):(1'h0)]);
            end
          for (forvar2465 = (1'h0); (forvar2465 < (1'h0)); forvar2465 = (forvar2465 + (1'h1)))
            begin
              for (forvar2466 = (1'h0); (forvar2466 < (2'h2)); forvar2466 = (forvar2466 + (1'h1)))
                begin
                  reg2467 <= "0vzlzDf9wv1O0vt8Jb53kz";
                  reg2468 = $signed("ZSg");
                  reg2469 = (forvar2406[(1'h0):(1'h0)] ?
                      {((forvar2328[(3'h6):(1'h0)] ?
                                  (8'hb3) : reg2359[(5'h11):(4'h9)]) ?
                              ((forvar2445 - forvar2466) ?
                                  (forvar2448 ?
                                      reg2394 : reg2316) : forvar2378[(1'h0):(1'h0)]) : reg2371),
                          (reg2446 >>> ($unsigned(reg2372) + reg2412[(5'h15):(2'h3)]))} : reg2401[(4'h8):(3'h7)]);
                  reg2470 <= ("96mffRZNwZiMQ8" | reg2415);
                  reg2471 <= $unsigned((reg2333 ?
                      (+$unsigned(reg2354)) : {reg2390}));
                  reg2472 = reg2303;
                end
              reg2473 <= $unsigned((reg2337[(1'h0):(1'h0)] ?
                  $signed((~reg2432[(4'hc):(4'h8)])) : ($unsigned((reg2394 ?
                          (8'hb1) : reg2370)) ?
                      ((reg2305 > reg2363) == "7pBHhfmOAq8hngQQ21xAR3q") : forvar2465)));
              reg2474 <= (!{"qJnh1c8qUY6SzVuVnFaQsSh3F", forvar2310});
            end
          reg2475 = (reg2470[(4'hb):(1'h0)] ?
              reg2342[(4'h8):(3'h7)] : (+(reg2362 ?
                  ((reg2436 ? reg2303 : (8'hb2)) ?
                      (+reg2437) : forvar2328) : ("kR" ?
                      forvar2299[(4'h8):(3'h7)] : (8'h9e)))));
          reg2476 <= {(!{"S0SgaldXB"}), (7'h40)};
        end
    end
  always
    @(posedge clk) begin
      reg2477 <= ("RegEk1z1ErHV" ?
          ($unsigned(reg2452) ^~ "2KmPcc6cU5iCI4vaFQaF1UyL") : forvar2296);
      reg2478 <= ((reg2474[(4'hc):(4'h8)] | "h4ICnrW2EJ8Kx9") - ($signed((&$signed(forvar2431))) << (($unsigned(forvar2378) ?
              $unsigned(wire2351) : reg2414[(2'h3):(2'h2)]) ?
          reg2339[(3'h6):(3'h6)] : reg2434)));
      reg2479 <= (&(({"QgR74mMzna3oap6BkqavwhY",
              (reg2337 ? (8'haa) : forvar2431)} ?
          $unsigned($signed((7'h4d))) : (reg2290 ?
              (reg2387 ?
                  forvar2453 : (8'ha2)) : (reg2399 | reg2442))) + (reg2463 < $unsigned(forvar2386))));
    end
  always
    @(posedge clk) begin
      if (reg2354[(1'h1):(1'h0)])
        begin
          if (($unsigned($unsigned($unsigned((reg2410 && reg2349)))) ?
              ($unsigned("5rMZKbt0") ?
                  {"CnDt0Psbr0vUdrikD",
                      ((reg2463 ? reg2295 : wire2351) ?
                          reg2391[(4'hf):(1'h0)] : (~|wire2285))} : reg2454[(1'h1):(1'h1)]) : ($unsigned($unsigned(forvar2378[(1'h1):(1'h1)])) < (reg2290 ?
                  $signed($unsigned(forvar2406)) : ("k3Y4YRcVKXKT9PzEBKoE" * $signed(reg2437))))))
            begin
              reg2480 = ($unsigned(reg2450[(3'h7):(1'h0)]) ?
                  reg2337 : (("" ?
                      (^"56J1LQMePWzTnOnRkd0gXnbH0") : ((reg2469 <= reg2463) ?
                          (reg2301 || reg2402) : {forvar2358})) || "f8JxQuBpe1XN"));
              for (forvar2481 = (1'h0); (forvar2481 < (3'h5)); forvar2481 = (forvar2481 + (1'h1)))
                begin
                  reg2482 <= "FYztkKQ2pRRJ";
                  reg2483 <= $unsigned(((forvar2425 ?
                      reg2480[(1'h1):(1'h1)] : reg2458) & forvar2445[(5'h10):(3'h5)]));
                  reg2484 = $signed({{reg2319, reg2349[(2'h2):(2'h2)]}});
                  reg2485 = "wsptPuVINDph4wPqUe1ohktf";
                end
              reg2486 <= $signed($signed((~^({reg2367,
                  reg2305} != ((7'h4a) ^ reg2345)))));
              for (forvar2487 = (1'h0); (forvar2487 < (2'h3)); forvar2487 = (forvar2487 + (1'h1)))
                begin
                  reg2488 <= "uQKN";
                  reg2489 <= $signed((reg2354[(2'h2):(1'h1)] ?
                      $signed($unsigned($signed(reg2387))) : forvar2445));
                end
              reg2490 <= $signed(reg2441[(4'hd):(4'h9)]);
              reg2491 <= reg2490[(2'h3):(1'h0)];
            end
          else
            begin
              for (forvar2480 = (1'h0); (forvar2480 < (1'h1)); forvar2480 = (forvar2480 + (1'h1)))
                begin
                  reg2481 <= $signed((~&(-("tFUBxSOXJIHrxSJVf5J57f" ?
                      $signed(forvar2465) : {wire2314, reg2458}))));
                end
              reg2482 <= "5VTKTLx8hwk";
            end
          reg2492 <= "4frz";
          for (forvar2493 = (1'h0); (forvar2493 < (2'h2)); forvar2493 = (forvar2493 + (1'h1)))
            begin
              reg2494 <= $unsigned((forvar2339[(4'hd):(4'h9)] ?
                  $unsigned($unsigned($unsigned(reg2440))) : $unsigned("1Doxn7KfXi7cP")));
              for (forvar2495 = (1'h0); (forvar2495 < (1'h1)); forvar2495 = (forvar2495 + (1'h1)))
                begin
                  reg2496 <= "0qVEKwO6nT0LO";
                end
              reg2497 <= reg2423;
              reg2498 <= $signed($unsigned(forvar2449));
            end
          reg2499 <= (&$unsigned(((-forvar2481) ?
              reg2379 : forvar2447[(3'h5):(3'h5)])));
        end
      else
        begin
          reg2480 <= "adEIXSYEf7DsJJNpIA2";
          for (forvar2481 = (1'h0); (forvar2481 < (2'h2)); forvar2481 = (forvar2481 + (1'h1)))
            begin
              reg2482 <= reg2464;
              reg2483 <= reg2345[(5'h14):(3'h5)];
            end
          reg2484 <= (8'hbd);
          reg2485 = reg2497[(4'h9):(1'h0)];
        end
      reg2500 <= ((8'hae) ^~ "5EyaKImApxWW6FFLXp3R");
    end
  always
    @(posedge clk) begin
      reg2501 <= $unsigned((forvar2320 ?
          "pqNS50NUoTzEKtRxBCck" : $signed((8'h9f))));
      reg2502 = reg2312[(3'h6):(1'h0)];
      reg2503 <= forvar2493[(1'h1):(1'h0)];
      for (forvar2504 = (1'h0); (forvar2504 < (2'h3)); forvar2504 = (forvar2504 + (1'h1)))
        begin
          reg2505 <= ("OYFLK5" ~^ reg2354[(3'h6):(1'h0)]);
          reg2506 <= (~|$unsigned(reg2472));
        end
      reg2507 <= (($unsigned(reg2410) ?
              $unsigned(reg2450[(4'h9):(3'h5)]) : "SK3Z0PEmU8VzbwO0UqB") ?
          {reg2360} : $signed(reg2478[(2'h2):(2'h2)]));
      reg2508 <= ($signed(reg2400[(2'h2):(1'h0)]) ?
          $signed("N0edJ54r4yJKhU8YAQvLHVzY") : wire2285);
    end
  always
    @(posedge clk) begin
      reg2509 <= reg2343;
      reg2510 <= $unsigned(($signed({(reg2421 ? reg2477 : reg2360), reg2395}) ?
          ($signed("2Mbgd7ecn5mpHZwy") ?
              {(reg2394 >> reg2355)} : (+$unsigned(reg2442))) : "tu"));
      for (forvar2511 = (1'h0); (forvar2511 < (2'h3)); forvar2511 = (forvar2511 + (1'h1)))
        begin
          for (forvar2512 = (1'h0); (forvar2512 < (2'h2)); forvar2512 = (forvar2512 + (1'h1)))
            begin
              reg2513 <= reg2414[(4'h9):(4'h8)];
              reg2514 <= (~^(^reg2479));
              reg2515 = reg2295;
              reg2516 <= ($unsigned("mq8ILpctSvLBBhECdcZ8QAy") ^~ (reg2316 && ($signed((reg2419 ?
                  reg2366 : reg2486)) >>> (reg2471[(3'h6):(3'h4)] ?
                  (reg2381 ? reg2338 : reg2461) : (~reg2300)))));
              reg2517 = $signed(((!(!$unsigned(reg2509))) ?
                  $unsigned("SIbpg3zH5trRP9") : "xx6nQIE2bHg5"));
            end
          reg2518 <= "Glymkx";
          for (forvar2519 = (1'h0); (forvar2519 < (3'h4)); forvar2519 = (forvar2519 + (1'h1)))
            begin
              reg2520 <= (&(reg2411[(3'h4):(3'h4)] & ((^~"BxEGf15O1PiOCz3") ?
                  $signed(((8'hb5) ?
                      reg2492 : forvar2380)) : $unsigned(((8'ha0) ^ reg2409)))));
              reg2521 <= reg2467[(1'h0):(1'h0)];
              reg2522 <= (reg2384 <= ({"AQAo",
                  "uI8TQh2z"} ~^ $unsigned($unsigned((8'hb6)))));
              reg2523 <= $unsigned(wire2315);
              reg2524 <= (~|wire2284[(3'h6):(3'h6)]);
            end
          reg2525 <= $signed($unsigned({{(reg2475 ? reg2455 : forvar2322)},
              ($signed(reg2414) ? (~&reg2507) : "uFs15dkJIQ")}));
        end
      reg2526 = $signed(forvar2288);
      for (forvar2527 = (1'h0); (forvar2527 < (3'h5)); forvar2527 = (forvar2527 + (1'h1)))
        begin
          reg2528 <= (+reg2486[(3'h7):(3'h5)]);
          reg2529 <= $signed({(("E" ?
                      (reg2424 ? reg2376 : forvar2380) : $signed(reg2363)) ?
                  "vzmnksKmYvP" : ((reg2337 ? wire2315 : reg2455) ?
                      "VG" : $signed((7'h4c))))});
        end
    end
  assign wire2530 = (($unsigned(((|reg2523) >> (^~reg2498))) ?
                            $signed(reg2459[(5'h10):(1'h0)]) : "MCztp3") ?
                        "DUauVxQWOD" : (^~"q3ayR7X4aP7LhcVriv"));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2090
#(parameter param2277 = (8'h9f), parameter param2278 = param2277)
(y, clk, wire2095, wire2094, wire2093, wire2092, wire2091);
  output wire [(32'ha40):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h1a):(1'h0)] wire2095;
  input wire [(5'h19):(1'h0)] wire2094;
  input wire [(2'h2):(1'h0)] wire2093;
  input wire signed [(4'ha):(1'h0)] wire2092;
  input wire signed [(5'h18):(1'h0)] wire2091;
  reg [(5'h14):(1'h0)] reg2276 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2275 = (1'h0);
  reg [(4'ha):(1'h0)] reg2274 = (1'h0);
  reg [(4'hb):(1'h0)] reg2273 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2272 = (1'h0);
  reg [(3'h5):(1'h0)] reg2271 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2270 = (1'h0);
  reg [(4'hc):(1'h0)] reg2269 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2268 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2267 = (1'h0);
  reg [(5'h16):(1'h0)] reg2266 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2265 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2264 = (1'h0);
  reg [(4'h9):(1'h0)] reg2263 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2262 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2261 = (1'h0);
  reg [(5'h12):(1'h0)] reg2260 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2259 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2258 = (1'h0);
  reg [(4'ha):(1'h0)] reg2257 = (1'h0);
  reg [(4'hd):(1'h0)] reg2256 = (1'h0);
  reg [(5'h17):(1'h0)] reg2255 = (1'h0);
  reg [(5'h10):(1'h0)] reg2254 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2253 = (1'h0);
  reg [(4'ha):(1'h0)] reg2252 = (1'h0);
  reg [(5'h10):(1'h0)] reg2251 = (1'h0);
  reg [(5'h19):(1'h0)] forvar2250 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2249 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2248 = (1'h0);
  reg [(5'h11):(1'h0)] reg2247 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire2246;
  reg [(2'h3):(1'h0)] reg2245 = (1'h0);
  reg [(5'h13):(1'h0)] reg2244 = (1'h0);
  reg [(3'h5):(1'h0)] reg2243 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2242 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2241 = (1'h0);
  reg [(4'hf):(1'h0)] reg2240 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2239 = (1'h0);
  reg [(4'hd):(1'h0)] reg2238 = (1'h0);
  reg [(4'h9):(1'h0)] reg2237 = (1'h0);
  reg [(2'h3):(1'h0)] reg2236 = (1'h0);
  reg [(4'hd):(1'h0)] reg2235 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2234 = (1'h0);
  reg [(3'h7):(1'h0)] reg2233 = (1'h0);
  reg [(4'hf):(1'h0)] reg2232 = (1'h0);
  reg [(4'hf):(1'h0)] reg2231 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2230 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2229 = (1'h0);
  reg [(2'h3):(1'h0)] reg2228 = (1'h0);
  reg [(4'he):(1'h0)] reg2227 = (1'h0);
  reg [(4'hd):(1'h0)] reg2226 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2225 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2224 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2223 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2222 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2221 = (1'h0);
  reg [(4'ha):(1'h0)] reg2220 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2219 = (1'h0);
  reg [(2'h3):(1'h0)] reg2218 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2217 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2216 = (1'h0);
  reg [(4'hc):(1'h0)] reg2215 = (1'h0);
  reg [(5'h10):(1'h0)] reg2214 = (1'h0);
  reg [(4'hb):(1'h0)] reg2213 = (1'h0);
  reg [(5'h10):(1'h0)] reg2212 = (1'h0);
  reg [(5'h13):(1'h0)] reg2211 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2210 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2209 = (1'h0);
  reg [(2'h2):(1'h0)] reg2208 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2207 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2206 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2205 = (1'h0);
  reg [(5'h13):(1'h0)] reg2204 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2203 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2202 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2201 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2200 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire2199;
  reg [(3'h7):(1'h0)] forvar2197 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2196 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2198 = (1'h0);
  reg [(4'h8):(1'h0)] reg2197 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2196 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2195 = (1'h0);
  reg [(4'he):(1'h0)] reg2194 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2193 = (1'h0);
  reg [(5'h19):(1'h0)] forvar2192 = (1'h0);
  reg [(5'h11):(1'h0)] reg2191 = (1'h0);
  reg [(5'h15):(1'h0)] reg2190 = (1'h0);
  reg [(4'hb):(1'h0)] reg2189 = (1'h0);
  reg [(2'h3):(1'h0)] reg2188 = (1'h0);
  reg [(5'h11):(1'h0)] reg2187 = (1'h0);
  reg [(3'h7):(1'h0)] reg2186 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2185 = (1'h0);
  reg [(4'hd):(1'h0)] reg2184 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2183 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2182 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2181 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2180 = (1'h0);
  reg [(4'h8):(1'h0)] reg2179 = (1'h0);
  reg [(3'h6):(1'h0)] reg2178 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2177 = (1'h0);
  reg [(5'h17):(1'h0)] reg2176 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2175 = (1'h0);
  reg [(5'h14):(1'h0)] reg2174 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2173 = (1'h0);
  reg [(5'h15):(1'h0)] reg2172 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2171 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2170 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2169 = (1'h0);
  reg [(5'h17):(1'h0)] reg2168 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2167 = (1'h0);
  reg [(3'h5):(1'h0)] reg2166 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2165 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2164 = (1'h0);
  reg [(4'hb):(1'h0)] reg2163 = (1'h0);
  reg [(5'h13):(1'h0)] reg2162 = (1'h0);
  reg [(3'h7):(1'h0)] reg2161 = (1'h0);
  reg [(5'h13):(1'h0)] reg2160 = (1'h0);
  reg [(4'h9):(1'h0)] reg2159 = (1'h0);
  reg [(2'h2):(1'h0)] reg2158 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2157 = (1'h0);
  reg [(5'h16):(1'h0)] reg2156 = (1'h0);
  reg [(4'h8):(1'h0)] reg2155 = (1'h0);
  reg [(5'h18):(1'h0)] reg2154 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2153 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2152 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2151 = (1'h0);
  reg [(5'h15):(1'h0)] reg2150 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2149 = (1'h0);
  wire [(5'h10):(1'h0)] wire2148;
  wire [(2'h2):(1'h0)] wire2147;
  reg [(3'h6):(1'h0)] reg2146 = (1'h0);
  reg [(5'h17):(1'h0)] reg2145 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2144 = (1'h0);
  wire [(5'h12):(1'h0)] wire2143;
  reg signed [(5'h15):(1'h0)] reg2142 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2141 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2140 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2139 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2138 = (1'h0);
  reg [(4'hf):(1'h0)] reg2137 = (1'h0);
  reg [(5'h17):(1'h0)] reg2136 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2135 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2134 = (1'h0);
  reg [(5'h12):(1'h0)] forvar2133 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2132 = (1'h0);
  reg [(5'h19):(1'h0)] reg2131 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2130 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2129 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2128 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2127 = (1'h0);
  reg [(2'h3):(1'h0)] reg2126 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2125 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2124 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2123 = (1'h0);
  reg [(2'h3):(1'h0)] reg2122 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2121 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2120 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2101 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2098 = (1'h0);
  reg [(3'h4):(1'h0)] reg2097 = (1'h0);
  reg [(5'h11):(1'h0)] reg2119 = (1'h0);
  reg [(3'h7):(1'h0)] reg2118 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2117 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2116 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2115 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2114 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2113 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2112 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2111 = (1'h0);
  reg [(5'h15):(1'h0)] reg2110 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2109 = (1'h0);
  reg [(4'he):(1'h0)] reg2108 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2107 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2106 = (1'h0);
  reg [(4'he):(1'h0)] reg2105 = (1'h0);
  reg [(4'hd):(1'h0)] reg2104 = (1'h0);
  reg [(5'h19):(1'h0)] reg2103 = (1'h0);
  reg [(3'h5):(1'h0)] reg2102 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2101 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2100 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2099 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2098 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2097 = (1'h0);
  reg [(4'hc):(1'h0)] reg2096 = (1'h0);
  assign y = {reg2276,
                 forvar2275,
                 reg2274,
                 reg2273,
                 reg2272,
                 reg2271,
                 reg2270,
                 reg2269,
                 reg2268,
                 forvar2267,
                 reg2266,
                 reg2265,
                 forvar2264,
                 reg2263,
                 reg2262,
                 forvar2261,
                 reg2260,
                 reg2259,
                 reg2258,
                 reg2257,
                 reg2256,
                 reg2255,
                 reg2254,
                 forvar2253,
                 reg2252,
                 reg2251,
                 forvar2250,
                 reg2249,
                 forvar2248,
                 reg2247,
                 wire2246,
                 reg2245,
                 reg2244,
                 reg2243,
                 reg2242,
                 reg2241,
                 reg2240,
                 reg2239,
                 reg2238,
                 reg2237,
                 reg2236,
                 reg2235,
                 forvar2234,
                 reg2233,
                 reg2232,
                 reg2231,
                 reg2230,
                 reg2229,
                 reg2228,
                 reg2227,
                 reg2226,
                 reg2225,
                 reg2224,
                 forvar2223,
                 reg2222,
                 forvar2221,
                 reg2220,
                 reg2219,
                 reg2218,
                 reg2217,
                 reg2216,
                 reg2215,
                 reg2214,
                 reg2213,
                 reg2212,
                 reg2211,
                 forvar2210,
                 reg2209,
                 reg2208,
                 reg2207,
                 reg2206,
                 reg2205,
                 reg2204,
                 reg2203,
                 reg2202,
                 forvar2201,
                 forvar2200,
                 wire2199,
                 forvar2197,
                 reg2196,
                 reg2198,
                 reg2197,
                 forvar2196,
                 reg2195,
                 reg2194,
                 reg2193,
                 forvar2192,
                 reg2191,
                 reg2190,
                 reg2189,
                 reg2188,
                 reg2187,
                 reg2186,
                 reg2185,
                 reg2184,
                 reg2183,
                 forvar2182,
                 reg2181,
                 forvar2180,
                 reg2179,
                 reg2178,
                 forvar2177,
                 reg2176,
                 reg2175,
                 reg2174,
                 reg2173,
                 reg2172,
                 forvar2171,
                 reg2170,
                 reg2169,
                 reg2168,
                 forvar2167,
                 reg2166,
                 forvar2165,
                 reg2164,
                 reg2163,
                 reg2162,
                 reg2161,
                 reg2160,
                 reg2159,
                 reg2158,
                 reg2157,
                 reg2156,
                 reg2155,
                 reg2154,
                 forvar2153,
                 forvar2152,
                 reg2151,
                 reg2150,
                 reg2149,
                 wire2148,
                 wire2147,
                 reg2146,
                 reg2145,
                 reg2144,
                 wire2143,
                 reg2142,
                 reg2141,
                 reg2140,
                 reg2139,
                 reg2138,
                 reg2137,
                 reg2136,
                 reg2135,
                 reg2134,
                 forvar2133,
                 reg2132,
                 reg2131,
                 reg2130,
                 reg2129,
                 forvar2128,
                 reg2127,
                 reg2126,
                 forvar2125,
                 reg2124,
                 reg2123,
                 reg2122,
                 reg2121,
                 forvar2120,
                 reg2101,
                 forvar2098,
                 reg2097,
                 reg2119,
                 reg2118,
                 reg2117,
                 reg2116,
                 reg2115,
                 reg2114,
                 reg2113,
                 reg2112,
                 reg2111,
                 reg2110,
                 forvar2109,
                 reg2108,
                 forvar2107,
                 reg2106,
                 reg2105,
                 reg2104,
                 reg2103,
                 reg2102,
                 forvar2101,
                 reg2100,
                 reg2099,
                 reg2098,
                 forvar2097,
                 reg2096,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg2096 <= (wire2093[(1'h0):(1'h0)] ^~ {(|$signed((wire2092 ?
              (8'ha9) : wire2091)))});
      if ({"punnNnroBMJ0SfMwuEcZUldD", (+wire2095)})
        begin
          for (forvar2097 = (1'h0); (forvar2097 < (1'h0)); forvar2097 = (forvar2097 + (1'h1)))
            begin
              reg2098 <= (|reg2096[(4'hc):(3'h7)]);
              reg2099 <= ($unsigned((($signed(reg2098) ?
                  wire2091[(3'h5):(1'h0)] : wire2095[(1'h1):(1'h1)]) | (+$signed(forvar2097)))) != (reg2096 ?
                  (~|(~|wire2094)) : ((8'ha7) <= {wire2094,
                      (reg2098 ? wire2092 : forvar2097)})));
              reg2100 <= $signed((-wire2092));
              for (forvar2101 = (1'h0); (forvar2101 < (2'h3)); forvar2101 = (forvar2101 + (1'h1)))
                begin
                  reg2102 <= "4LJOO80JR3r";
                  reg2103 <= "SwIO351A0I";
                  reg2104 <= $unsigned((^reg2096[(1'h1):(1'h1)]));
                  reg2105 <= ($signed(reg2098[(5'h11):(1'h0)]) | $unsigned($signed({"MGQb3dHqqJykVdP"})));
                end
            end
          reg2106 <= (~&{$unsigned("xzG96bSohTsYlOXXsW3HlrmJ")});
          for (forvar2107 = (1'h0); (forvar2107 < (3'h5)); forvar2107 = (forvar2107 + (1'h1)))
            begin
              reg2108 <= (~|"SyEP2E6BGBDrIz");
              for (forvar2109 = (1'h0); (forvar2109 < (3'h5)); forvar2109 = (forvar2109 + (1'h1)))
                begin
                  reg2110 = $signed(reg2099[(1'h1):(1'h1)]);
                  reg2111 <= reg2108[(4'hb):(3'h5)];
                  reg2112 <= (^~$signed((+($unsigned(reg2102) ?
                      reg2103[(4'hb):(4'h9)] : ""))));
                  reg2113 <= ((+"AIi7m6dNseyl") ?
                      ({forvar2109[(1'h1):(1'h0)]} ?
                          (|{reg2105[(4'hb):(3'h7)]}) : (reg2103[(5'h12):(1'h1)] ~^ (wire2092[(4'ha):(4'h9)] ^~ $signed(wire2093)))) : forvar2101);
                end
              reg2114 <= forvar2101[(3'h4):(2'h2)];
              reg2115 <= (((~&(reg2114[(1'h0):(1'h0)] ?
                  "i" : $unsigned(reg2103))) >>> reg2106) > ({$unsigned($signed(forvar2097))} << {"bPsGb3YJbG1bVFssubItX",
                  $unsigned((wire2093 <= reg2096))}));
              reg2116 <= reg2114[(5'h11):(4'h9)];
              reg2117 <= wire2091[(4'hf):(3'h7)];
            end
          reg2118 <= $unsigned(reg2112[(4'h8):(3'h4)]);
          reg2119 <= (("a0hqDaksQ1Y" < "Eh85Ih") >> ((8'ha3) ?
              $signed(($signed(reg2105) ?
                  (reg2118 ? reg2098 : reg2108) : {reg2096,
                      (8'ha4)})) : {$signed({wire2094}),
                  {(7'h4b), $signed(wire2094)}}));
        end
      else
        begin
          reg2097 <= (reg2114 ?
              $unsigned(reg2116) : $signed((~{$unsigned(reg2099)})));
          for (forvar2098 = (1'h0); (forvar2098 < (2'h3)); forvar2098 = (forvar2098 + (1'h1)))
            begin
              reg2099 <= "v5TnWdh5cr";
              reg2100 <= ($signed(({(reg2108 ? reg2103 : forvar2097),
                          {reg2097, reg2100}} ?
                      wire2092[(3'h5):(2'h3)] : (forvar2109[(2'h2):(1'h0)] ?
                          $signed(forvar2098) : $unsigned(forvar2097)))) ?
                  {({$unsigned(forvar2097),
                          $unsigned(forvar2109)} <= reg2097)} : reg2114);
              reg2101 <= (reg2112[(3'h7):(3'h6)] ?
                  "Qi89Z1hmAioAf" : {{(|(^reg2108))}});
              reg2102 <= (~((reg2118[(1'h0):(1'h0)] ~^ (&(^~reg2102))) ?
                  $unsigned((~&wire2094)) : ($signed(reg2099[(1'h1):(1'h0)]) ?
                      {{reg2115}} : $unsigned((wire2092 ^ reg2115)))));
            end
          reg2103 = reg2102[(1'h0):(1'h0)];
          reg2104 = reg2113[(3'h5):(3'h5)];
        end
      for (forvar2120 = (1'h0); (forvar2120 < (2'h2)); forvar2120 = (forvar2120 + (1'h1)))
        begin
          reg2121 = "YzZBkumTbMMqrqB9tMCZdtra";
        end
      reg2122 <= (|reg2102[(2'h2):(1'h1)]);
      reg2123 <= $signed(((~|reg2119[(1'h0):(1'h0)]) ?
          ($signed($unsigned(reg2119)) != (8'ha8)) : wire2091[(4'hd):(3'h6)]));
    end
  always
    @(posedge clk) begin
      reg2124 <= $signed(forvar2098[(4'h8):(4'h8)]);
      for (forvar2125 = (1'h0); (forvar2125 < (2'h3)); forvar2125 = (forvar2125 + (1'h1)))
        begin
          reg2126 <= $unsigned(reg2097[(1'h0):(1'h0)]);
          reg2127 = ({reg2099,
              $unsigned($unsigned(reg2113[(5'h17):(4'h8)]))} >= "gxhHmHak");
          for (forvar2128 = (1'h0); (forvar2128 < (3'h5)); forvar2128 = (forvar2128 + (1'h1)))
            begin
              reg2129 <= $signed("cBtF4BG");
              reg2130 <= $signed(reg2112);
              reg2131 = reg2097;
              reg2132 <= "LlGhvwH19rZawELElc";
              for (forvar2133 = (1'h0); (forvar2133 < (3'h5)); forvar2133 = (forvar2133 + (1'h1)))
                begin
                  reg2134 <= $unsigned(reg2100[(2'h3):(2'h2)]);
                  reg2135 <= ("obcUMbvJQID5x6TzN" ? ("8XrZ" <= "TD") : (8'ha4));
                  reg2136 <= reg2096;
                  reg2137 <= (reg2117 + $signed("mbQzEN4ERkYFO6Plf"));
                  reg2138 <= reg2110[(3'h4):(2'h3)];
                end
            end
          reg2139 <= $unsigned(({"uqYSfTfWM8IZq",
                  ((reg2117 + reg2110) ?
                      (wire2095 ? reg2124 : (7'h46)) : "Hk8ZGMDl")} ?
              $unsigned({"ePR91SW", {reg2111, reg2119}}) : "FQhqxTSCfZecWHZL"));
          reg2140 <= {$unsigned($signed(((~|reg2130) != forvar2101[(4'h8):(1'h0)]))),
              $unsigned(({""} ? (!(reg2132 || reg2106)) : reg2106))};
          reg2141 <= (("X8IEPA4F4Ng4ObtK3EBp" ?
              ((reg2115 ?
                  reg2140[(4'hf):(4'h9)] : (reg2112 ?
                      reg2137 : reg2139)) != (reg2123[(4'h8):(2'h2)] <= $unsigned(forvar2133))) : reg2115) >>> "26KafXLagYkrtQLdhZ2F7Sh");
        end
      reg2142 = {{$unsigned("tq"), ($unsigned(reg2138) ~^ reg2130)},
          ("QGACMJ1vOFXfdUtHRKurI" >>> (!$unsigned((wire2092 <<< reg2099))))};
    end
  assign wire2143 = (8'hb2);
  always
    @(posedge clk) begin
      reg2144 = $signed($signed((^($unsigned(reg2101) >= $signed(reg2105)))));
      reg2145 <= "rFpWvBGbipk93sf4gEBeY";
      reg2146 = reg2118;
    end
  assign wire2147 = $unsigned(forvar2128);
  assign wire2148 = $signed($unsigned(reg2142));
  always
    @(posedge clk) begin
      reg2149 <= $unsigned($unsigned((|forvar2097)));
      reg2150 <= reg2119;
      reg2151 <= "aK";
      for (forvar2152 = (1'h0); (forvar2152 < (1'h1)); forvar2152 = (forvar2152 + (1'h1)))
        begin
          for (forvar2153 = (1'h0); (forvar2153 < (1'h1)); forvar2153 = (forvar2153 + (1'h1)))
            begin
              reg2154 <= reg2150;
              reg2155 <= reg2099[(4'he):(3'h5)];
              reg2156 = ((-reg2124) >> (~|$signed(($unsigned((8'ha3)) ?
                  "BVYb6Raix9zz9mcP45rKrio" : "u70k6R3DtQrNLLr"))));
            end
        end
      reg2157 <= {{"Y9Yo4UlS", forvar2098[(3'h7):(1'h0)]},
          $signed(reg2136[(4'hc):(3'h4)])};
    end
  always
    @(posedge clk) begin
      reg2158 = ((^~wire2093[(2'h2):(1'h1)]) ^~ ($signed($unsigned(reg2111[(5'h14):(4'hf)])) ?
          ($signed(((8'ha2) == (8'ha7))) ?
              $signed((reg2141 ?
                  reg2126 : (8'h9f))) : wire2092[(1'h0):(1'h0)]) : $unsigned(reg2157[(4'hd):(4'ha)])));
      reg2159 = "NR2";
      reg2160 <= (&((~$signed("mJ6BfrVvWldOl")) ?
          "ytZ5ZmBIu6mni4nhTRgRy5P" : reg2156));
      reg2161 <= $unsigned(($unsigned((&(reg2135 ? reg2115 : forvar2097))) ?
          wire2091[(5'h15):(5'h10)] : $unsigned($signed((reg2150 ?
              reg2132 : reg2124)))));
    end
  always
    @(posedge clk) begin
      reg2162 = ($unsigned($signed(wire2093)) ?
          (~("GQ9yWEtJYq" ?
              (~^$unsigned((7'h43))) : ($signed(forvar2133) ?
                  $signed(reg2112) : reg2118))) : ("u9GxK2ed25" ~^ $signed(((reg2146 ?
                  forvar2128 : reg2160) ?
              $unsigned(wire2094) : "sOhEnlFW"))));
      reg2163 <= {(reg2117 >= "w5N")};
      reg2164 = $signed($signed((reg2138[(3'h7):(1'h1)] ?
          {(reg2158 ? reg2149 : reg2116),
              (forvar2097 ? forvar2153 : reg2162)} : {"gmB5mDNgBnigApR"})));
      for (forvar2165 = (1'h0); (forvar2165 < (1'h0)); forvar2165 = (forvar2165 + (1'h1)))
        begin
          reg2166 <= reg2121;
          for (forvar2167 = (1'h0); (forvar2167 < (3'h5)); forvar2167 = (forvar2167 + (1'h1)))
            begin
              reg2168 <= {(7'h48)};
              reg2169 <= {(+(($unsigned(reg2166) >> (forvar2153 >>> reg2104)) ?
                      reg2157[(5'h15):(4'hf)] : ($signed(reg2137) ?
                          ((8'hbc) && reg2111) : {reg2151, reg2166})))};
              reg2170 <= reg2097;
              for (forvar2171 = (1'h0); (forvar2171 < (2'h2)); forvar2171 = (forvar2171 + (1'h1)))
                begin
                  reg2172 <= $signed($signed($signed((reg2156[(3'h7):(3'h7)] && {reg2110}))));
                  reg2173 <= reg2144[(4'ha):(3'h5)];
                  reg2174 <= $signed(forvar2152);
                  reg2175 <= $signed("UPPL7PAB6rqbMB68Ng0cMdrET");
                  reg2176 = "muagyVPBi9";
                end
              for (forvar2177 = (1'h0); (forvar2177 < (3'h4)); forvar2177 = (forvar2177 + (1'h1)))
                begin
                  reg2178 <= {({reg2175} ?
                          ($unsigned($unsigned((8'haf))) ?
                              reg2106[(4'h8):(3'h6)] : $unsigned((&reg2122))) : (reg2134[(3'h7):(3'h7)] ?
                              {(reg2131 ? forvar2125 : (8'hb7)),
                                  $unsigned(reg2172)} : "bcOVUVHFkD"))};
                  reg2179 <= ($unsigned(($unsigned((!reg2102)) ?
                      $signed(((8'ha3) ?
                          reg2116 : reg2132)) : ($unsigned(reg2112) > "ry1WYJhMQ"))) == $signed("WTBtUSx"));
                end
            end
          for (forvar2180 = (1'h0); (forvar2180 < (1'h1)); forvar2180 = (forvar2180 + (1'h1)))
            begin
              reg2181 <= ($signed(reg2178) ?
                  ("RIhFBKBcY574Z8qz" ?
                      forvar2101 : (7'h4c)) : ((&(reg2170[(2'h2):(2'h2)] + {(8'ha2)})) ?
                      $signed(forvar2097) : $signed((8'hb4))));
              for (forvar2182 = (1'h0); (forvar2182 < (3'h5)); forvar2182 = (forvar2182 + (1'h1)))
                begin
                  reg2183 <= reg2103[(3'h7):(3'h4)];
                  reg2184 <= $unsigned(forvar2120);
                  reg2185 <= {forvar2177, (!reg2169)};
                  reg2186 <= (+"c4fupS4ISbUUswWTiG");
                  reg2187 <= reg2158;
                end
              reg2188 <= reg2134[(4'hc):(4'hb)];
              reg2189 <= $unsigned($unsigned($signed((((8'hb0) * forvar2098) ?
                  reg2188[(1'h0):(1'h0)] : (!reg2173)))));
              reg2190 <= reg2134;
            end
          reg2191 <= ((-(+("JT86m1ev" ?
              (~|reg2144) : $unsigned(forvar2153)))) ^ "");
          for (forvar2192 = (1'h0); (forvar2192 < (1'h0)); forvar2192 = (forvar2192 + (1'h1)))
            begin
              reg2193 <= reg2160[(5'h13):(3'h5)];
            end
        end
      if ("yVQQ4GsC4SGlxe2oVcY017R")
        begin
          reg2194 = reg2186;
          reg2195 = ($signed(($signed($unsigned(reg2105)) <= {"WQC7iEv3h7SJqY9rgAfZOqA"})) > reg2110);
          for (forvar2196 = (1'h0); (forvar2196 < (3'h4)); forvar2196 = (forvar2196 + (1'h1)))
            begin
              reg2197 = ("rcxXZSGDMF2B1009MCbqFV3E" | reg2150);
            end
          reg2198 <= (((~&{{reg2178, reg2140},
                  forvar2120}) >> (($signed(reg2183) <<< "JtzGLUauMzMywx2tV") ?
                  (~|$unsigned(reg2140)) : ((forvar2177 >>> reg2194) < $signed(wire2091)))) ?
              reg2138 : ((+{(reg2186 ? reg2113 : reg2102)}) ?
                  "8p0G0yxaJWnS" : ($unsigned((reg2178 << reg2135)) != ((reg2142 - (8'hbf)) ?
                      reg2175 : $signed(reg2116)))));
        end
      else
        begin
          reg2194 <= $signed((&{(|reg2131),
              ((^reg2169) ? "H9sbLME05" : reg2175[(1'h0):(1'h0)])}));
          reg2195 <= (($signed($signed($signed((8'ha7)))) ?
                  ({{forvar2152}} ^~ reg2130[(3'h6):(1'h0)]) : reg2188) ?
              reg2105 : forvar2167[(2'h2):(2'h2)]);
          reg2196 <= (~|"1JgcIoYP");
          for (forvar2197 = (1'h0); (forvar2197 < (1'h0)); forvar2197 = (forvar2197 + (1'h1)))
            begin
              reg2198 <= (8'ha4);
            end
        end
    end
  assign wire2199 = forvar2192[(5'h10):(4'h9)];
  always
    @(posedge clk) begin
      for (forvar2200 = (1'h0); (forvar2200 < (2'h3)); forvar2200 = (forvar2200 + (1'h1)))
        begin
          for (forvar2201 = (1'h0); (forvar2201 < (2'h3)); forvar2201 = (forvar2201 + (1'h1)))
            begin
              reg2202 <= reg2116;
              reg2203 <= $signed(("sZrCzYp9lD7MsSPQPW" ?
                  reg2116[(4'hd):(2'h3)] : $unsigned(reg2170)));
              reg2204 <= ((-({reg2121,
                  (-(8'haa))} || reg2113[(5'h1a):(1'h1)])) ^ $signed(forvar2201));
              reg2205 <= (($unsigned($unsigned(((8'h9f) << reg2157))) & "F2WICcrrsST9YrKITD") ?
                  (($unsigned($unsigned(forvar2128)) ? reg2134 : reg2185) ?
                      reg2169[(5'h10):(4'hf)] : $signed(reg2105)) : "MqRp");
              reg2206 = ((reg2181[(4'h8):(3'h4)] ?
                  (((reg2106 ? reg2134 : reg2106) >> reg2136) ?
                      $unsigned(reg2168) : reg2175) : (-forvar2098)) | "lLBhbI3HYXvBTVz7q");
              reg2207 <= $unsigned((forvar2107[(3'h7):(3'h6)] ?
                  $unsigned($signed({reg2198, (7'h40)})) : reg2146));
            end
          reg2208 <= "D0yFgmNyRrhtzzHuYfepF1c";
          reg2209 <= ("hFJ" << $unsigned({(~^wire2148[(3'h7):(3'h4)]),
              "5qbakiFWsFmycgcFwpNvX6BN"}));
        end
      for (forvar2210 = (1'h0); (forvar2210 < (2'h3)); forvar2210 = (forvar2210 + (1'h1)))
        begin
          reg2211 = reg2207[(2'h3):(2'h2)];
        end
    end
  always
    @(posedge clk) begin
      reg2212 <= {reg2191};
      reg2213 = reg2149;
      reg2214 = forvar2200;
    end
  always
    @(posedge clk) begin
      reg2215 <= $unsigned((("5my7zMlQrCuKTLLmadm" + reg2098) != $unsigned($unsigned((^reg2202)))));
      reg2216 = ((reg2184[(4'h8):(1'h0)] ?
          (~&reg2198) : reg2127[(1'h0):(1'h0)]) & $unsigned($signed((~|$unsigned(reg2204)))));
      reg2217 <= (("tY0ARLQiIWeJ6PYnvzhG4DC54" == $unsigned((!{wire2095}))) ?
          reg2150[(3'h7):(3'h4)] : wire2092);
      reg2218 <= (&(~|(~|$signed((!forvar2200)))));
    end
  always
    @(posedge clk) begin
      reg2219 <= reg2099[(3'h7):(3'h7)];
      reg2220 <= (^~$unsigned({{$unsigned(forvar2098)},
          (forvar2182[(3'h7):(3'h4)] >= (8'hb9))}));
    end
  always
    @(posedge clk) begin
      for (forvar2221 = (1'h0); (forvar2221 < (3'h4)); forvar2221 = (forvar2221 + (1'h1)))
        begin
          reg2222 <= reg2163;
          for (forvar2223 = (1'h0); (forvar2223 < (2'h2)); forvar2223 = (forvar2223 + (1'h1)))
            begin
              reg2224 <= $signed("9pZ1rOhJF5Vxn51Jf66Ba");
            end
          reg2225 <= $unsigned($signed(reg2116));
          reg2226 <= {$signed($unsigned((((8'hbe) ?
                  reg2187 : (8'hbf)) == $unsigned(reg2115))))};
          if (reg2136[(2'h2):(1'h1)])
            begin
              reg2227 = $signed({$signed(("X2JE" ?
                      forvar2120[(2'h3):(1'h1)] : reg2166[(1'h1):(1'h0)]))});
              reg2228 <= "DsP8KWvkHhXlnG8cXiI";
              reg2229 <= reg2208[(1'h1):(1'h0)];
            end
          else
            begin
              reg2227 <= ("rhH1YK2IPhGQFKRJFRqqC" ^ reg2169[(4'h9):(3'h7)]);
              reg2228 <= forvar2152[(3'h4):(2'h2)];
              if (("o1zXfBiO" >>> ("QHiyQ7wHq1J" ?
                  {{{reg2168}},
                      reg2166[(1'h0):(1'h0)]} : reg2151[(2'h2):(1'h1)])))
                begin
                  reg2229 <= $unsigned(reg2103[(4'hc):(1'h1)]);
                  reg2230 <= {$unsigned(reg2197[(1'h1):(1'h1)]),
                      (($signed(reg2137[(4'hc):(2'h2)]) * (~^$signed(reg2146))) ?
                          reg2215 : (!"k"))};
                  reg2231 = ({forvar2192} ?
                      $signed(reg2115[(1'h0):(1'h0)]) : (("YkPMdVI" ?
                              $signed((reg2136 ?
                                  reg2175 : reg2102)) : reg2127) ?
                          ("5Ek0R09" ?
                              reg2151 : ("P8h" != $signed(reg2181))) : ({(~|reg2160),
                              (forvar2200 ?
                                  reg2123 : (7'h47))} || $signed(((7'h46) ?
                              forvar2101 : (8'ha9))))));
                  reg2232 <= "m8YBmitNm4dzH";
                  reg2233 <= (+$unsigned((~^reg2179)));
                end
              else
                begin
                  reg2229 = $unsigned(reg2174);
                  reg2230 <= (-(wire2148[(4'ha):(3'h7)] ?
                      "0dyZ9N3CFPIybbNWZycowUA" : reg2151));
                  reg2231 <= reg2138;
                  reg2232 = ("vhofsRIDmkRSc" == reg2172[(2'h2):(2'h2)]);
                end
              for (forvar2234 = (1'h0); (forvar2234 < (3'h5)); forvar2234 = (forvar2234 + (1'h1)))
                begin
                  reg2235 = forvar2197;
                  reg2236 <= $unsigned(reg2231);
                  reg2237 <= (("prk9rEsJygGcCfttyM18b" ?
                      $unsigned(reg2204) : reg2149[(1'h1):(1'h1)]) <= "JNKoHQMdyntb5oZ");
                  reg2238 <= (8'hb3);
                  reg2239 <= ((reg2183[(4'h8):(1'h0)] + ($signed(((8'hbb) >> (8'ha9))) - $unsigned(((8'hb3) > reg2098)))) ?
                      $signed(reg2158[(1'h1):(1'h0)]) : $unsigned(((!(reg2101 ?
                          reg2121 : (8'ha3))) ~^ $unsigned((reg2190 ?
                          wire2199 : reg2217)))));
                  reg2240 <= $signed((~&$signed("JW1AQHpdMTRCG2gOrG37yr")));
                end
            end
          reg2241 <= "10zUxQlQud8UKJUp8w6lBeJLO";
        end
      reg2242 <= {(((|$unsigned(wire2143)) - wire2092[(4'ha):(3'h6)]) ?
              "rMvp" : (^~$signed((reg2226 <= reg2169))))};
      reg2243 = "QvFq0avc6QUYKlt";
      reg2244 <= "ieNdiR78ZdmkDluEUyDcZRu";
      reg2245 <= reg2214[(4'he):(3'h6)];
    end
  assign wire2246 = ("Cy7Utp3sXNo2M709hO1NUYaIU" ^ $unsigned((("cHWYrE" + (forvar2152 * reg2237)) ^ "tzKaSHUZz7g85qJ7KuhcFuG5")));
  always
    @(posedge clk) begin
      reg2247 <= reg2185;
    end
  always
    @(posedge clk) begin
      for (forvar2248 = (1'h0); (forvar2248 < (3'h5)); forvar2248 = (forvar2248 + (1'h1)))
        begin
          reg2249 <= reg2174;
          for (forvar2250 = (1'h0); (forvar2250 < (1'h0)); forvar2250 = (forvar2250 + (1'h1)))
            begin
              reg2251 <= (&(8'haf));
              reg2252 <= reg2240;
              for (forvar2253 = (1'h0); (forvar2253 < (3'h5)); forvar2253 = (forvar2253 + (1'h1)))
                begin
                  reg2254 <= $signed($signed(""));
                  reg2255 <= $signed(reg2155);
                  reg2256 = reg2244[(4'he):(3'h4)];
                  reg2257 <= (!$signed($unsigned(("ih53drqL3sglkHsA6MRgsnR" ?
                      (forvar2153 ? reg2116 : reg2103) : "Xmo9G10acFRDhn7N"))));
                  reg2258 = $unsigned($signed((((reg2164 ?
                      forvar2171 : reg2174) > "ZqoSYGLm") ~^ "hKXlgoroK4KDA9")));
                  reg2259 = $signed(reg2158);
                end
              reg2260 <= {(&((^(reg2186 ^ reg2208)) ?
                      "qtiD05J" : {$signed((8'hbb)), $signed(reg2114)}))};
            end
          for (forvar2261 = (1'h0); (forvar2261 < (1'h1)); forvar2261 = (forvar2261 + (1'h1)))
            begin
              reg2262 <= $signed($unsigned((^"tS")));
              reg2263 <= ("siL3tlEQ1NuWRh" | $signed((!reg2166)));
              for (forvar2264 = (1'h0); (forvar2264 < (2'h2)); forvar2264 = (forvar2264 + (1'h1)))
                begin
                  reg2265 <= forvar2120;
                  reg2266 = "nIn9yO";
                end
              for (forvar2267 = (1'h0); (forvar2267 < (2'h2)); forvar2267 = (forvar2267 + (1'h1)))
                begin
                  reg2268 <= (~|"6N1rqw4v8EMlNoJwdTiJkNk");
                  reg2269 = (reg2266 || $signed($signed(reg2162[(4'hd):(4'hb)])));
                  reg2270 <= ("dg6EFiJnedbrAWAaznWlK" > (~&("1UtktBnJR" && $unsigned($unsigned(reg2140)))));
                  reg2271 <= "7cGVexzZTXz580t2PFYXPNCl";
                end
              reg2272 <= $unsigned((((|$signed(reg2215)) ?
                  "irlah1Mf92abQgho5S4ayIb" : $unsigned(((8'hb2) ?
                      reg2112 : (8'hae)))) == (((reg2265 ?
                      forvar2250 : (8'hbf)) | reg2216) ?
                  {$signed(reg2172)} : $signed(reg2121))));
            end
          reg2273 <= (reg2112 ? forvar2098[(2'h2):(1'h1)] : "JVlRqgYeC3XZD3");
        end
      reg2274 <= (8'h9e);
    end
  always
    @(posedge clk) begin
      for (forvar2275 = (1'h0); (forvar2275 < (2'h3)); forvar2275 = (forvar2275 + (1'h1)))
        begin
          reg2276 <= (~^$unsigned(""));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1914  (y, clk, wire1918, wire1917, wire1916, wire1915);
  output wire [(32'h848):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h17):(1'h0)] wire1918;
  input wire signed [(2'h2):(1'h0)] wire1917;
  input wire signed [(3'h7):(1'h0)] wire1916;
  input wire signed [(4'hd):(1'h0)] wire1915;
  reg [(5'h17):(1'h0)] reg2067 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2066 = (1'h0);
  reg [(4'ha):(1'h0)] reg2065 = (1'h0);
  reg [(5'h18):(1'h0)] reg2064 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2063 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2062 = (1'h0);
  reg [(4'h8):(1'h0)] reg2061 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2060 = (1'h0);
  reg [(3'h6):(1'h0)] reg2059 = (1'h0);
  reg [(5'h14):(1'h0)] reg2058 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2057 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2056 = (1'h0);
  reg [(4'he):(1'h0)] reg2055 = (1'h0);
  reg [(5'h13):(1'h0)] reg2054 = (1'h0);
  reg [(4'h9):(1'h0)] reg2053 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2052 = (1'h0);
  reg [(5'h13):(1'h0)] reg2051 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2050 = (1'h0);
  reg [(3'h5):(1'h0)] reg2049 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2048 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2047 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2046 = (1'h0);
  reg [(4'h8):(1'h0)] reg2045 = (1'h0);
  reg [(4'ha):(1'h0)] reg2044 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2043 = (1'h0);
  wire [(3'h6):(1'h0)] wire2042;
  reg [(5'h17):(1'h0)] reg2041 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2040 = (1'h0);
  reg [(5'h12):(1'h0)] forvar2039 = (1'h0);
  reg [(5'h10):(1'h0)] reg2038 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2037 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2036 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2035 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2034 = (1'h0);
  reg [(4'hf):(1'h0)] reg2033 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2032 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2031 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2030 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2029 = (1'h0);
  reg [(5'h10):(1'h0)] reg2028 = (1'h0);
  reg [(5'h15):(1'h0)] reg2027 = (1'h0);
  reg [(2'h3):(1'h0)] reg2026 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2025 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2024 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2023 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2022 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2021 = (1'h0);
  reg [(4'ha):(1'h0)] reg2020 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2019 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2018 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2017 = (1'h0);
  reg [(4'hb):(1'h0)] reg2016 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2015 = (1'h0);
  reg [(4'h9):(1'h0)] reg2014 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2013 = (1'h0);
  wire signed [(4'he):(1'h0)] wire2012;
  reg signed [(2'h3):(1'h0)] reg2011 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2010 = (1'h0);
  wire [(4'h9):(1'h0)] wire2009;
  reg [(3'h6):(1'h0)] reg2008 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2007 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2006 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2005 = (1'h0);
  wire [(4'hf):(1'h0)] wire2004;
  reg [(3'h6):(1'h0)] reg2003 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2002 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2001 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2000 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1999 = (1'h0);
  reg [(5'h17):(1'h0)] reg1998 = (1'h0);
  reg [(4'ha):(1'h0)] reg1993 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1988 = (1'h0);
  reg [(5'h11):(1'h0)] reg1997 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1996 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1995 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1994 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1993 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1992 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1991 = (1'h0);
  reg [(5'h11):(1'h0)] reg1990 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1989 = (1'h0);
  reg [(3'h4):(1'h0)] reg1988 = (1'h0);
  reg [(3'h6):(1'h0)] reg1987 = (1'h0);
  reg [(5'h19):(1'h0)] reg1986 = (1'h0);
  reg [(3'h4):(1'h0)] reg1985 = (1'h0);
  reg [(4'h8):(1'h0)] reg1984 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1983 = (1'h0);
  reg [(4'h8):(1'h0)] reg1982 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1981 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1980 = (1'h0);
  reg [(5'h12):(1'h0)] reg1979 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1978 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1977 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1976 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1975 = (1'h0);
  reg [(5'h15):(1'h0)] reg1974 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1973 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1972 = (1'h0);
  reg [(4'hb):(1'h0)] reg1971 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1970 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1969 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1968 = (1'h0);
  reg [(4'h9):(1'h0)] reg1967 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1966 = (1'h0);
  reg [(5'h17):(1'h0)] reg1965 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1964 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1963 = (1'h0);
  reg [(4'hc):(1'h0)] reg1962 = (1'h0);
  reg [(5'h19):(1'h0)] reg1961 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1960 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1959 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1958 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1957 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1956 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1955 = (1'h0);
  reg [(5'h15):(1'h0)] reg1954 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1953 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1952 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1951 = (1'h0);
  reg [(2'h2):(1'h0)] reg1950 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1949 = (1'h0);
  reg [(4'h8):(1'h0)] reg1948 = (1'h0);
  reg [(4'ha):(1'h0)] reg1947 = (1'h0);
  reg [(3'h7):(1'h0)] reg1946 = (1'h0);
  reg [(5'h18):(1'h0)] reg1945 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1944 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1943 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1942 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1941 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1940 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1939 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1938 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1937 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1936 = (1'h0);
  reg [(4'hc):(1'h0)] reg1935 = (1'h0);
  reg [(5'h17):(1'h0)] reg1934 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1933 = (1'h0);
  reg [(5'h10):(1'h0)] reg1932 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1931 = (1'h0);
  reg [(5'h18):(1'h0)] reg1930 = (1'h0);
  reg [(2'h3):(1'h0)] reg1929 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1928 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1927 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1927 = (1'h0);
  reg [(5'h14):(1'h0)] reg1926 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1925 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1924 = (1'h0);
  reg [(5'h11):(1'h0)] reg1923 = (1'h0);
  reg [(4'hd):(1'h0)] reg1922 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1921 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1920 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1919 = (1'h0);
  assign y = {reg2067,
                 reg2066,
                 reg2065,
                 reg2064,
                 reg2063,
                 reg2062,
                 reg2061,
                 reg2060,
                 reg2059,
                 reg2058,
                 forvar2057,
                 reg2056,
                 reg2055,
                 reg2054,
                 reg2053,
                 reg2052,
                 reg2051,
                 forvar2050,
                 reg2049,
                 forvar2048,
                 reg2047,
                 forvar2046,
                 reg2045,
                 reg2044,
                 reg2043,
                 wire2042,
                 reg2041,
                 reg2040,
                 forvar2039,
                 reg2038,
                 reg2037,
                 reg2036,
                 reg2035,
                 reg2034,
                 reg2033,
                 reg2032,
                 reg2031,
                 reg2030,
                 forvar2029,
                 reg2028,
                 reg2027,
                 reg2026,
                 reg2025,
                 reg2024,
                 forvar2023,
                 reg2022,
                 forvar2021,
                 reg2020,
                 reg2019,
                 reg2018,
                 forvar2017,
                 reg2016,
                 reg2015,
                 reg2014,
                 forvar2013,
                 wire2012,
                 reg2011,
                 reg2010,
                 wire2009,
                 reg2008,
                 reg2007,
                 reg2006,
                 reg2005,
                 wire2004,
                 reg2003,
                 reg2002,
                 reg2001,
                 reg2000,
                 reg1999,
                 reg1998,
                 reg1993,
                 forvar1988,
                 reg1997,
                 reg1996,
                 reg1995,
                 reg1994,
                 forvar1993,
                 reg1992,
                 forvar1991,
                 reg1990,
                 reg1989,
                 reg1988,
                 reg1987,
                 reg1986,
                 reg1985,
                 reg1984,
                 reg1983,
                 reg1982,
                 reg1981,
                 reg1980,
                 reg1979,
                 forvar1978,
                 forvar1977,
                 reg1976,
                 reg1975,
                 reg1974,
                 reg1973,
                 reg1972,
                 reg1971,
                 reg1970,
                 reg1969,
                 reg1968,
                 reg1967,
                 forvar1966,
                 reg1965,
                 forvar1964,
                 reg1963,
                 reg1962,
                 reg1961,
                 reg1960,
                 reg1959,
                 forvar1958,
                 forvar1957,
                 reg1956,
                 forvar1955,
                 reg1954,
                 reg1953,
                 forvar1952,
                 forvar1951,
                 reg1950,
                 reg1949,
                 reg1948,
                 reg1947,
                 reg1946,
                 reg1945,
                 reg1944,
                 reg1943,
                 reg1942,
                 forvar1941,
                 reg1940,
                 reg1939,
                 forvar1938,
                 forvar1937,
                 reg1936,
                 reg1935,
                 reg1934,
                 reg1933,
                 reg1932,
                 reg1931,
                 reg1930,
                 reg1929,
                 reg1928,
                 forvar1927,
                 reg1927,
                 reg1926,
                 reg1925,
                 reg1924,
                 reg1923,
                 reg1922,
                 reg1921,
                 reg1920,
                 forvar1919,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar1919 = (1'h0); (forvar1919 < (1'h1)); forvar1919 = (forvar1919 + (1'h1)))
        begin
          reg1920 <= (|$unsigned($unsigned("Q")));
          reg1921 <= ("B6M7wVknAnT3pvYqUQB" ?
              ((wire1918[(2'h3):(2'h2)] ?
                  (wire1916[(1'h0):(1'h0)] ?
                      (-wire1916) : $unsigned(reg1920)) : wire1918[(1'h1):(1'h1)]) && ({(!(8'hbe)),
                      (8'ha6)} ?
                  "xc8gMp" : {wire1918, "f1M"})) : (~&{"M8eGYsmBE1"}));
          reg1922 <= $unsigned((("" ?
              {(reg1921 * wire1917),
                  (reg1921 ? wire1915 : (8'hae))} : ($unsigned(reg1920) ?
                  (wire1918 != reg1921) : $unsigned(wire1917))) >> "BCfIoq6"));
        end
      if (((wire1917 ?
              $unsigned($signed((!reg1922))) : (reg1920[(3'h4):(1'h1)] & {wire1918[(5'h10):(3'h4)],
                  $signed(wire1915)})) ?
          {"ciY7bVrh"} : (|"O74cTYGLm")))
        begin
          reg1923 <= wire1918[(4'hc):(3'h4)];
          reg1924 = wire1916[(3'h7):(2'h3)];
          reg1925 <= $unsigned($signed(wire1916));
          reg1926 = $signed(({"Omb7bmm4eo", wire1917} ?
              $unsigned({reg1920[(3'h4):(1'h1)],
                  $unsigned((8'ha6))}) : reg1925));
          reg1927 <= "OrYoHsdUm3c8kyC44f3Q8h";
        end
      else
        begin
          reg1923 <= ((wire1918 ?
              (!$signed((8'ha3))) : $unsigned($signed((reg1923 ?
                  reg1927 : wire1918)))) >= forvar1919);
          reg1924 <= $unsigned($unsigned(($unsigned(reg1924) ?
              (reg1924[(4'hb):(3'h7)] ?
                  "fFbbLy09ywV82XzUC0gfJHQ" : (reg1922 < reg1927)) : $signed((wire1917 & wire1916)))));
          reg1925 <= {reg1927[(1'h1):(1'h1)],
              {((&forvar1919[(4'h8):(4'h8)]) - "u"),
                  (~^$unsigned(forvar1919[(2'h3):(1'h1)]))}};
          if (reg1924)
            begin
              reg1926 <= ($signed(($signed($signed(reg1924)) ?
                  "JMM7M9dGh8qIsLHT65t4y" : $signed((|(7'h43))))) ~^ (^~{reg1927[(4'hc):(1'h1)]}));
              for (forvar1927 = (1'h0); (forvar1927 < (1'h1)); forvar1927 = (forvar1927 + (1'h1)))
                begin
                  reg1928 <= reg1921[(3'h5):(3'h4)];
                  reg1929 = (+$unsigned({wire1916, "kOAsJr9UsqnygH2dzPZH6QX"}));
                  reg1930 = "Dshk9XR3";
                  reg1931 = (!forvar1919);
                  reg1932 <= (($unsigned((wire1915[(4'h9):(4'h9)] >= (reg1923 ?
                          reg1920 : forvar1927))) == $signed($signed(reg1922))) ?
                      $unsigned($unsigned(($signed(reg1921) & "P0EmtymOvH"))) : forvar1927[(3'h6):(1'h0)]);
                end
              reg1933 = $signed(reg1924[(3'h4):(2'h3)]);
              reg1934 = "KcUfFAV";
              reg1935 <= $unsigned((((!$signed(forvar1927)) ?
                      $signed(reg1922) : reg1933) ?
                  ((!reg1925) <= (((8'h9e) >= (7'h45)) ^~ (~|reg1934))) : ((8'ha4) ^~ "ZU1YKoXl56")));
            end
          else
            begin
              reg1926 <= wire1915[(4'hb):(3'h6)];
              for (forvar1927 = (1'h0); (forvar1927 < (3'h4)); forvar1927 = (forvar1927 + (1'h1)))
                begin
                  reg1928 <= reg1928[(4'h8):(4'h8)];
                  reg1929 <= (($unsigned($signed("au")) ?
                      ($signed((reg1930 <= reg1934)) ?
                          (+((8'hb1) ?
                              (8'h9e) : reg1920)) : $signed((8'h9f))) : "nb1T6fDmpUHq") >>> "L9XOL06L");
                  reg1930 <= (|($unsigned($signed($signed(forvar1927))) <= ((|(reg1926 ?
                          reg1928 : wire1916)) ?
                      "ShVK3EOTXZkJt0U2I" : {(8'ha7)})));
                  reg1931 <= (reg1920 - $unsigned(reg1933));
                  reg1932 <= (((-reg1922) ?
                          wire1916[(2'h2):(1'h0)] : reg1932[(2'h3):(1'h1)]) ?
                      $unsigned($signed($signed($signed(reg1933)))) : "tkJ6YM6MKCm2s");
                end
              reg1933 <= (reg1928[(4'hb):(4'hb)] ?
                  (reg1921 || reg1922) : reg1926);
              reg1934 = ($signed((8'had)) ?
                  reg1934 : (({$unsigned(reg1930),
                      reg1921[(5'h16):(5'h16)]} - reg1924[(2'h2):(2'h2)]) ~^ wire1915[(4'h8):(3'h7)]));
              reg1935 <= forvar1919[(4'ha):(4'ha)];
              reg1936 <= {"SHfPs8lZzEsCrkD6qbMOF"};
            end
          for (forvar1937 = (1'h0); (forvar1937 < (3'h5)); forvar1937 = (forvar1937 + (1'h1)))
            begin
              for (forvar1938 = (1'h0); (forvar1938 < (2'h2)); forvar1938 = (forvar1938 + (1'h1)))
                begin
                  reg1939 <= reg1929[(2'h3):(1'h0)];
                end
              reg1940 <= $unsigned($unsigned((~{(reg1939 ?
                      (8'hb3) : reg1932)})));
              for (forvar1941 = (1'h0); (forvar1941 < (2'h3)); forvar1941 = (forvar1941 + (1'h1)))
                begin
                  reg1942 = (reg1935[(3'h5):(2'h2)] ?
                      reg1931[(3'h6):(3'h6)] : (($unsigned((wire1916 ?
                              wire1918 : reg1920)) <= ((^~reg1936) ^~ (reg1936 << (7'h4b)))) ?
                          (reg1920[(3'h6):(3'h4)] ?
                              ($signed((8'hbc)) - {reg1926}) : ((~^wire1916) ?
                                  (~^reg1926) : $unsigned(wire1918))) : ("PaxzIO7IBeSB" ?
                              (((8'hb2) ?
                                  forvar1937 : (8'ha9)) <<< "49GBstT07oDY9ynEYb8bX5zZ") : $signed((|reg1929)))));
                  reg1943 <= "9yGma1aD2X8790uH";
                end
              reg1944 <= $signed({{"aLPVWcmD73SoaP8h11WJd"}});
              if (("Nh9VL6VXbuUFhoaAX" ? $signed(reg1926) : "DAF7w8qSyt"))
                begin
                  reg1945 = (8'haa);
                  reg1946 <= $signed((-(reg1933[(4'hb):(4'h9)] ?
                      {(~^reg1940)} : (7'h47))));
                  reg1947 <= $signed(reg1943[(1'h0):(1'h0)]);
                  reg1948 <= (-{(~&((reg1940 ? reg1920 : reg1924) ?
                          $unsigned((7'h4b)) : $signed(reg1921))),
                      $unsigned((reg1926 == forvar1919[(3'h5):(3'h4)]))});
                  reg1949 <= reg1939[(3'h4):(1'h0)];
                  reg1950 <= ("fzcHoJG83T" ?
                      (($signed(forvar1941) ?
                          (-(reg1928 << reg1946)) : ($signed(reg1920) ?
                              "UsegKKP7Nnkpe9" : ((8'hb9) & reg1942))) | reg1944) : reg1939);
                end
              else
                begin
                  reg1945 <= (reg1943[(2'h2):(1'h1)] + reg1925);
                  reg1946 = "oJH3tTkQSiBpBVValNYfbDXd";
                  reg1947 <= ($signed("sNqNHidc30fZ5W9z") ?
                      (^reg1929[(1'h1):(1'h1)]) : reg1944);
                  reg1948 <= {"VQEeULhc6STCi6manM2g1JdXk"};
                  reg1949 <= reg1923[(4'h8):(4'h8)];
                end
            end
          for (forvar1951 = (1'h0); (forvar1951 < (2'h3)); forvar1951 = (forvar1951 + (1'h1)))
            begin
              for (forvar1952 = (1'h0); (forvar1952 < (3'h4)); forvar1952 = (forvar1952 + (1'h1)))
                begin
                  reg1953 <= (~(^$signed("827")));
                end
              reg1954 <= (("QkvM00t006mpba0HA74Y" ?
                  {$unsigned({reg1942,
                          reg1922})} : (~reg1934)) <= $signed(reg1934));
            end
        end
      for (forvar1955 = (1'h0); (forvar1955 < (1'h0)); forvar1955 = (forvar1955 + (1'h1)))
        begin
          reg1956 <= reg1943[(1'h1):(1'h1)];
          for (forvar1957 = (1'h0); (forvar1957 < (1'h0)); forvar1957 = (forvar1957 + (1'h1)))
            begin
              for (forvar1958 = (1'h0); (forvar1958 < (1'h0)); forvar1958 = (forvar1958 + (1'h1)))
                begin
                  reg1959 <= ((($unsigned($unsigned((8'ha8))) && "FtPLr6AUUZ") ?
                          {reg1944[(4'h9):(3'h7)]} : (&$unsigned($signed(reg1934)))) ?
                      ((~&(+(reg1926 ? reg1930 : (8'hbb)))) ?
                          reg1944 : "SllZdAgzq51zUQEatvmI") : "U");
                end
              reg1960 <= {"2fsayrYpRD"};
              reg1961 <= (((^forvar1955[(2'h3):(1'h0)]) ?
                  (7'h4c) : "ZeRp3CgFZvts3NC54HY") >= (~"nWMMBmtA9xQQBrv2Pd9HNW"));
              reg1962 <= reg1921;
            end
          reg1963 = (reg1953[(3'h4):(1'h0)] >= (^~reg1950));
          for (forvar1964 = (1'h0); (forvar1964 < (1'h0)); forvar1964 = (forvar1964 + (1'h1)))
            begin
              reg1965 = (!(|reg1930));
              for (forvar1966 = (1'h0); (forvar1966 < (3'h4)); forvar1966 = (forvar1966 + (1'h1)))
                begin
                  reg1967 <= ((^({$signed(forvar1955)} ~^ ((reg1936 ?
                              reg1926 : wire1918) ?
                          $signed(wire1918) : $signed(reg1927)))) ?
                      (reg1935 == (("AKtPqhV" || (8'ha4)) * $unsigned($signed(reg1925)))) : "nlw70EReISsOqC21hT6");
                  reg1968 <= (($signed($unsigned((&wire1917))) ?
                          reg1962 : (forvar1951[(3'h4):(1'h1)] ?
                              $unsigned((forvar1919 ?
                                  forvar1964 : (7'h42))) : ((~reg1930) == reg1936))) ?
                      $unsigned(reg1962[(3'h5):(3'h5)]) : (7'h40));
                  reg1969 = (^reg1967[(3'h5):(1'h1)]);
                  reg1970 = $signed({{({reg1948,
                              reg1924} >= (reg1922 & (8'ha3)))}});
                  reg1971 <= $unsigned(($unsigned((reg1929 ?
                      (~^reg1949) : {wire1918})) >> $signed($unsigned("0XpngNBrgpTg"))));
                  reg1972 <= {({"zhhm0fXtNrFCR", reg1942[(2'h2):(1'h0)]} ?
                          ("FmzOy2q2UCPQ5Xah" ?
                              ((7'h48) ?
                                  wire1916 : {reg1947}) : $signed($unsigned((8'hb7)))) : (forvar1937[(2'h3):(2'h2)] | (~reg1960[(4'hd):(1'h1)])))};
                end
              reg1973 = $signed(("GA" ? "Fh7xv6qcF3lcE7" : reg1961));
              reg1974 = ((reg1953[(1'h0):(1'h0)] ?
                      {{(~^reg1931)}} : ("Lyuh70Ms20SIMnosXE" ^~ reg1940)) ?
                  (($unsigned($signed(reg1949)) ?
                      (~&{reg1970}) : {(reg1973 ? (8'haf) : (8'h9d)),
                          $signed(reg1965)}) < wire1917) : (("2YedmiGDaYphHgAK93AT" >> (^~reg1950[(1'h0):(1'h0)])) > {reg1948[(2'h3):(1'h1)]}));
              reg1975 <= "lPzuii";
              reg1976 <= (|wire1915[(4'h9):(2'h3)]);
            end
          for (forvar1977 = (1'h0); (forvar1977 < (2'h3)); forvar1977 = (forvar1977 + (1'h1)))
            begin
              for (forvar1978 = (1'h0); (forvar1978 < (3'h4)); forvar1978 = (forvar1978 + (1'h1)))
                begin
                  reg1979 = $unsigned("92IdYP");
                  reg1980 <= ($unsigned($unsigned($signed((reg1954 << reg1922)))) ?
                      ((~{$unsigned((8'ha2))}) >> (((+(8'hb0)) ?
                          "y" : $signed((8'ha8))) >>> $unsigned((reg1950 | reg1960)))) : "iaIDkb7xkiaRzcJlbJA");
                  reg1981 <= $unsigned(($signed(((&reg1962) ?
                      reg1970 : "NWt")) || reg1974[(4'hc):(2'h2)]));
                  reg1982 <= (^~"Q");
                  reg1983 <= forvar1938[(2'h2):(1'h1)];
                end
              reg1984 <= (&((~^reg1947) < $unsigned($signed($unsigned(reg1976)))));
            end
          reg1985 <= (~reg1926);
        end
      reg1986 <= (reg1928 ?
          (^~(~^(8'ha1))) : (~^$signed("rbGAM5xii4JLl9QPFMkA3IJUP")));
      if (forvar1966[(1'h0):(1'h0)])
        begin
          reg1987 = (+(~|$signed(($unsigned(reg1981) > ((8'had) ?
              reg1920 : reg1947)))));
          reg1988 = (("" ~^ $signed({reg1922})) ~^ (^~(|$unsigned("LK"))));
          reg1989 <= reg1931[(3'h5):(1'h1)];
          reg1990 = $signed($unsigned(reg1987));
          for (forvar1991 = (1'h0); (forvar1991 < (1'h0)); forvar1991 = (forvar1991 + (1'h1)))
            begin
              reg1992 <= reg1933;
              for (forvar1993 = (1'h0); (forvar1993 < (2'h3)); forvar1993 = (forvar1993 + (1'h1)))
                begin
                  reg1994 = "3B4ZXcqzPJT";
                  reg1995 <= "EG9kdXPyJkq5cMTxHc";
                end
              reg1996 <= $unsigned((^~(((reg1972 > reg1959) ^ $unsigned(reg1933)) << "h")));
              reg1997 <= reg1939;
            end
        end
      else
        begin
          reg1987 <= $unsigned(("mVPHThcS1wiluYBsLcc4Nl3MX" ?
              (+(((8'hbf) >> reg1965) ?
                  $unsigned(forvar1958) : reg1990[(1'h1):(1'h0)])) : (~&(reg1962 < ((7'h48) ?
                  reg1983 : (8'ha2))))));
          for (forvar1988 = (1'h0); (forvar1988 < (3'h4)); forvar1988 = (forvar1988 + (1'h1)))
            begin
              reg1989 = $signed("inLBErMANBzMmeDJiYTiKsM");
              reg1990 = (^~(reg1924[(3'h5):(1'h1)] << forvar1951));
              for (forvar1991 = (1'h0); (forvar1991 < (2'h3)); forvar1991 = (forvar1991 + (1'h1)))
                begin
                  reg1992 <= reg1956[(2'h3):(2'h2)];
                end
              reg1993 <= ("0WXGMV" ?
                  ((reg1929[(2'h2):(1'h0)] ? forvar1919 : forvar1964) ?
                      $signed("tfDhCNpDaRaRWl1d") : (~^"")) : ((~^(+(^reg1984))) ?
                      ((~{forvar1977}) + forvar1993) : "zEI"));
              reg1994 <= $unsigned(("2pyy70dHdT9T0Jiuu7N5HTWp" == reg1971[(1'h1):(1'h1)]));
              reg1995 = ((((~|(forvar1952 ?
                  reg1980 : reg1922)) <<< "WmSBtcqH5s9ImIblJHtzd") - $unsigned(forvar1978)) <= reg1933);
            end
          reg1996 <= (((~(-$signed(reg1970))) ?
                  "QcHwQysQwhuXcrFQRZnho" : (+($unsigned(forvar1938) & $signed(reg1976)))) ?
              ("dv" ?
                  $unsigned(reg1954[(4'h9):(4'h9)]) : (-($unsigned(reg1979) ?
                      reg1996[(4'hc):(4'h9)] : $unsigned(reg1944)))) : ("lNrGb0gkCPSWi5OqPZ" ?
                  "SB9zNY" : (((~^reg1934) == (reg1939 || (7'h42))) ?
                      forvar1938[(1'h0):(1'h0)] : (^~(-reg1963)))));
          reg1997 <= $unsigned("YNz5NJxssk0TnaN8honG");
          reg1998 <= ({reg1930[(5'h14):(4'ha)]} - $signed(forvar1938[(2'h2):(1'h1)]));
        end
    end
  always
    @(posedge clk) begin
      reg1999 <= $signed(reg1962[(3'h7):(3'h4)]);
      reg2000 = reg1953;
      reg2001 <= {(|(($signed(forvar1977) >>> "NcPcnquPQep8nABU0Ju6O6") & (^((8'hbb) ?
              forvar1955 : (8'h9d))))),
          ((("7vZdIxzweq4t" ?
                      reg1949[(4'he):(1'h1)] : (reg1986 <= forvar1955)) ?
                  ("w" == $signed(reg1944)) : reg1993[(1'h0):(1'h0)]) ?
              "BJUvrHlFdC4smwldRFV" : (reg1980 | reg1980[(3'h6):(3'h5)]))};
    end
  always
    @(posedge clk) begin
      reg2002 <= $signed($unsigned(((reg1927 & (+(8'hbf))) & "4agKSkuoXhH2QYDn4hPze")));
      reg2003 <= $signed((-reg1996));
    end
  assign wire2004 = reg1950[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      reg2005 = $unsigned((reg1954 * (~&$unsigned("aOS7w1EW"))));
      reg2006 <= reg1994;
      reg2007 <= wire1917[(1'h0):(1'h0)];
      reg2008 <= reg1956;
    end
  assign wire2009 = reg1963[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg2010 = $unsigned($signed(reg1973[(4'hf):(2'h3)]));
      reg2011 <= $unsigned("LZIJhHlJ6kEGqPSOWRe9Qznx");
    end
  assign wire2012 = "Fb5gX";
  always
    @(posedge clk) begin
      for (forvar2013 = (1'h0); (forvar2013 < (1'h0)); forvar2013 = (forvar2013 + (1'h1)))
        begin
          reg2014 <= (($unsigned($unsigned((reg1997 ?
                  forvar1952 : wire1917))) | reg1997) ?
              forvar1941 : reg1983[(2'h2):(1'h1)]);
          reg2015 = "m409pcA9uXGaTWH5oeHK4A";
          reg2016 = "eWa9cCkCltl3YTfT18";
        end
      for (forvar2017 = (1'h0); (forvar2017 < (3'h5)); forvar2017 = (forvar2017 + (1'h1)))
        begin
          reg2018 <= $unsigned((~^{reg1988[(2'h2):(1'h1)], ""}));
          reg2019 <= "PDFPbKemBQg";
          reg2020 <= (reg1990 ?
              ({reg1992} << (8'haf)) : ((((wire2004 ^~ reg2015) >= (reg1931 & (8'hbb))) ?
                      ($unsigned(reg1981) ?
                          $unsigned(reg2015) : (reg1998 ?
                              reg2003 : forvar1991)) : $unsigned($signed(forvar1958))) ?
                  forvar1955[(2'h2):(1'h0)] : (~|reg1931)));
          for (forvar2021 = (1'h0); (forvar2021 < (3'h5)); forvar2021 = (forvar2021 + (1'h1)))
            begin
              reg2022 <= forvar2017[(4'h8):(2'h2)];
              for (forvar2023 = (1'h0); (forvar2023 < (1'h1)); forvar2023 = (forvar2023 + (1'h1)))
                begin
                  reg2024 = reg1981;
                  reg2025 = (~(~^$unsigned($signed((forvar1978 ?
                      reg2001 : wire1916)))));
                  reg2026 <= reg2024;
                  reg2027 = {($signed($signed($signed(reg1942))) || {(-(reg2001 ?
                              reg1998 : reg1970)),
                          reg1979[(4'ha):(4'h9)]}),
                      $signed(reg1983[(3'h4):(2'h3)])};
                  reg2028 <= $unsigned("f4FYrQE63VpYZyyC0XXtpuI");
                end
            end
          for (forvar2029 = (1'h0); (forvar2029 < (1'h1)); forvar2029 = (forvar2029 + (1'h1)))
            begin
              reg2030 <= reg1982;
              reg2031 = (~^$signed(($signed((reg1973 ? reg1935 : (8'h9e))) ?
                  (~|(^(7'h46))) : "D4N3I9t3GZmNNY0gvdgvpJ")));
              reg2032 <= $signed(forvar1937[(1'h0):(1'h0)]);
            end
        end
      reg2033 <= {$signed(reg1986)};
    end
  always
    @(posedge clk) begin
      reg2034 <= (~($signed((~$unsigned(reg1979))) ? "DXbLbcTi" : reg1947));
      reg2035 <= "aiJrnoFINeGi";
      reg2036 <= $unsigned(reg2033);
      reg2037 = reg1944;
      reg2038 <= forvar1978;
      for (forvar2039 = (1'h0); (forvar2039 < (3'h5)); forvar2039 = (forvar2039 + (1'h1)))
        begin
          reg2040 <= $unsigned((8'hb2));
          reg2041 <= reg2025;
        end
    end
  assign wire2042 = (-$signed(((reg1947[(4'h8):(1'h1)] >= "96NduM") ?
                        $signed("YaTrX2DeD5lcHod") : $signed((forvar1958 ?
                            reg1922 : reg1925)))));
  always
    @(posedge clk) begin
      reg2043 <= (((&forvar1919[(4'h9):(1'h0)]) ~^ $unsigned($unsigned((reg2014 ?
          reg1927 : reg2028)))) >> "FEr6bEeBJT6KJcW6gX");
      reg2044 = $unsigned(((~(((8'hab) ? reg2020 : wire1918) != reg2018)) ?
          $signed($signed((reg1954 ?
              (8'hb5) : reg1926))) : ("i9p3X" * wire1917)));
      reg2045 <= "FWe3hQfDRY82Qsh9";
      for (forvar2046 = (1'h0); (forvar2046 < (3'h5)); forvar2046 = (forvar2046 + (1'h1)))
        begin
          reg2047 <= "4yRPa9WPOo8";
          for (forvar2048 = (1'h0); (forvar2048 < (3'h5)); forvar2048 = (forvar2048 + (1'h1)))
            begin
              reg2049 <= $unsigned(wire1915[(3'h4):(2'h2)]);
              for (forvar2050 = (1'h0); (forvar2050 < (3'h4)); forvar2050 = (forvar2050 + (1'h1)))
                begin
                  reg2051 = $signed(((("TW3xt8q6mwO0evbWF" <= reg2015[(1'h1):(1'h1)]) - (!$unsigned(reg1926))) < $unsigned(reg2041)));
                  reg2052 <= $unsigned("qIQSHhIB1");
                  reg2053 <= "EwTcTLMUlrTgComq7";
                  reg2054 <= (^(reg1981 ?
                      reg1944[(3'h7):(1'h0)] : (reg1996 & (^~(reg2027 ?
                          forvar1957 : forvar1941)))));
                  reg2055 <= $signed({{((reg1927 ?
                              wire1918 : reg2027) & "yE4Tg8bKWC2WwE")},
                      ((^~(~^reg1935)) <<< (reg2024[(2'h3):(2'h3)] ?
                          (8'hab) : {forvar1964, reg2027}))});
                  reg2056 <= "5kHHumP";
                end
              for (forvar2057 = (1'h0); (forvar2057 < (3'h4)); forvar2057 = (forvar2057 + (1'h1)))
                begin
                  reg2058 <= reg2015[(3'h5):(2'h3)];
                  reg2059 <= ($signed($signed(forvar1951[(1'h1):(1'h0)])) ?
                      ($unsigned(((8'ha8) + reg2001[(5'h18):(5'h16)])) * $unsigned(reg1984[(2'h3):(1'h0)])) : "LGzYQgVHIcy");
                  reg2060 <= reg2026[(2'h3):(1'h0)];
                  reg2061 <= (!(&(~^({reg2010, forvar1988} ?
                      ((7'h48) <<< forvar1937) : $signed(reg2015)))));
                  reg2062 <= $unsigned({({forvar1952} ?
                          (7'h4d) : {(reg1936 || reg1976), reg2041})});
                end
              reg2063 <= $signed(reg1974[(1'h1):(1'h0)]);
              reg2064 <= "VsvRUqUlWNeXaEpe9B";
            end
          reg2065 <= reg2034[(5'h11):(4'ha)];
          reg2066 <= ($signed(reg2055) ?
              forvar2023[(1'h1):(1'h0)] : (({(~reg1925),
                  "OD2Hbz3BUX2pv3RuGo"} >= (^~reg2038)) - ({(reg1982 && (8'hb6))} | (~|(8'hb0)))));
          reg2067 <= $signed($signed($signed({$unsigned(reg1987)})));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1872
#( parameter param1911 = (^((~|(~(&(7'h4a)))) << (~((-(8'hbf)) >>> ((8'hb7) != (7'h47)))))) )
(y, clk, wire1877, wire1876, wire1875, wire1874, wire1873);
  output wire [(32'h1c4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire1877;
  input wire signed [(3'h5):(1'h0)] wire1876;
  input wire signed [(2'h3):(1'h0)] wire1875;
  input wire [(5'h17):(1'h0)] wire1874;
  input wire signed [(5'h16):(1'h0)] wire1873;
  reg [(4'hb):(1'h0)] reg1910 = (1'h0);
  reg [(4'h9):(1'h0)] reg1909 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1908;
  reg [(5'h11):(1'h0)] reg1907 = (1'h0);
  reg [(5'h19):(1'h0)] reg1906 = (1'h0);
  reg [(3'h7):(1'h0)] reg1905 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1904 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1903 = (1'h0);
  reg [(2'h2):(1'h0)] reg1902 = (1'h0);
  reg [(4'ha):(1'h0)] reg1901 = (1'h0);
  reg [(5'h12):(1'h0)] reg1900 = (1'h0);
  reg [(4'h9):(1'h0)] reg1899 = (1'h0);
  reg [(5'h10):(1'h0)] reg1898 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1897 = (1'h0);
  reg [(4'ha):(1'h0)] reg1896 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1895 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1894 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1893 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1892 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1891 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1890 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1889 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1888 = (1'h0);
  reg [(3'h4):(1'h0)] reg1887 = (1'h0);
  reg [(5'h15):(1'h0)] reg1886 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1885 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire1884;
  reg signed [(2'h3):(1'h0)] reg1883 = (1'h0);
  reg [(2'h3):(1'h0)] reg1882 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1881 = (1'h0);
  reg [(3'h6):(1'h0)] reg1880 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1879 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1878 = (1'h0);
  assign y = {reg1910,
                 reg1909,
                 wire1908,
                 reg1907,
                 reg1906,
                 reg1905,
                 reg1904,
                 forvar1903,
                 reg1902,
                 reg1901,
                 reg1900,
                 reg1899,
                 reg1898,
                 reg1897,
                 reg1896,
                 reg1895,
                 forvar1894,
                 reg1893,
                 forvar1892,
                 reg1891,
                 reg1890,
                 forvar1889,
                 reg1888,
                 reg1887,
                 reg1886,
                 reg1885,
                 wire1884,
                 reg1883,
                 reg1882,
                 reg1881,
                 reg1880,
                 reg1879,
                 forvar1878,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar1878 = (1'h0); (forvar1878 < (1'h1)); forvar1878 = (forvar1878 + (1'h1)))
        begin
          reg1879 <= (^("aEAwUAYDpm4vq0m8AmQAhe4" >>> (^((wire1876 ?
                  wire1876 : wire1876) ?
              {(7'h4a)} : wire1876))));
          reg1880 = $unsigned(reg1879);
          reg1881 <= {($unsigned("rYYJwUHF23J") ^ "yK23gUWgAigdyouJg5Ay6bUm")};
        end
      reg1882 <= "WhmD9vIOp5pPFJC";
      reg1883 = reg1880;
    end
  assign wire1884 = "Nxp7VZHoQvfCAV5KMFb7";
  always
    @(posedge clk) begin
      reg1885 = {($signed(wire1875) ?
              {(!{(7'h45), (7'h44)}), forvar1878} : wire1875),
          $signed(("VLNC4MUec9e5W1WescABnsUS" ?
              (~^$signed(wire1884)) : "afs5m"))};
      reg1886 <= ($signed(($signed((+wire1876)) ?
              wire1876 : reg1882[(2'h3):(1'h0)])) ?
          $unsigned(wire1876) : reg1879[(3'h5):(2'h3)]);
      reg1887 <= reg1879[(3'h5):(3'h4)];
    end
  always
    @(posedge clk) begin
      reg1888 = {$unsigned({$unsigned("EB64lb51IESvv4VMNB8HDpF"),
              (-forvar1878)})};
      for (forvar1889 = (1'h0); (forvar1889 < (3'h5)); forvar1889 = (forvar1889 + (1'h1)))
        begin
          reg1890 <= $signed("9TDfsF9");
          reg1891 <= reg1880[(2'h3):(2'h2)];
          for (forvar1892 = (1'h0); (forvar1892 < (2'h2)); forvar1892 = (forvar1892 + (1'h1)))
            begin
              reg1893 <= (+(|(8'ha0)));
              for (forvar1894 = (1'h0); (forvar1894 < (1'h0)); forvar1894 = (forvar1894 + (1'h1)))
                begin
                  reg1895 <= $signed($signed(wire1875));
                  reg1896 <= "dJiQgiXcPie6lZ9mt";
                  reg1897 <= (((((~|reg1891) * (~&reg1890)) ?
                      (-forvar1889[(3'h7):(1'h1)]) : (-reg1887[(2'h3):(1'h0)])) || forvar1894) < (^~reg1887));
                end
              reg1898 <= wire1876[(1'h0):(1'h0)];
            end
        end
      reg1899 <= {((&(!(wire1876 ?
              (8'hac) : reg1883))) >>> reg1883[(2'h3):(1'h0)]),
          (!reg1885[(5'h18):(3'h7)])};
      reg1900 <= (7'h44);
      reg1901 <= $signed(reg1883);
      reg1902 <= (^~{(($unsigned(reg1899) >>> "tXKQRPh2aRRPiXQITLD1") ?
              "WbdmkdViYebGzUP6RidHqSWPk" : ($signed(reg1880) ?
                  (|reg1880) : forvar1878)),
          ((|reg1896) - ((|reg1883) ? reg1898 : $signed(reg1885)))});
    end
  always
    @(posedge clk) begin
      for (forvar1903 = (1'h0); (forvar1903 < (1'h0)); forvar1903 = (forvar1903 + (1'h1)))
        begin
          reg1904 <= (("lKTzRqLYEeK1CLcWt" ^~ (8'hb9)) ?
              (((7'h4d) > reg1896) <= (~^((7'h46) | forvar1903[(5'h10):(4'hd)]))) : reg1896[(1'h0):(1'h0)]);
        end
      reg1905 <= (~|$signed(((((8'hb8) ?
              forvar1892 : (8'hbe)) >= "GTxhyB49grno7IHLJLYYlXM") ?
          $signed($unsigned(reg1880)) : "BCM")));
      reg1906 <= reg1899;
      reg1907 = reg1895;
    end
  assign wire1908 = (!(((wire1877 ? reg1881 : reg1905[(3'h5):(1'h1)]) ?
                            reg1898 : "Rdtg2gXUs") ?
                        $signed(reg1905) : $signed(($unsigned((8'hb9)) ?
                            "ef" : ((7'h43) << forvar1894)))));
  always
    @(posedge clk) begin
      reg1909 <= (~|((wire1874[(1'h0):(1'h0)] ~^ (reg1897[(4'hd):(3'h4)] & $unsigned(wire1875))) ?
          (((reg1898 >> forvar1894) <<< $signed(reg1895)) ?
              reg1887[(2'h2):(2'h2)] : "SydZrRemVJo0BR") : (reg1880[(3'h4):(3'h4)] >>> ((~wire1876) ?
              $unsigned((8'had)) : (~^reg1898)))));
      reg1910 <= reg1887[(2'h3):(2'h3)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1674
#( parameter param1833 = (({(|((8'ha1) < (8'ha5))), ({(8'ha0), (8'hbc)} ? {(8'had), (7'h43)} : (+(8'ha5)))} ? (({(7'h4b)} ? (~&(7'h4a)) : ((8'hba) ? (8'hb3) : (8'haf))) ^~ ((~|(7'h4d)) ^ (~&(7'h46)))) : (((~&(7'h41)) ? ((7'h43) <<< (8'ha7)) : (~|(8'h9f))) != (((8'hb9) >> (7'h4a)) ? (~|(8'haa)) : ((7'h46) ? (7'h47) : (7'h47))))) ? (8'hac) : ((+(((7'h4c) != (8'h9c)) != ((7'h42) ? (8'hb5) : (7'h48)))) ? (^(((8'h9f) >> (8'hb4)) < {(7'h44), (7'h45)})) : {(-((8'hbc) ? (7'h4e) : (7'h47))), (((7'h4e) > (8'hae)) << ((8'ha4) ? (8'hb4) : (7'h45)))}))
, parameter param1834 = (((((param1833 < param1833) ? ((8'hbf) * param1833) : param1833) ? (~^(param1833 >>> param1833)) : param1833) ? (+((param1833 ? param1833 : param1833) ~^ (~param1833))) : param1833) != (^~(-(!param1833)))) )
(y, clk, wire1679, wire1678, wire1677, wire1676, wire1675);
  output wire [(32'h8fe):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire1679;
  input wire signed [(5'h13):(1'h0)] wire1678;
  input wire [(5'h16):(1'h0)] wire1677;
  input wire signed [(2'h2):(1'h0)] wire1676;
  input wire [(5'h11):(1'h0)] wire1675;
  reg signed [(5'h14):(1'h0)] reg1832 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1831 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1830 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1829 = (1'h0);
  reg [(5'h11):(1'h0)] reg1828 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1827 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1826 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1825 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1824 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1823 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1822 = (1'h0);
  reg [(4'h8):(1'h0)] reg1821 = (1'h0);
  reg [(5'h18):(1'h0)] reg1820 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1819 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1818 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1817 = (1'h0);
  reg [(5'h11):(1'h0)] reg1816 = (1'h0);
  reg [(5'h11):(1'h0)] reg1815 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1814 = (1'h0);
  reg [(3'h7):(1'h0)] reg1813 = (1'h0);
  reg [(5'h19):(1'h0)] reg1812 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1811 = (1'h0);
  reg [(5'h12):(1'h0)] reg1810 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1809 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1808 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1807 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1806 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1805 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1804 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1803 = (1'h0);
  reg [(5'h12):(1'h0)] reg1802 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1801 = (1'h0);
  reg [(4'hc):(1'h0)] reg1800 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1799 = (1'h0);
  reg [(5'h15):(1'h0)] reg1798 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1797 = (1'h0);
  wire signed [(5'h16):(1'h0)] wire1796;
  reg signed [(5'h17):(1'h0)] reg1795 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1794 = (1'h0);
  reg [(5'h14):(1'h0)] reg1793 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1792 = (1'h0);
  reg [(4'hf):(1'h0)] reg1791 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1790 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1789 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1788 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1787 = (1'h0);
  reg [(4'ha):(1'h0)] reg1786 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1785 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1784 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1783 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1782 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1781 = (1'h0);
  reg [(5'h11):(1'h0)] reg1780 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1779 = (1'h0);
  reg [(5'h15):(1'h0)] reg1778 = (1'h0);
  reg [(5'h19):(1'h0)] reg1777 = (1'h0);
  reg [(2'h2):(1'h0)] reg1776 = (1'h0);
  reg [(5'h19):(1'h0)] reg1775 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1774 = (1'h0);
  reg [(4'h9):(1'h0)] reg1773 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1772 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1771 = (1'h0);
  reg [(4'hf):(1'h0)] reg1770 = (1'h0);
  wire [(3'h5):(1'h0)] wire1769;
  reg signed [(4'h9):(1'h0)] reg1768 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1767 = (1'h0);
  reg [(4'h9):(1'h0)] reg1766 = (1'h0);
  reg [(4'hb):(1'h0)] reg1765 = (1'h0);
  wire [(3'h4):(1'h0)] wire1764;
  reg signed [(5'h19):(1'h0)] reg1763 = (1'h0);
  reg [(4'ha):(1'h0)] reg1762 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1761 = (1'h0);
  reg [(5'h14):(1'h0)] reg1760 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1759 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1758 = (1'h0);
  reg [(5'h11):(1'h0)] reg1757 = (1'h0);
  reg [(2'h2):(1'h0)] reg1756 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1755 = (1'h0);
  wire [(5'h12):(1'h0)] wire1754;
  reg signed [(5'h19):(1'h0)] reg1753 = (1'h0);
  wire [(5'h15):(1'h0)] wire1752;
  reg signed [(5'h18):(1'h0)] reg1751 = (1'h0);
  reg [(3'h6):(1'h0)] reg1750 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1749 = (1'h0);
  reg [(5'h19):(1'h0)] reg1748 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1747 = (1'h0);
  reg [(5'h16):(1'h0)] reg1746 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1745 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1744 = (1'h0);
  reg [(4'hf):(1'h0)] reg1743 = (1'h0);
  reg [(5'h18):(1'h0)] reg1742 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1741 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1740 = (1'h0);
  reg [(4'hc):(1'h0)] reg1739 = (1'h0);
  reg [(4'hc):(1'h0)] reg1738 = (1'h0);
  reg [(4'h9):(1'h0)] reg1737 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1736 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1735 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1734 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1733 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1732 = (1'h0);
  reg [(5'h18):(1'h0)] reg1731 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1730 = (1'h0);
  reg [(5'h11):(1'h0)] reg1729 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1728 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1727 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1726 = (1'h0);
  reg [(3'h7):(1'h0)] reg1725 = (1'h0);
  reg [(5'h16):(1'h0)] reg1724 = (1'h0);
  reg [(2'h3):(1'h0)] reg1723 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1722 = (1'h0);
  reg [(5'h19):(1'h0)] reg1721 = (1'h0);
  reg [(2'h2):(1'h0)] reg1720 = (1'h0);
  reg [(4'hf):(1'h0)] reg1719 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1718 = (1'h0);
  wire [(4'hc):(1'h0)] wire1717;
  reg [(3'h7):(1'h0)] reg1716 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1715 = (1'h0);
  reg [(5'h13):(1'h0)] reg1714 = (1'h0);
  reg [(5'h14):(1'h0)] reg1713 = (1'h0);
  reg [(3'h6):(1'h0)] reg1712 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1711 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1710 = (1'h0);
  reg [(4'hd):(1'h0)] reg1709 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1708 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1707 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1706 = (1'h0);
  reg [(5'h15):(1'h0)] reg1705 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1704 = (1'h0);
  wire [(5'h17):(1'h0)] wire1703;
  reg [(4'h9):(1'h0)] reg1690 = (1'h0);
  reg [(2'h2):(1'h0)] reg1688 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1686 = (1'h0);
  reg [(5'h19):(1'h0)] reg1702 = (1'h0);
  reg [(5'h10):(1'h0)] reg1701 = (1'h0);
  reg [(5'h17):(1'h0)] reg1700 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1699 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1698 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1697 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1696 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1695 = (1'h0);
  reg [(4'ha):(1'h0)] reg1694 = (1'h0);
  reg [(3'h7):(1'h0)] reg1693 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1692 = (1'h0);
  reg [(2'h2):(1'h0)] reg1691 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1690 = (1'h0);
  reg [(4'h9):(1'h0)] reg1689 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1688 = (1'h0);
  reg [(3'h6):(1'h0)] reg1687 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1686 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1685 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1684 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1683 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1682 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1681 = (1'h0);
  wire [(4'ha):(1'h0)] wire1680;
  assign y = {reg1832,
                 reg1831,
                 reg1830,
                 reg1829,
                 reg1828,
                 forvar1827,
                 reg1826,
                 reg1825,
                 reg1824,
                 reg1823,
                 forvar1822,
                 reg1821,
                 reg1820,
                 reg1819,
                 reg1818,
                 reg1817,
                 reg1816,
                 reg1815,
                 reg1814,
                 reg1813,
                 reg1812,
                 reg1811,
                 reg1810,
                 forvar1809,
                 forvar1808,
                 reg1807,
                 reg1806,
                 reg1805,
                 forvar1804,
                 forvar1803,
                 reg1802,
                 reg1801,
                 reg1800,
                 reg1799,
                 reg1798,
                 forvar1797,
                 wire1796,
                 reg1795,
                 reg1794,
                 reg1793,
                 reg1792,
                 reg1791,
                 reg1790,
                 forvar1789,
                 forvar1788,
                 reg1787,
                 reg1786,
                 reg1785,
                 reg1784,
                 reg1783,
                 reg1782,
                 forvar1781,
                 reg1780,
                 forvar1779,
                 reg1778,
                 reg1777,
                 reg1776,
                 reg1775,
                 forvar1774,
                 reg1773,
                 reg1772,
                 forvar1771,
                 reg1770,
                 wire1769,
                 reg1768,
                 forvar1767,
                 reg1766,
                 reg1765,
                 wire1764,
                 reg1763,
                 reg1762,
                 reg1761,
                 reg1760,
                 reg1759,
                 reg1758,
                 reg1757,
                 reg1756,
                 forvar1755,
                 wire1754,
                 reg1753,
                 wire1752,
                 reg1751,
                 reg1750,
                 reg1749,
                 reg1748,
                 forvar1747,
                 reg1746,
                 reg1745,
                 forvar1744,
                 reg1743,
                 reg1742,
                 forvar1741,
                 reg1740,
                 reg1739,
                 reg1738,
                 reg1737,
                 forvar1736,
                 reg1735,
                 forvar1734,
                 reg1733,
                 reg1732,
                 reg1731,
                 reg1730,
                 reg1729,
                 reg1728,
                 reg1727,
                 forvar1726,
                 reg1725,
                 reg1724,
                 reg1723,
                 forvar1722,
                 reg1721,
                 reg1720,
                 reg1719,
                 forvar1718,
                 wire1717,
                 reg1716,
                 reg1715,
                 reg1714,
                 reg1713,
                 reg1712,
                 forvar1711,
                 reg1710,
                 reg1709,
                 reg1708,
                 forvar1707,
                 reg1706,
                 reg1705,
                 reg1704,
                 wire1703,
                 reg1690,
                 reg1688,
                 forvar1686,
                 reg1702,
                 reg1701,
                 reg1700,
                 reg1699,
                 forvar1698,
                 forvar1697,
                 reg1696,
                 reg1695,
                 reg1694,
                 reg1693,
                 reg1692,
                 reg1691,
                 forvar1690,
                 reg1689,
                 forvar1688,
                 reg1687,
                 reg1686,
                 reg1685,
                 reg1684,
                 forvar1683,
                 reg1682,
                 reg1681,
                 wire1680,
                 (1'h0)};
  assign wire1680 = $unsigned((wire1676 ? "NhD3Uphog1PGhNypXxUt" : wire1675));
  always
    @(posedge clk) begin
      reg1681 <= wire1678[(3'h7):(3'h7)];
      reg1682 <= $signed($signed($unsigned((~|$signed(reg1681)))));
      for (forvar1683 = (1'h0); (forvar1683 < (1'h1)); forvar1683 = (forvar1683 + (1'h1)))
        begin
          reg1684 = "oKIINN1LzDGWh94CvBAA0u19";
        end
      if (wire1675[(2'h2):(1'h0)])
        begin
          reg1685 <= (reg1682 <<< {(~^(8'ha6))});
          reg1686 <= wire1678[(4'hb):(3'h7)];
          reg1687 <= reg1684[(5'h12):(1'h0)];
          for (forvar1688 = (1'h0); (forvar1688 < (3'h4)); forvar1688 = (forvar1688 + (1'h1)))
            begin
              reg1689 = ((~&$signed($unsigned("UBUI4Wz"))) ?
                  $signed("c6qQKOSao8B") : "gHJ3qzhwlYLUCX5c58lP");
              for (forvar1690 = (1'h0); (forvar1690 < (3'h4)); forvar1690 = (forvar1690 + (1'h1)))
                begin
                  reg1691 <= reg1686[(2'h3):(1'h0)];
                  reg1692 <= ($unsigned((7'h44)) >= (~^wire1678));
                end
              reg1693 = {($signed($signed($signed(wire1680))) ?
                      ($signed($unsigned(wire1677)) ?
                          $unsigned((+reg1687)) : wire1679[(1'h0):(1'h0)]) : $signed((reg1681 != ((8'hab) > wire1675))))};
              reg1694 = (+(^(~|(((7'h44) ?
                  reg1687 : reg1693) == reg1689[(3'h5):(3'h4)]))));
              reg1695 <= $signed((reg1682[(1'h1):(1'h0)] ?
                  (((+forvar1683) != ((8'h9f) ?
                      (8'hab) : reg1691)) && forvar1690) : wire1675));
              reg1696 <= (forvar1690 & (reg1694[(1'h1):(1'h0)] ?
                  reg1691[(2'h2):(1'h0)] : ("RZT1NZFWs4xayWH1LpCXSQ6e" != "L1XriKdmcz")));
            end
          for (forvar1697 = (1'h0); (forvar1697 < (3'h4)); forvar1697 = (forvar1697 + (1'h1)))
            begin
              for (forvar1698 = (1'h0); (forvar1698 < (1'h0)); forvar1698 = (forvar1698 + (1'h1)))
                begin
                  reg1699 = (^~(reg1686[(2'h3):(2'h2)] || ({reg1685[(3'h6):(2'h3)]} ?
                      "8o0BSV5XnbBCmt6mOLr05ud6s" : forvar1688)));
                  reg1700 <= wire1677;
                  reg1701 <= (({$unsigned({forvar1690, reg1692}),
                          (~|$unsigned(reg1695))} != forvar1688) ?
                      "RAagNycXQ0DZHKpAGHgx" : "sNwing08G4ec");
                end
              reg1702 <= "qhoAkkptGL2PMxTtHHWq";
            end
        end
      else
        begin
          reg1685 = (~&((7'h47) ?
              $unsigned(forvar1688) : ($signed((reg1681 ?
                  reg1695 : reg1684)) <<< forvar1690)));
          for (forvar1686 = (1'h0); (forvar1686 < (1'h1)); forvar1686 = (forvar1686 + (1'h1)))
            begin
              reg1687 <= ((reg1694 > reg1692) ?
                  $signed(reg1699[(1'h0):(1'h0)]) : {(+({wire1680} ?
                          "elLqyZWmFJ1uRJKklwi8l" : (-forvar1690))),
                      $signed("3cgzRD68")});
              reg1688 <= forvar1698;
              reg1689 = wire1679[(4'ha):(3'h4)];
              reg1690 <= {$unsigned({{(reg1699 || wire1679)}, wire1680}),
                  forvar1698[(2'h3):(1'h1)]};
              reg1691 <= {$unsigned(($signed(reg1701[(1'h1):(1'h1)]) || $signed((-reg1691)))),
                  "odoN"};
            end
          reg1692 <= (^~{reg1700[(3'h4):(2'h2)]});
          reg1693 <= (~^{{"eeNS3wRNQCRAGeOIRv"}, reg1696});
          reg1694 <= (~wire1680);
          reg1695 = forvar1686[(1'h1):(1'h0)];
        end
    end
  assign wire1703 = "Ap7nTn3Lg";
  always
    @(posedge clk) begin
      reg1704 = $signed((^~($signed(reg1687[(3'h6):(3'h6)]) ?
          ((reg1696 ?
              forvar1690 : reg1690) != reg1681[(4'hc):(3'h6)]) : $unsigned((wire1676 ?
              reg1684 : reg1695)))));
      reg1705 <= ("WgrH" ^ ((8'ha2) < $signed(reg1691)));
    end
  always
    @(posedge clk) begin
      reg1706 = $unsigned((wire1676[(1'h0):(1'h0)] > $signed("c21G")));
      for (forvar1707 = (1'h0); (forvar1707 < (2'h2)); forvar1707 = (forvar1707 + (1'h1)))
        begin
          reg1708 <= ((7'h4c) >= $unsigned((7'h4e)));
          reg1709 <= (8'hb6);
          reg1710 <= $unsigned("1kVcRScrmhV3SLFaxe");
          for (forvar1711 = (1'h0); (forvar1711 < (3'h4)); forvar1711 = (forvar1711 + (1'h1)))
            begin
              reg1712 <= reg1705[(4'hb):(3'h4)];
              reg1713 <= reg1695[(3'h5):(3'h4)];
              reg1714 <= $signed((|(7'h40)));
              reg1715 = {("EgsYYziBEylBc" & (&$unsigned("8vxJbq"))),
                  wire1678[(3'h5):(1'h1)]};
              reg1716 <= reg1700[(1'h1):(1'h0)];
            end
        end
    end
  assign wire1717 = $signed(reg1714[(5'h11):(2'h2)]);
  always
    @(posedge clk) begin
      for (forvar1718 = (1'h0); (forvar1718 < (3'h5)); forvar1718 = (forvar1718 + (1'h1)))
        begin
          reg1719 <= "ncO8B9IKk31wh2a6";
          reg1720 <= (8'hbb);
          reg1721 = forvar1686[(2'h3):(1'h0)];
          for (forvar1722 = (1'h0); (forvar1722 < (3'h4)); forvar1722 = (forvar1722 + (1'h1)))
            begin
              reg1723 <= "PDsR7qRqGh";
              reg1724 <= $unsigned("NT9E0AkkhdoQR3W6JOO8");
              reg1725 <= forvar1718;
              for (forvar1726 = (1'h0); (forvar1726 < (3'h4)); forvar1726 = (forvar1726 + (1'h1)))
                begin
                  reg1727 <= "KOTneBziTI";
                  reg1728 <= {wire1717, reg1705[(4'h8):(2'h2)]};
                  reg1729 <= "b1aM6ds19SuChVeZ7f9gNI6wR";
                  reg1730 <= (!((((reg1691 ? (8'ha4) : forvar1686) ?
                          (-(8'hac)) : reg1704) ?
                      reg1699 : ((reg1687 * (8'haa)) == "cPT1BPEtgtERMD0H")) < reg1684[(5'h11):(3'h4)]));
                end
              reg1731 = ("" ?
                  (~&$signed(reg1699[(1'h1):(1'h0)])) : $unsigned((("rLNC31tnQTVefJhk14" ?
                          "Eh7U927uo7kG0COo5Jfh" : $unsigned((8'h9c))) ?
                      ($unsigned(reg1720) || $signed(forvar1697)) : reg1728[(5'h10):(4'hc)])));
              reg1732 <= $unsigned((~^reg1691[(1'h0):(1'h0)]));
            end
        end
      reg1733 <= (|$signed("q6DHW4bn8wKGlkBd"));
    end
  always
    @(posedge clk) begin
      for (forvar1734 = (1'h0); (forvar1734 < (2'h2)); forvar1734 = (forvar1734 + (1'h1)))
        begin
          reg1735 <= $signed((reg1696 ?
              ($unsigned({forvar1734}) ?
                  ($signed(reg1712) || (&reg1694)) : (reg1701[(3'h4):(3'h4)] ?
                      {wire1717, reg1704} : reg1689)) : (-((reg1685 | reg1728) ?
                  (forvar1688 & forvar1734) : reg1690[(3'h6):(2'h2)]))));
        end
      for (forvar1736 = (1'h0); (forvar1736 < (3'h5)); forvar1736 = (forvar1736 + (1'h1)))
        begin
          reg1737 <= ((reg1719 ?
                  wire1678 : $signed((wire1675[(4'hc):(4'h8)] ?
                      forvar1722 : (reg1721 ? reg1716 : reg1733)))) ?
              $signed($signed($signed("Tg"))) : $signed($signed("EB0UHCm")));
          reg1738 = (^$signed(reg1732));
          reg1739 = forvar1722[(5'h13):(5'h12)];
          reg1740 <= $signed((-forvar1734));
        end
      for (forvar1741 = (1'h0); (forvar1741 < (3'h5)); forvar1741 = (forvar1741 + (1'h1)))
        begin
          reg1742 <= reg1715;
          reg1743 = (~^$signed($signed(reg1737[(2'h3):(1'h0)])));
          for (forvar1744 = (1'h0); (forvar1744 < (3'h5)); forvar1744 = (forvar1744 + (1'h1)))
            begin
              reg1745 <= (~&reg1738);
              reg1746 <= ((reg1682 >= (|(((8'h9c) ?
                      forvar1707 : reg1682) + (~forvar1683)))) ?
                  reg1740[(4'hb):(3'h7)] : forvar1736);
            end
          for (forvar1747 = (1'h0); (forvar1747 < (2'h2)); forvar1747 = (forvar1747 + (1'h1)))
            begin
              reg1748 = (reg1743 ? forvar1688[(2'h2):(2'h2)] : "GQWzqIV");
              reg1749 <= reg1720;
            end
        end
      reg1750 <= $unsigned($signed("ni0DVv"));
      reg1751 <= ((^"yRUCAQhplE2siZXG") ?
          ({((wire1677 ? reg1714 : (7'h43)) ?
                      forvar1734 : reg1710[(4'hc):(1'h1)]),
                  "NPbMH"} ?
              (^$unsigned((reg1702 ?
                  (7'h48) : reg1746))) : $unsigned((|(reg1690 - reg1694)))) : (^~(-{$signed(reg1687)})));
    end
  assign wire1752 = (8'ha8);
  always
    @(posedge clk) begin
      reg1753 <= $signed(reg1694[(3'h6):(3'h4)]);
    end
  assign wire1754 = reg1720[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar1755 = (1'h0); (forvar1755 < (2'h2)); forvar1755 = (forvar1755 + (1'h1)))
        begin
          reg1756 <= ((8'hb3) ? ("htFF" * {$unsigned((^wire1703))}) : (^"7oO"));
          reg1757 = $signed($unsigned((reg1708 ?
              reg1695[(3'h6):(3'h5)] : "KEkxxWuGPX")));
          reg1758 = ($unsigned((!((^reg1723) ^ "12CHUN3DH8"))) ^~ ($signed(("SQWbWRcRmGEI9cMYeVtLVP" > reg1733[(1'h0):(1'h0)])) ?
              forvar1690 : reg1706));
          reg1759 <= (~^wire1754);
        end
    end
  always
    @(posedge clk) begin
      reg1760 = (~|$signed((reg1750 + (reg1695[(4'h9):(1'h1)] ?
          (reg1714 ? forvar1734 : reg1753) : (reg1699 ?
              (7'h4e) : forvar1686)))));
      reg1761 = (reg1695[(4'ha):(4'ha)] && (-{$signed(reg1757[(4'h9):(1'h0)]),
          ((|forvar1726) || $signed(reg1689))}));
      reg1762 <= ("dZZCk9edUcNdS" ?
          $unsigned((8'ha0)) : {$unsigned("Qz37"),
              $signed(wire1677[(5'h15):(4'hb)])});
      reg1763 <= {"yimnfeLzdipzeAbU2x"};
    end
  assign wire1764 = "71M";
  always
    @(posedge clk) begin
      reg1765 <= (wire1764[(3'h4):(2'h3)] >>> {$signed(reg1729)});
      reg1766 <= ($signed({$signed((reg1725 ? reg1706 : reg1724)),
              ("" ? $unsigned(forvar1686) : forvar1688[(5'h15):(4'h8)])}) ?
          ($unsigned(reg1682[(1'h0):(1'h0)]) ?
              reg1749 : "eIaWG") : reg1765[(4'ha):(3'h7)]);
    end
  always
    @(posedge clk) begin
      for (forvar1767 = (1'h0); (forvar1767 < (3'h4)); forvar1767 = (forvar1767 + (1'h1)))
        begin
          reg1768 = ((forvar1736[(4'ha):(4'h8)] != (~forvar1688)) ?
              (^(reg1732 ?
                  reg1735 : "yrYoeKrpsNESH")) : $unsigned(("qHCi5Cd9Rdl1VaifBhd4P" >= {$unsigned(reg1762)})));
        end
    end
  assign wire1769 = forvar1690[(4'h9):(4'h9)];
  always
    @(posedge clk) begin
      reg1770 <= ($signed($signed(reg1728[(4'hf):(4'hc)])) ?
          $signed($unsigned(({(8'ha6), forvar1686} ~^ (forvar1718 ?
              reg1746 : reg1762)))) : ($signed(($signed(reg1693) ^ (+wire1717))) >= reg1750));
      for (forvar1771 = (1'h0); (forvar1771 < (1'h0)); forvar1771 = (forvar1771 + (1'h1)))
        begin
          reg1772 = ((reg1762[(4'h9):(1'h1)] ?
                  (&reg1692[(2'h3):(1'h0)]) : (forvar1747[(5'h10):(4'ha)] >>> $signed("yEqZadQwxAg0EpV8FnSr"))) ?
              reg1700 : reg1701);
          reg1773 <= reg1727[(2'h3):(2'h2)];
        end
      for (forvar1774 = (1'h0); (forvar1774 < (2'h2)); forvar1774 = (forvar1774 + (1'h1)))
        begin
          reg1775 <= reg1706[(3'h7):(2'h3)];
          reg1776 <= ($unsigned($signed(reg1773)) ?
              ((~|forvar1690[(2'h2):(1'h1)]) ?
                  (forvar1718[(4'h8):(1'h0)] * reg1737) : reg1724) : $unsigned((7'h4a)));
        end
    end
  always
    @(posedge clk) begin
      reg1777 <= $unsigned(($unsigned(forvar1734) ? $unsigned(reg1692) : "o"));
      reg1778 <= {forvar1734[(1'h1):(1'h0)]};
      for (forvar1779 = (1'h0); (forvar1779 < (3'h4)); forvar1779 = (forvar1779 + (1'h1)))
        begin
          reg1780 <= $signed((8'hb1));
          for (forvar1781 = (1'h0); (forvar1781 < (2'h2)); forvar1781 = (forvar1781 + (1'h1)))
            begin
              reg1782 <= ($signed($signed((~&reg1710))) == "JTKJO0wM");
              if ($unsigned(wire1680))
                begin
                  reg1783 = (&reg1760[(5'h13):(5'h13)]);
                end
              else
                begin
                  reg1783 = ((!$unsigned("APLaB5hcAm0Ve7hHWe0CsL8US")) | (|reg1687));
                  reg1784 <= "09usW3cOQZ3";
                end
              reg1785 <= $unsigned(forvar1736[(3'h5):(1'h0)]);
              reg1786 <= (7'h41);
            end
          reg1787 <= $unsigned(reg1713);
        end
      for (forvar1788 = (1'h0); (forvar1788 < (3'h4)); forvar1788 = (forvar1788 + (1'h1)))
        begin
          for (forvar1789 = (1'h0); (forvar1789 < (1'h1)); forvar1789 = (forvar1789 + (1'h1)))
            begin
              reg1790 <= reg1693;
              reg1791 <= "lXe6Ktrl";
            end
          reg1792 <= reg1772[(2'h3):(2'h3)];
          reg1793 <= "Oz2JytDryzNtnRQLPAxTl";
          reg1794 <= (^~reg1750);
          reg1795 <= $unsigned((8'hb4));
        end
    end
  assign wire1796 = reg1727[(2'h3):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar1797 = (1'h0); (forvar1797 < (2'h3)); forvar1797 = (forvar1797 + (1'h1)))
        begin
          reg1798 <= (~&reg1704[(3'h4):(1'h1)]);
          reg1799 <= reg1763;
          reg1800 = (+reg1795[(4'h8):(2'h2)]);
          reg1801 <= (wire1679 ?
              reg1729[(4'h9):(1'h0)] : ((|$signed(reg1758)) == ("" || reg1733)));
        end
      reg1802 <= (^reg1751[(3'h5):(2'h3)]);
      for (forvar1803 = (1'h0); (forvar1803 < (1'h1)); forvar1803 = (forvar1803 + (1'h1)))
        begin
          for (forvar1804 = (1'h0); (forvar1804 < (3'h4)); forvar1804 = (forvar1804 + (1'h1)))
            begin
              reg1805 <= "bAwimuVkeHIOOs8zVRpvT96";
              reg1806 = ($unsigned(reg1773[(3'h5):(2'h3)]) ?
                  $unsigned($unsigned(forvar1736)) : (reg1783[(1'h1):(1'h1)] * forvar1726));
            end
          reg1807 <= ("b9WJEw9ssyPbDUtg6VXSsAdg" ^~ $signed((((reg1778 >> wire1754) - (reg1738 ?
              wire1717 : reg1714)) == $signed("fGgZZvWRUXh27NqMOm8tNH9Gz"))));
          for (forvar1808 = (1'h0); (forvar1808 < (2'h2)); forvar1808 = (forvar1808 + (1'h1)))
            begin
              for (forvar1809 = (1'h0); (forvar1809 < (3'h5)); forvar1809 = (forvar1809 + (1'h1)))
                begin
                  reg1810 <= "PEFW1";
                  reg1811 <= ($unsigned($unsigned(forvar1789[(3'h6):(2'h3)])) ?
                      $unsigned(reg1756[(1'h0):(1'h0)]) : {(-reg1695[(3'h5):(3'h5)]),
                          ($unsigned((forvar1804 & forvar1788)) || $signed((~^reg1798)))});
                  reg1812 <= (|reg1756[(2'h2):(1'h1)]);
                  reg1813 = {(!reg1748[(4'hd):(3'h6)]),
                      (((~|$unsigned(wire1717)) ?
                              $signed(((8'haa) ?
                                  reg1738 : reg1806)) : reg1732[(3'h5):(3'h5)]) ?
                          ("s6dgRIJMnycFN6O" ?
                              forvar1771 : (wire1717 >>> (reg1748 | reg1699))) : reg1784[(3'h6):(3'h4)])};
                  reg1814 = ($unsigned(reg1723[(1'h0):(1'h0)]) ?
                      ((!((~&(8'ha3)) ? wire1717 : "1w")) ?
                          reg1806 : {$unsigned((reg1745 ?
                                  reg1738 : reg1800))}) : ("ywtP" ?
                          ((reg1708 ?
                              "QQqCG5HiXMgPIdIqgmz" : $signed(reg1753)) | ((reg1773 - reg1790) ^~ "")) : (~^((^~forvar1774) >>> $unsigned(reg1706)))));
                end
              reg1815 = (~^reg1794[(4'hc):(4'hc)]);
              reg1816 <= $unsigned(("6RewKCWTqmpRE" | ("wwN" ?
                  ("TrQq" >>> (reg1750 ?
                      (8'hac) : forvar1804)) : (~&$unsigned(reg1693)))));
              reg1817 <= $signed(($unsigned("") <= {{((8'hb8) ?
                          reg1728 : (8'hbe)),
                      "xhhFvhroI0WhlpS"},
                  reg1699}));
              reg1818 = "gNTCM7adNL";
            end
        end
      reg1819 <= $signed({$signed($unsigned(((7'h4a) ? reg1750 : reg1742))),
          reg1792[(3'h6):(3'h5)]});
      reg1820 <= (^"");
      reg1821 <= reg1753;
    end
  always
    @(posedge clk) begin
      for (forvar1822 = (1'h0); (forvar1822 < (3'h4)); forvar1822 = (forvar1822 + (1'h1)))
        begin
          reg1823 <= $signed(forvar1718);
        end
      reg1824 <= $signed(reg1806[(3'h4):(2'h2)]);
      reg1825 <= (^reg1748[(4'h9):(2'h3)]);
      reg1826 <= (reg1823 >>> $signed(((^~(reg1816 ~^ reg1733)) | forvar1789)));
    end
  always
    @(posedge clk) begin
      for (forvar1827 = (1'h0); (forvar1827 < (1'h0)); forvar1827 = (forvar1827 + (1'h1)))
        begin
          reg1828 <= (8'ha4);
          reg1829 = {"nDlMyoV9FT7", "a"};
          reg1830 <= $signed(forvar1711);
        end
      reg1831 <= ($signed((((+(7'h46)) ?
              {reg1791} : "zyJIVLNG") < $unsigned($unsigned(reg1791)))) ?
          $unsigned(reg1682) : $signed((~|reg1710)));
      reg1832 <= $unsigned(({("3T7nsmXnJKZQgTU" * reg1738[(4'h8):(1'h0)])} ?
          (~&((~&reg1830) ?
              forvar1722[(5'h17):(4'ha)] : {reg1716, reg1807})) : ((reg1762 ?
                  forvar1736 : reg1800[(4'h9):(2'h3)]) ?
              "v5" : "2IfmEwSxocLoSSxDTg")));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1483  (y, clk, wire1487, wire1486, wire1485, wire1484);
  output wire [(32'haa1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire1487;
  input wire [(5'h11):(1'h0)] wire1486;
  input wire signed [(5'h19):(1'h0)] wire1485;
  input wire [(3'h5):(1'h0)] wire1484;
  reg signed [(3'h5):(1'h0)] reg1671 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1670 = (1'h0);
  reg [(5'h13):(1'h0)] reg1669 = (1'h0);
  reg [(5'h17):(1'h0)] reg1668 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1667 = (1'h0);
  wire [(4'hc):(1'h0)] wire1666;
  reg signed [(3'h6):(1'h0)] reg1665 = (1'h0);
  reg [(5'h12):(1'h0)] reg1664 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1642 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1663 = (1'h0);
  reg [(5'h19):(1'h0)] reg1662 = (1'h0);
  reg [(5'h16):(1'h0)] reg1661 = (1'h0);
  reg [(5'h12):(1'h0)] reg1660 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1659 = (1'h0);
  reg [(5'h12):(1'h0)] reg1658 = (1'h0);
  reg [(5'h15):(1'h0)] reg1657 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1656 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1655 = (1'h0);
  reg [(4'h8):(1'h0)] reg1654 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1653 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1652 = (1'h0);
  reg [(2'h3):(1'h0)] reg1651 = (1'h0);
  reg [(4'h8):(1'h0)] reg1650 = (1'h0);
  reg [(4'ha):(1'h0)] reg1649 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1648 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1647 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1646 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1645 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1644 = (1'h0);
  reg [(3'h7):(1'h0)] reg1643 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1642 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1641 = (1'h0);
  reg [(5'h13):(1'h0)] reg1640 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1639 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1638 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1637 = (1'h0);
  reg [(4'h9):(1'h0)] reg1636 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1635 = (1'h0);
  reg [(5'h14):(1'h0)] reg1634 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1633 = (1'h0);
  reg [(5'h17):(1'h0)] reg1632 = (1'h0);
  reg [(3'h7):(1'h0)] reg1631 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1630 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1629 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1628 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1627 = (1'h0);
  reg [(2'h3):(1'h0)] reg1626 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1625 = (1'h0);
  reg [(4'hb):(1'h0)] reg1624 = (1'h0);
  reg [(5'h10):(1'h0)] reg1623 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1622 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1621 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1620 = (1'h0);
  reg [(5'h17):(1'h0)] reg1619 = (1'h0);
  reg [(5'h10):(1'h0)] reg1618 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1617 = (1'h0);
  reg [(5'h15):(1'h0)] reg1616 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1615 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1614 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1613 = (1'h0);
  reg [(2'h2):(1'h0)] reg1612 = (1'h0);
  reg [(3'h5):(1'h0)] reg1611 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1610 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1609 = (1'h0);
  reg [(4'hb):(1'h0)] reg1608 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1607 = (1'h0);
  reg [(4'h9):(1'h0)] reg1606 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1605 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1604 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1603 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1602 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire1601;
  reg signed [(4'hd):(1'h0)] reg1600 = (1'h0);
  reg [(2'h3):(1'h0)] reg1599 = (1'h0);
  reg [(3'h5):(1'h0)] reg1598 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1597 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1596 = (1'h0);
  reg [(2'h3):(1'h0)] reg1595 = (1'h0);
  reg [(5'h16):(1'h0)] reg1594 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1593 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1592 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1591 = (1'h0);
  reg [(5'h11):(1'h0)] reg1590 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1589 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1588 = (1'h0);
  reg [(4'he):(1'h0)] reg1587 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1586 = (1'h0);
  reg [(4'he):(1'h0)] forvar1585 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1584 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1583 = (1'h0);
  reg [(4'he):(1'h0)] reg1582 = (1'h0);
  reg [(5'h16):(1'h0)] reg1581 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire1580;
  reg [(3'h5):(1'h0)] reg1579 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1578 = (1'h0);
  reg [(2'h3):(1'h0)] reg1577 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1576 = (1'h0);
  reg [(5'h16):(1'h0)] reg1575 = (1'h0);
  reg [(3'h5):(1'h0)] reg1574 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1573 = (1'h0);
  reg [(3'h7):(1'h0)] reg1572 = (1'h0);
  reg [(3'h6):(1'h0)] reg1571 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1570 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1569 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1568 = (1'h0);
  reg [(5'h15):(1'h0)] reg1567 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1566 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1565 = (1'h0);
  reg [(5'h12):(1'h0)] reg1564 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1563 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1562 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1561 = (1'h0);
  reg [(4'ha):(1'h0)] reg1560 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1559 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1558 = (1'h0);
  wire [(5'h16):(1'h0)] wire1557;
  reg [(3'h4):(1'h0)] reg1556 = (1'h0);
  reg [(4'h8):(1'h0)] reg1555 = (1'h0);
  wire [(4'hf):(1'h0)] wire1554;
  reg [(5'h15):(1'h0)] reg1553 = (1'h0);
  reg [(4'h8):(1'h0)] reg1552 = (1'h0);
  reg [(5'h19):(1'h0)] reg1551 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1550 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1549 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1548 = (1'h0);
  reg [(2'h3):(1'h0)] reg1547 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1546 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1545 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1544 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1543 = (1'h0);
  reg [(5'h16):(1'h0)] reg1542 = (1'h0);
  reg [(5'h16):(1'h0)] reg1541 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1540 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1539 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1538 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1537 = (1'h0);
  reg [(5'h10):(1'h0)] reg1536 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1535 = (1'h0);
  reg [(2'h2):(1'h0)] reg1534 = (1'h0);
  reg [(4'hc):(1'h0)] reg1533 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1532 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1531 = (1'h0);
  wire signed [(5'h18):(1'h0)] wire1530;
  reg signed [(5'h17):(1'h0)] reg1529 = (1'h0);
  reg [(5'h13):(1'h0)] reg1528 = (1'h0);
  reg [(4'hd):(1'h0)] reg1527 = (1'h0);
  reg [(5'h17):(1'h0)] reg1526 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1525 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1524 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1523 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1522 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1521 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1520 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1519 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1518 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1517 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1516 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1515 = (1'h0);
  reg [(2'h2):(1'h0)] reg1514 = (1'h0);
  reg [(3'h6):(1'h0)] reg1513 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1512 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1511 = (1'h0);
  reg [(4'ha):(1'h0)] reg1510 = (1'h0);
  reg [(5'h15):(1'h0)] reg1509 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1508 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1507 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1506 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1504 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1502 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1505 = (1'h0);
  reg [(4'hb):(1'h0)] reg1504 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1503 = (1'h0);
  reg [(3'h7):(1'h0)] reg1502 = (1'h0);
  reg [(5'h11):(1'h0)] reg1501 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1500 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1499 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1498 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1497 = (1'h0);
  reg [(3'h4):(1'h0)] reg1496 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1495 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1494 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1493 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1492 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1491 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1490 = (1'h0);
  reg [(5'h12):(1'h0)] reg1489 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1488 = (1'h0);
  assign y = {reg1671,
                 reg1670,
                 reg1669,
                 reg1668,
                 forvar1667,
                 wire1666,
                 reg1665,
                 reg1664,
                 reg1642,
                 reg1663,
                 reg1662,
                 reg1661,
                 reg1660,
                 reg1659,
                 reg1658,
                 reg1657,
                 reg1656,
                 forvar1655,
                 reg1654,
                 forvar1653,
                 reg1652,
                 reg1651,
                 reg1650,
                 reg1649,
                 reg1648,
                 reg1647,
                 reg1646,
                 reg1645,
                 forvar1644,
                 reg1643,
                 forvar1642,
                 reg1641,
                 reg1640,
                 reg1639,
                 reg1638,
                 forvar1637,
                 reg1636,
                 reg1635,
                 reg1634,
                 forvar1633,
                 reg1632,
                 reg1631,
                 reg1630,
                 forvar1629,
                 reg1628,
                 forvar1627,
                 reg1626,
                 forvar1625,
                 reg1624,
                 reg1623,
                 reg1622,
                 reg1621,
                 reg1620,
                 reg1619,
                 reg1618,
                 forvar1617,
                 reg1616,
                 reg1615,
                 reg1614,
                 reg1613,
                 reg1612,
                 reg1611,
                 reg1610,
                 forvar1609,
                 reg1608,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1604,
                 reg1603,
                 forvar1602,
                 wire1601,
                 reg1600,
                 reg1599,
                 reg1598,
                 reg1597,
                 forvar1596,
                 reg1595,
                 reg1594,
                 reg1593,
                 forvar1592,
                 forvar1591,
                 reg1590,
                 forvar1589,
                 reg1588,
                 reg1587,
                 reg1586,
                 forvar1585,
                 reg1584,
                 reg1583,
                 reg1582,
                 reg1581,
                 wire1580,
                 reg1579,
                 reg1578,
                 reg1577,
                 reg1576,
                 reg1575,
                 reg1574,
                 forvar1573,
                 reg1572,
                 reg1571,
                 reg1570,
                 reg1569,
                 reg1568,
                 reg1567,
                 forvar1566,
                 forvar1565,
                 reg1564,
                 reg1563,
                 forvar1562,
                 reg1561,
                 reg1560,
                 reg1559,
                 reg1558,
                 wire1557,
                 reg1556,
                 reg1555,
                 wire1554,
                 reg1553,
                 reg1552,
                 reg1551,
                 reg1550,
                 reg1549,
                 forvar1548,
                 reg1547,
                 reg1546,
                 reg1545,
                 reg1544,
                 reg1543,
                 reg1542,
                 reg1541,
                 reg1540,
                 reg1539,
                 forvar1538,
                 reg1537,
                 reg1536,
                 forvar1535,
                 reg1534,
                 reg1533,
                 reg1532,
                 forvar1531,
                 wire1530,
                 reg1529,
                 reg1528,
                 reg1527,
                 reg1526,
                 reg1525,
                 reg1524,
                 reg1523,
                 reg1522,
                 reg1521,
                 forvar1520,
                 reg1519,
                 forvar1518,
                 reg1517,
                 reg1516,
                 reg1515,
                 reg1514,
                 reg1513,
                 forvar1512,
                 forvar1511,
                 reg1510,
                 reg1509,
                 reg1508,
                 reg1507,
                 reg1506,
                 forvar1504,
                 forvar1502,
                 reg1505,
                 reg1504,
                 reg1503,
                 reg1502,
                 reg1501,
                 reg1500,
                 reg1499,
                 reg1498,
                 reg1497,
                 reg1496,
                 reg1495,
                 reg1494,
                 reg1493,
                 reg1492,
                 reg1491,
                 reg1490,
                 reg1489,
                 forvar1488,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar1488 = (1'h0); (forvar1488 < (1'h1)); forvar1488 = (forvar1488 + (1'h1)))
        begin
          reg1489 <= $signed(("07NP" <= {"AU76Ie"}));
          reg1490 <= $unsigned($signed("HJT3ZXR6NUozeZMCWa6mDQ2w2"));
          reg1491 = (reg1490[(3'h7):(2'h3)] != $signed((reg1490 ?
              (wire1485[(5'h15):(5'h11)] || "o53FyLBGUPTL") : reg1489[(4'hf):(4'h9)])));
          reg1492 <= wire1486;
          reg1493 <= forvar1488;
          reg1494 <= (&(-$unsigned(($unsigned((8'haa)) ^~ $unsigned(reg1490)))));
        end
      reg1495 <= (+("W" ? reg1490 : wire1486[(2'h3):(2'h2)]));
      reg1496 <= ("V4AihNZ7" ^ (!(~$unsigned("6faP"))));
      reg1497 <= {$unsigned((($signed(wire1485) ?
                  $unsigned(reg1494) : "irxqD") ?
              ($signed(reg1495) ?
                  wire1487 : ((7'h46) >> reg1489)) : reg1489[(5'h11):(2'h3)])),
          {(reg1490 ? wire1487 : reg1495[(5'h14):(4'ha)])}};
      reg1498 <= reg1497;
      reg1499 = {wire1484[(3'h5):(3'h4)],
          ("kzsLmW0pRAGT31" && {$signed((|(7'h47))),
              ({reg1494, reg1491} ~^ "GYTzJMcxUaTMqZyIRcmpfgm")})};
    end
  always
    @(posedge clk) begin
      reg1500 <= "2q";
      if (reg1494[(5'h10):(4'ha)])
        begin
          reg1501 <= (reg1500 ?
              $unsigned((~&{$signed(wire1484),
                  reg1491})) : "BoDIROubP3bIUZAGlzUhI1eVQ");
          reg1502 <= ($signed({wire1487,
              $signed($signed(reg1492))}) <= (({$unsigned(reg1493),
                  $signed(reg1492)} <<< (wire1486 ?
                  $signed(reg1492) : "xkZ0XqyLBMuWU0")) ?
              "Dia8EgKVpCbZ3" : $signed(forvar1488)));
          reg1503 <= "IpTYs8uBFm4sGGpDL";
          reg1504 <= (8'hbe);
          reg1505 <= reg1503[(4'ha):(3'h5)];
        end
      else
        begin
          reg1501 <= ($signed((8'hbf)) && $unsigned((~($signed((8'ha6)) ?
              reg1493[(4'he):(3'h7)] : reg1495[(4'hb):(3'h6)]))));
          for (forvar1502 = (1'h0); (forvar1502 < (1'h0)); forvar1502 = (forvar1502 + (1'h1)))
            begin
              reg1503 = {("0duzbcrMNXYtQoCwdFt" ?
                      $signed(((wire1484 ^ reg1489) ^~ (forvar1488 <= wire1486))) : "HOv1Wa5ns4"),
                  reg1501[(5'h11):(1'h0)]};
              for (forvar1504 = (1'h0); (forvar1504 < (3'h5)); forvar1504 = (forvar1504 + (1'h1)))
                begin
                  reg1505 <= reg1491[(1'h0):(1'h0)];
                  reg1506 = wire1487[(3'h5):(1'h0)];
                  reg1507 <= reg1504;
                end
              reg1508 <= reg1489;
            end
        end
      reg1509 <= "g8Q7mbKDiQIwRAoYntemcQS";
      reg1510 = $unsigned(reg1491[(3'h4):(3'h4)]);
      for (forvar1511 = (1'h0); (forvar1511 < (3'h4)); forvar1511 = (forvar1511 + (1'h1)))
        begin
          for (forvar1512 = (1'h0); (forvar1512 < (3'h5)); forvar1512 = (forvar1512 + (1'h1)))
            begin
              reg1513 <= (((^~reg1491[(2'h3):(1'h1)]) ?
                  reg1495[(5'h12):(4'h8)] : ($unsigned((^~reg1505)) ?
                      $signed($unsigned(reg1501)) : "vcwwwWwYSB")) - (8'hac));
              reg1514 = ((($unsigned("C") ?
                      $unsigned(reg1503) : reg1493) >> "Oi5EhD5dyb3h622") ?
                  $unsigned(reg1500[(4'h8):(1'h1)]) : (+$signed(reg1504[(3'h7):(1'h0)])));
            end
          reg1515 <= "ZTCXEhENeksRUYHVgnxCwE";
          reg1516 <= "1sWvJa0xKS";
          reg1517 <= "V8dtQFfFyJZMMBJehKn";
        end
    end
  always
    @(posedge clk) begin
      for (forvar1518 = (1'h0); (forvar1518 < (1'h1)); forvar1518 = (forvar1518 + (1'h1)))
        begin
          reg1519 <= ((reg1496 - ($signed($unsigned(wire1485)) ?
              (&reg1504) : reg1514[(1'h1):(1'h0)])) > (8'hae));
          for (forvar1520 = (1'h0); (forvar1520 < (2'h3)); forvar1520 = (forvar1520 + (1'h1)))
            begin
              reg1521 <= $unsigned(($unsigned({(reg1493 & reg1515)}) ?
                  $signed($unsigned((^reg1493))) : $unsigned("v8ZGHvXJbMu")));
              reg1522 = (forvar1504[(2'h2):(1'h0)] ?
                  ({$signed(forvar1518[(1'h1):(1'h0)])} ?
                      (8'h9f) : $signed((reg1514 ?
                          "lBrQs1T0AUF5KdQ" : (reg1513 ?
                              reg1509 : reg1503)))) : "h2hGrmKkPnUYwtfc8g8sO");
              reg1523 <= $unsigned($unsigned($signed({$signed(reg1509)})));
              reg1524 = (7'h4e);
              reg1525 = (&"");
            end
          reg1526 <= $signed($signed((reg1522[(4'he):(4'ha)] && forvar1502)));
          reg1527 = reg1503[(3'h6):(1'h0)];
          reg1528 <= (^((+((wire1486 || wire1487) | $signed(wire1484))) ?
              reg1501[(3'h7):(3'h7)] : reg1499[(4'h9):(4'h8)]));
          reg1529 <= forvar1520[(3'h5):(3'h4)];
        end
    end
  assign wire1530 = {$signed("31Ie"), reg1525};
  always
    @(posedge clk) begin
      for (forvar1531 = (1'h0); (forvar1531 < (1'h1)); forvar1531 = (forvar1531 + (1'h1)))
        begin
          reg1532 <= $signed(reg1519[(1'h0):(1'h0)]);
          reg1533 <= $unsigned(("ogrfOB3v7VJVyZ" ?
              $signed($unsigned(reg1528)) : (((reg1513 | (7'h4b)) ?
                  ((7'h44) < reg1497) : "PorD4Mr") >> "hViDZlzOCKhl7Msp7WQ")));
          reg1534 <= (~^{$signed((8'ha7)), reg1506});
          for (forvar1535 = (1'h0); (forvar1535 < (3'h5)); forvar1535 = (forvar1535 + (1'h1)))
            begin
              reg1536 = "JveFxx";
              reg1537 <= {reg1494, ($unsigned(reg1523) ? reg1523 : forvar1502)};
              for (forvar1538 = (1'h0); (forvar1538 < (3'h4)); forvar1538 = (forvar1538 + (1'h1)))
                begin
                  reg1539 <= "VNDQczbcQXmAJZYlU";
                  reg1540 <= $unsigned(reg1506);
                end
              if ((reg1529 ? $signed(reg1501) : (8'ha0)))
                begin
                  reg1541 = (^reg1496[(3'h4):(3'h4)]);
                end
              else
                begin
                  reg1541 <= ("MiP6sU7l9DhAV8RyB" == $signed(reg1501[(4'hd):(2'h2)]));
                  reg1542 = ((^~{reg1490[(2'h3):(2'h2)]}) ?
                      ((~|forvar1518[(1'h1):(1'h0)]) ?
                          $signed("l9cqm0") : ($signed((reg1524 ?
                              reg1505 : forvar1502)) - "s")) : reg1516[(4'h8):(3'h5)]);
                  reg1543 <= ((!reg1524) >> wire1485[(1'h0):(1'h0)]);
                  reg1544 = reg1495[(2'h2):(1'h1)];
                end
              reg1545 = "F3rcvWmFukoaMTrkdHKvf5qz";
            end
          reg1546 <= ($unsigned("Qkh9fFE27tBamxRNC6wrmUaP1") ?
              $unsigned(($signed($unsigned(reg1501)) ?
                  ("0afla5VEUimEJhkI6" <<< (forvar1502 <<< reg1497)) : $signed($signed(reg1539)))) : reg1501);
          reg1547 <= "MysJ";
        end
      for (forvar1548 = (1'h0); (forvar1548 < (2'h2)); forvar1548 = (forvar1548 + (1'h1)))
        begin
          reg1549 = forvar1538[(1'h0):(1'h0)];
          reg1550 = $signed((reg1517 ?
              (reg1547[(1'h1):(1'h0)] ?
                  {((7'h42) >>> reg1544),
                      $signed(reg1490)} : $signed($unsigned(reg1514))) : (~|(7'h49))));
          reg1551 <= (!$signed((^~(~|reg1496))));
        end
      reg1552 <= reg1544[(4'h9):(3'h5)];
      reg1553 <= (~|"WNh72V7P6z2uMzulzpiq");
    end
  assign wire1554 = $unsigned("MzxdIXwpUglAzpBzaRn8c5");
  always
    @(posedge clk) begin
      reg1555 <= reg1544[(4'hc):(4'h8)];
      reg1556 = $unsigned(reg1526[(3'h7):(3'h5)]);
    end
  assign wire1557 = {"oFRfF"};
  always
    @(posedge clk) begin
      reg1558 = forvar1538;
      reg1559 <= (~$unsigned($unsigned(reg1516[(4'hd):(3'h6)])));
      reg1560 <= (8'ha3);
    end
  always
    @(posedge clk) begin
      reg1561 <= $signed($signed($unsigned(wire1530[(4'hc):(2'h3)])));
      for (forvar1562 = (1'h0); (forvar1562 < (3'h5)); forvar1562 = (forvar1562 + (1'h1)))
        begin
          reg1563 <= {($unsigned(forvar1531[(3'h6):(2'h3)]) * "IEDRPbELk64LF"),
              ("7J0X" <<< (8'hb0))};
        end
      reg1564 <= (~|reg1547[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      for (forvar1565 = (1'h0); (forvar1565 < (3'h4)); forvar1565 = (forvar1565 + (1'h1)))
        begin
          for (forvar1566 = (1'h0); (forvar1566 < (3'h5)); forvar1566 = (forvar1566 + (1'h1)))
            begin
              reg1567 <= (((-forvar1518[(1'h0):(1'h0)]) << reg1544) && reg1553[(4'h9):(3'h7)]);
            end
          reg1568 <= $unsigned((|reg1505[(1'h0):(1'h0)]));
          reg1569 = reg1500;
          reg1570 = ($unsigned("WPRiMQ3aHU09DZg8") ?
              (reg1522 ? "a1L8qP6bak1GPrGzBXgbv" : (!reg1515)) : "cwMfS");
          reg1571 <= ({{$signed($unsigned(reg1515)), reg1517},
                  reg1550[(5'h18):(5'h15)]} ?
              reg1541[(5'h15):(5'h14)] : (((((8'ha8) ~^ wire1487) ?
                      (8'ha6) : $signed(reg1528)) ?
                  ((!reg1551) > {reg1500,
                      reg1491}) : "Tqf8rPcsE3Flu") >= reg1545));
          reg1572 <= ("wc" || {{($signed(reg1541) * (!reg1501)),
                  (!((8'haf) ? (8'hb3) : reg1532))}});
        end
      for (forvar1573 = (1'h0); (forvar1573 < (3'h5)); forvar1573 = (forvar1573 + (1'h1)))
        begin
          reg1574 <= (!(^~$signed($unsigned("rlp7thpZJwOc93"))));
        end
      reg1575 <= (("WGwEcRDqrFNipXX" > forvar1502) > (7'h45));
    end
  always
    @(posedge clk) begin
      reg1576 <= "5gX4";
      reg1577 <= ($signed((-($signed(reg1523) | reg1560[(1'h0):(1'h0)]))) ?
          $unsigned($signed(($signed(reg1576) ^ {wire1557}))) : $signed("GuyvU9zh4fu1cGFZ"));
      reg1578 = (-reg1524[(4'hf):(1'h0)]);
      reg1579 <= reg1576;
    end
  assign wire1580 = $signed($unsigned($unsigned(wire1484)));
  always
    @(posedge clk) begin
      reg1581 <= ({(~forvar1562[(4'he):(4'hd)])} | "9RDh1Imt0SO2qifN");
      reg1582 <= $signed(reg1494);
    end
  always
    @(posedge clk) begin
      reg1583 <= (("V3s8o" * reg1541) ?
          $signed($unsigned(forvar1562[(1'h1):(1'h0)])) : $signed(("" ?
              "P9xVpOUD9Su8qn1NGVary" : reg1560)));
      reg1584 <= {((reg1522[(4'hb):(4'h9)] != $signed((~&(7'h48)))) || {$signed($signed(reg1528)),
              ($signed(reg1581) + reg1499[(3'h4):(3'h4)])}),
          (+"z85JZZpaoWrnkxu1")};
      for (forvar1585 = (1'h0); (forvar1585 < (3'h5)); forvar1585 = (forvar1585 + (1'h1)))
        begin
          reg1586 = "Eb2";
          reg1587 <= wire1554[(4'ha):(2'h3)];
          reg1588 = ($signed((^~{$unsigned((7'h4e))})) ? reg1560 : (8'hb3));
          for (forvar1589 = (1'h0); (forvar1589 < (2'h3)); forvar1589 = (forvar1589 + (1'h1)))
            begin
              reg1590 <= ((^wire1484[(3'h5):(1'h1)]) == reg1536);
            end
        end
      for (forvar1591 = (1'h0); (forvar1591 < (2'h2)); forvar1591 = (forvar1591 + (1'h1)))
        begin
          for (forvar1592 = (1'h0); (forvar1592 < (3'h4)); forvar1592 = (forvar1592 + (1'h1)))
            begin
              reg1593 <= reg1494[(5'h11):(4'ha)];
            end
          reg1594 <= "UOHSmtN";
          reg1595 <= $unsigned((reg1576 * {reg1547[(1'h1):(1'h1)],
              {(forvar1585 ? reg1510 : reg1524), (!(7'h4b))}}));
        end
      for (forvar1596 = (1'h0); (forvar1596 < (1'h0)); forvar1596 = (forvar1596 + (1'h1)))
        begin
          reg1597 <= ((reg1569 ?
                  forvar1573 : ((~|(forvar1535 != reg1491)) ?
                      $signed(reg1569) : (^forvar1562))) ?
              "wGHVAFZIZO" : "HNSy");
          reg1598 <= {$unsigned("FChnWt")};
          reg1599 <= $unsigned(((^(~|(~^reg1526))) ?
              reg1588[(5'h12):(1'h1)] : "gr"));
          reg1600 <= (~&{(~|"6id2"), forvar1565[(1'h1):(1'h0)]});
        end
    end
  assign wire1601 = (~&{"kyfyOLyY0e2xTeSZdfSL", (7'h47)});
  always
    @(posedge clk) begin
      for (forvar1602 = (1'h0); (forvar1602 < (1'h0)); forvar1602 = (forvar1602 + (1'h1)))
        begin
          reg1603 = (reg1498[(4'h8):(4'h8)] ?
              reg1503[(4'ha):(3'h6)] : reg1568[(1'h0):(1'h0)]);
          reg1604 <= (~^(~$unsigned($signed((reg1560 ? reg1578 : (8'haa))))));
          reg1605 <= "INDhg7Uwx";
          reg1606 = ($signed($signed("LYaWEhJ3aodZCG3dqsb")) ^ reg1529[(4'hd):(1'h1)]);
          reg1607 <= (reg1561[(4'h8):(2'h2)] ?
              (8'h9d) : ((7'h4b) ?
                  (($unsigned(reg1560) ?
                      (reg1491 ?
                          reg1567 : reg1559) : reg1532[(2'h2):(1'h0)]) - reg1521[(4'h9):(4'h8)]) : "F92vtESRUJ"));
          reg1608 = $signed($signed($unsigned(reg1493)));
        end
      for (forvar1609 = (1'h0); (forvar1609 < (3'h5)); forvar1609 = (forvar1609 + (1'h1)))
        begin
          reg1610 <= (~|reg1600[(4'hc):(3'h5)]);
          reg1611 <= {reg1549,
              {(reg1490[(2'h2):(1'h1)] <= (&reg1536)),
                  ("y" ?
                      (^~(reg1550 ? reg1533 : reg1599)) : ({reg1498, reg1597} ?
                          $unsigned(forvar1602) : $unsigned((7'h45))))}};
        end
      reg1612 <= reg1600[(4'hb):(2'h2)];
      reg1613 <= $unsigned(((-$unsigned((reg1604 ?
          reg1491 : reg1544))) << ((~^((7'h4b) | forvar1538)) | (reg1563[(2'h3):(2'h3)] ?
          (~(7'h4b)) : {wire1484, reg1568}))));
    end
  always
    @(posedge clk) begin
      reg1614 <= reg1516[(5'h13):(1'h1)];
      reg1615 <= {"1viLR8vldV1F"};
    end
  always
    @(posedge clk) begin
      reg1616 <= "8ohKud3w8WiJGdSunoctY7K";
      for (forvar1617 = (1'h0); (forvar1617 < (3'h5)); forvar1617 = (forvar1617 + (1'h1)))
        begin
          reg1618 <= $signed(reg1540[(2'h3):(2'h3)]);
          reg1619 = ($unsigned("7ZxDMwSOnWC") ?
              reg1544[(4'ha):(2'h3)] : (&$unsigned(({wire1485, (8'h9d)} ?
                  forvar1589[(4'hb):(1'h0)] : {reg1503, wire1580}))));
          reg1620 <= $signed(forvar1531[(3'h5):(3'h5)]);
          reg1621 <= ("" ? "kHxUzCJVWaV0KJWBTghGG" : "sK");
        end
      reg1622 <= reg1545[(1'h1):(1'h0)];
      reg1623 = (reg1586[(2'h3):(2'h3)] ?
          ({(reg1550[(2'h3):(1'h0)] && wire1487[(2'h3):(1'h1)]),
              "aiKSi7dTv"} >> $signed(reg1615)) : ((($signed(reg1586) & {reg1619,
                  reg1497}) ?
              $unsigned($unsigned((8'h9e))) : $signed($unsigned(reg1595))) > "cQM2q1"));
    end
  always
    @(posedge clk) begin
      reg1624 = reg1515;
      for (forvar1625 = (1'h0); (forvar1625 < (3'h4)); forvar1625 = (forvar1625 + (1'h1)))
        begin
          reg1626 = ($signed($signed($signed(((8'hac) - wire1580)))) ?
              "d5ZLIXHzSSuGUz2AYyAupO7" : {(reg1563[(2'h3):(1'h1)] ?
                      "3" : reg1618)});
          for (forvar1627 = (1'h0); (forvar1627 < (3'h4)); forvar1627 = (forvar1627 + (1'h1)))
            begin
              reg1628 <= (+(|((forvar1538[(1'h0):(1'h0)] <<< {(8'hb9)}) != reg1543)));
              for (forvar1629 = (1'h0); (forvar1629 < (3'h5)); forvar1629 = (forvar1629 + (1'h1)))
                begin
                  reg1630 = "KDNO6KhPcrxfoP";
                  reg1631 <= {"NGriC",
                      ($signed("FVNcFl8DvZMANZaFK") + reg1505[(4'hc):(3'h6)])};
                end
            end
        end
      reg1632 <= ($unsigned($signed(("RuD" && (reg1494 ?
          reg1583 : reg1509)))) >>> {{forvar1562[(2'h2):(2'h2)]},
          (&($unsigned(reg1519) ? $unsigned(reg1624) : {reg1613, reg1586}))});
      for (forvar1633 = (1'h0); (forvar1633 < (2'h2)); forvar1633 = (forvar1633 + (1'h1)))
        begin
          reg1634 <= reg1567[(5'h13):(4'he)];
          reg1635 <= ({$unsigned(({reg1604} ?
                      $signed(forvar1518) : (-forvar1625)))} ?
              (reg1568[(3'h4):(1'h1)] <<< reg1491) : $signed((reg1496[(1'h0):(1'h0)] != ((8'ha6) <= (reg1505 ?
                  reg1551 : reg1614)))));
          reg1636 <= ((8'ha5) - "iWC1cFcARkNu1ewQzz");
          for (forvar1637 = (1'h0); (forvar1637 < (3'h4)); forvar1637 = (forvar1637 + (1'h1)))
            begin
              reg1638 = reg1587;
              reg1639 <= reg1579[(2'h3):(2'h2)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg1640 <= $signed(((reg1497[(1'h1):(1'h0)] * $unsigned((reg1503 >> forvar1511))) ?
          (({reg1631} ?
              (wire1580 ?
                  (8'hb5) : (8'hb5)) : reg1513) == reg1616) : (~^"ZTu1AIoYe7UP")));
    end
  always
    @(posedge clk) begin
      reg1641 <= $signed("mxgHG7WNS79Ya8Urgv8");
    end
  always
    @(posedge clk) begin
      if ($signed(("ppSVTtOnZW" > (($signed(reg1503) ?
              (reg1534 ? reg1612 : reg1590) : "CL97S1bo7o") ?
          ($signed(reg1575) ?
              ((7'h4b) >>> reg1578) : wire1485) : "KXgLys4NLC1Gmlwsvf"))))
        begin
          for (forvar1642 = (1'h0); (forvar1642 < (2'h2)); forvar1642 = (forvar1642 + (1'h1)))
            begin
              reg1643 = $signed((({(reg1496 ?
                      reg1598 : forvar1573)} + ($signed(reg1492) && $signed((8'hb5)))) - (+(-$unsigned(forvar1538)))));
              for (forvar1644 = (1'h0); (forvar1644 < (2'h2)); forvar1644 = (forvar1644 + (1'h1)))
                begin
                  reg1645 <= (+(&(8'hb7)));
                  reg1646 <= "Qe9ce8";
                  reg1647 <= (|(!$signed($unsigned(reg1608[(2'h3):(2'h3)]))));
                  reg1648 <= ((("nccT" ?
                          $signed({reg1575}) : ($unsigned(forvar1538) ^ forvar1504)) <<< {$unsigned(reg1525)}) ?
                      ($unsigned("u") - $signed({(~&(8'hb8)),
                          reg1639})) : $unsigned((7'h44)));
                  reg1649 <= {({((reg1636 ? reg1499 : reg1632) ?
                                  reg1605[(1'h0):(1'h0)] : $signed((8'hb5))),
                              $signed($signed(reg1624))} ?
                          reg1610[(1'h0):(1'h0)] : $unsigned(((reg1515 && reg1583) >= $unsigned((7'h4d))))),
                      reg1555[(3'h6):(2'h2)]};
                  reg1650 = ((^(~^((reg1495 + reg1607) > $unsigned(reg1497)))) + $signed((!((reg1501 <<< reg1499) | "4lUJTWbeJ4zS"))));
                end
              reg1651 <= ($unsigned({(forvar1627[(3'h4):(1'h0)] | reg1504[(3'h7):(2'h2)]),
                  forvar1596[(4'he):(3'h5)]}) - reg1553[(5'h11):(4'hf)]);
              reg1652 <= ($unsigned(reg1525) ~^ $signed($signed(($unsigned(reg1552) ^ reg1567[(5'h15):(5'h13)]))));
            end
          for (forvar1653 = (1'h0); (forvar1653 < (2'h2)); forvar1653 = (forvar1653 + (1'h1)))
            begin
              reg1654 <= (wire1487 ?
                  (|reg1608) : ((reg1628 || {reg1576}) ?
                      (~^"lXnpak4h6LkNv") : reg1648[(4'hb):(3'h7)]));
              for (forvar1655 = (1'h0); (forvar1655 < (1'h0)); forvar1655 = (forvar1655 + (1'h1)))
                begin
                  reg1656 <= (reg1526[(3'h7):(1'h1)] ~^ (8'ha6));
                  reg1657 <= $unsigned("JLYr");
                  reg1658 <= $signed((($signed((reg1534 ? reg1559 : (8'hb2))) ?
                          ((wire1580 ^~ reg1641) >> $signed(reg1491)) : reg1492) ?
                      $signed((!reg1582[(3'h5):(3'h5)])) : forvar1573[(4'ha):(2'h3)]));
                  reg1659 <= wire1557[(3'h6):(3'h4)];
                  reg1660 = wire1484[(1'h0):(1'h0)];
                end
              reg1661 <= ((+(~|forvar1518[(1'h0):(1'h0)])) ?
                  reg1575[(5'h14):(4'hb)] : reg1556[(3'h4):(1'h1)]);
              reg1662 <= forvar1565;
            end
          reg1663 <= $unsigned("QPmT8tH5bKA");
        end
      else
        begin
          reg1642 <= "aIKprn";
        end
      reg1664 = $signed("M5SegUodW0");
      reg1665 <= reg1509;
    end
  assign wire1666 = $signed(((~|"m8DSZRe2qvkOPSZPe") ?
                        (7'h46) : "UibTlq8w60llq4KmUGXNfJ11"));
  always
    @(posedge clk) begin
      for (forvar1667 = (1'h0); (forvar1667 < (3'h4)); forvar1667 = (forvar1667 + (1'h1)))
        begin
          reg1668 <= $unsigned(reg1560);
          reg1669 = $unsigned("6T2eeJTuJ9ubQsrbU");
          reg1670 <= ((&$unsigned({"c2hUxmNTTo0TQTPSUk",
              $signed(reg1584)})) != ((^$unsigned((reg1582 >= forvar1629))) << "38cCWwuwJmz"));
          reg1671 <= $unsigned(({(reg1575 ?
                  (reg1619 ?
                      reg1496 : reg1490) : reg1583[(4'hc):(4'h9)])} != reg1594[(3'h6):(3'h6)]));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1250
#( parameter param1480 = (({({(8'hbf), (7'h46)} && ((7'h46) == (7'h47))), ({(8'hba)} << {(7'h46)})} ? (8'hb1) : (~^{((8'ha6) == (8'haf)), (~^(8'ha6))})) ? {{(((8'hb3) > (8'h9c)) ? (|(8'hba)) : ((8'hb4) ? (8'hbe) : (7'h4c)))}} : ((~&{((7'h49) + (8'h9c)), ((8'haf) ~^ (8'hae))}) * (((+(7'h42)) & (~^(8'hb2))) ? ((~(8'ha1)) - ((8'h9e) >>> (8'ha7))) : (((8'hbf) ? (8'had) : (8'hbc)) ? (^~(8'hbf)) : ((8'hac) ? (7'h4e) : (8'ha1)))))) )
(y, clk, wire1254, wire1253, wire1252, wire1251);
  output wire [(32'hc48):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire1254;
  input wire signed [(5'h13):(1'h0)] wire1253;
  input wire [(4'hf):(1'h0)] wire1252;
  input wire [(3'h5):(1'h0)] wire1251;
  wire [(5'h11):(1'h0)] wire1479;
  reg [(4'ha):(1'h0)] reg1478 = (1'h0);
  reg [(3'h4):(1'h0)] reg1477 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1476 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1475 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1474 = (1'h0);
  reg [(5'h15):(1'h0)] reg1473 = (1'h0);
  wire signed [(5'h1a):(1'h0)] wire1472;
  reg [(5'h12):(1'h0)] reg1471 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1470 = (1'h0);
  reg [(5'h13):(1'h0)] reg1469 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1468 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1467 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1466 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1465 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1464 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1463 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1462 = (1'h0);
  reg [(4'ha):(1'h0)] reg1461 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1460 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1459 = (1'h0);
  reg [(2'h2):(1'h0)] reg1458 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1457 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1456 = (1'h0);
  reg [(4'h8):(1'h0)] reg1455 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1454 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1453 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1452 = (1'h0);
  reg [(5'h18):(1'h0)] reg1451 = (1'h0);
  reg [(5'h18):(1'h0)] reg1450 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1449 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1448 = (1'h0);
  reg [(4'h8):(1'h0)] reg1447 = (1'h0);
  reg [(2'h3):(1'h0)] reg1446 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1445 = (1'h0);
  reg [(4'ha):(1'h0)] reg1444 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1443 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1442 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1441 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1440 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1439 = (1'h0);
  reg [(3'h6):(1'h0)] reg1438 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1437 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1436 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire1435;
  reg [(4'hf):(1'h0)] reg1434 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1433 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1432 = (1'h0);
  reg [(4'he):(1'h0)] reg1431 = (1'h0);
  reg [(5'h19):(1'h0)] reg1430 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1429 = (1'h0);
  reg [(5'h18):(1'h0)] reg1428 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1427 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1426 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1425 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1424 = (1'h0);
  reg [(4'h9):(1'h0)] reg1423 = (1'h0);
  reg [(4'h8):(1'h0)] reg1422 = (1'h0);
  reg [(3'h4):(1'h0)] reg1421 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1420 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1419 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1418 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1417 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1416 = (1'h0);
  reg [(5'h15):(1'h0)] reg1415 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1414 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1413 = (1'h0);
  reg [(5'h17):(1'h0)] reg1412 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1411 = (1'h0);
  reg [(4'hb):(1'h0)] reg1410 = (1'h0);
  reg [(5'h17):(1'h0)] reg1409 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1408 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1407 = (1'h0);
  reg [(4'h9):(1'h0)] reg1406 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1405 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1404 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1403 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1402 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1401 = (1'h0);
  reg [(5'h16):(1'h0)] reg1400 = (1'h0);
  reg [(5'h17):(1'h0)] reg1399 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1398 = (1'h0);
  reg [(5'h13):(1'h0)] reg1397 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1396 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1395 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1394 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1393 = (1'h0);
  reg [(4'he):(1'h0)] reg1392 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1391 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1390 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1389 = (1'h0);
  reg [(3'h7):(1'h0)] reg1388 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1387 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1386 = (1'h0);
  wire [(5'h11):(1'h0)] wire1385;
  reg signed [(4'h8):(1'h0)] reg1384 = (1'h0);
  reg [(4'h8):(1'h0)] reg1383 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1382 = (1'h0);
  reg [(4'hb):(1'h0)] reg1381 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1380 = (1'h0);
  reg [(4'hc):(1'h0)] reg1379 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1378 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1377 = (1'h0);
  reg [(5'h19):(1'h0)] reg1376 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1375 = (1'h0);
  reg [(4'hd):(1'h0)] reg1374 = (1'h0);
  reg [(4'h9):(1'h0)] reg1373 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1372 = (1'h0);
  reg [(5'h14):(1'h0)] reg1371 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1370 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1369 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1368 = (1'h0);
  reg [(5'h14):(1'h0)] reg1367 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1366 = (1'h0);
  reg [(4'ha):(1'h0)] reg1365 = (1'h0);
  reg [(3'h4):(1'h0)] reg1364 = (1'h0);
  reg [(4'hf):(1'h0)] reg1363 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1362 = (1'h0);
  reg [(5'h12):(1'h0)] reg1361 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1360 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1359 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1358 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1357 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1356 = (1'h0);
  reg [(4'hd):(1'h0)] reg1355 = (1'h0);
  reg [(3'h6):(1'h0)] reg1354 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1353 = (1'h0);
  reg [(5'h13):(1'h0)] reg1352 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1351 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1350 = (1'h0);
  reg [(2'h3):(1'h0)] reg1349 = (1'h0);
  reg [(4'hf):(1'h0)] reg1348 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1347 = (1'h0);
  reg [(5'h18):(1'h0)] reg1346 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1345 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1344 = (1'h0);
  reg [(2'h3):(1'h0)] reg1343 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1342 = (1'h0);
  reg [(4'he):(1'h0)] reg1341 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1340 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1339 = (1'h0);
  reg [(3'h4):(1'h0)] reg1338 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1337 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1336 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1335 = (1'h0);
  reg [(5'h19):(1'h0)] reg1334 = (1'h0);
  reg [(5'h10):(1'h0)] reg1333 = (1'h0);
  reg [(4'he):(1'h0)] reg1332 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1331 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1330 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1329 = (1'h0);
  reg [(5'h10):(1'h0)] reg1328 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1327 = (1'h0);
  reg [(4'hd):(1'h0)] reg1326 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1325 = (1'h0);
  reg [(5'h16):(1'h0)] reg1324 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1323 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1322 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1321 = (1'h0);
  reg [(3'h6):(1'h0)] reg1320 = (1'h0);
  reg [(5'h17):(1'h0)] reg1319 = (1'h0);
  reg [(4'h9):(1'h0)] reg1318 = (1'h0);
  reg [(5'h14):(1'h0)] reg1317 = (1'h0);
  reg [(5'h19):(1'h0)] reg1316 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire1315;
  reg signed [(4'h9):(1'h0)] reg1314 = (1'h0);
  reg [(4'hd):(1'h0)] reg1313 = (1'h0);
  reg [(5'h14):(1'h0)] reg1312 = (1'h0);
  reg [(4'h8):(1'h0)] reg1311 = (1'h0);
  reg [(4'ha):(1'h0)] reg1310 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1309 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1308 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1307 = (1'h0);
  reg [(4'h9):(1'h0)] reg1306 = (1'h0);
  reg [(4'hd):(1'h0)] reg1305 = (1'h0);
  reg [(5'h12):(1'h0)] reg1304 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1303 = (1'h0);
  reg [(3'h4):(1'h0)] reg1302 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1301 = (1'h0);
  reg [(5'h15):(1'h0)] reg1300 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1299 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1298 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1297 = (1'h0);
  reg [(4'h8):(1'h0)] reg1296 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1295 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1294 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1293 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1292 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1291 = (1'h0);
  reg [(5'h12):(1'h0)] reg1290 = (1'h0);
  reg [(5'h15):(1'h0)] reg1289 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1288 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1287 = (1'h0);
  reg [(5'h13):(1'h0)] reg1286 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1285 = (1'h0);
  reg [(4'h9):(1'h0)] reg1284 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1283 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1282 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1281 = (1'h0);
  reg [(3'h6):(1'h0)] reg1280 = (1'h0);
  reg [(4'ha):(1'h0)] reg1279 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1278 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1277 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1276 = (1'h0);
  reg [(4'hc):(1'h0)] reg1275 = (1'h0);
  reg [(4'hc):(1'h0)] reg1274 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1273 = (1'h0);
  reg [(3'h7):(1'h0)] reg1272 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1271 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1270 = (1'h0);
  reg [(5'h13):(1'h0)] reg1269 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1268 = (1'h0);
  reg [(5'h11):(1'h0)] reg1267 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1266 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1265 = (1'h0);
  reg [(3'h6):(1'h0)] reg1264 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1263 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1262 = (1'h0);
  reg [(4'hb):(1'h0)] reg1261 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1260 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1259 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1258 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1257 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1256 = (1'h0);
  wire signed [(5'h18):(1'h0)] wire1255;
  assign y = {wire1479,
                 reg1478,
                 reg1477,
                 reg1476,
                 reg1475,
                 reg1474,
                 reg1473,
                 wire1472,
                 reg1471,
                 reg1470,
                 reg1469,
                 reg1468,
                 reg1467,
                 reg1466,
                 reg1465,
                 reg1464,
                 reg1463,
                 forvar1462,
                 reg1461,
                 forvar1460,
                 reg1459,
                 reg1458,
                 forvar1457,
                 reg1456,
                 reg1455,
                 reg1454,
                 reg1453,
                 forvar1452,
                 reg1451,
                 reg1450,
                 reg1449,
                 reg1448,
                 reg1447,
                 reg1446,
                 reg1445,
                 reg1444,
                 forvar1443,
                 reg1442,
                 reg1441,
                 reg1440,
                 forvar1439,
                 reg1438,
                 forvar1437,
                 forvar1436,
                 wire1435,
                 reg1434,
                 reg1433,
                 reg1432,
                 reg1431,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1427,
                 forvar1426,
                 reg1425,
                 reg1424,
                 reg1423,
                 reg1422,
                 reg1421,
                 forvar1420,
                 reg1419,
                 reg1418,
                 reg1417,
                 forvar1416,
                 reg1415,
                 reg1414,
                 reg1413,
                 reg1412,
                 reg1411,
                 reg1410,
                 reg1409,
                 reg1408,
                 forvar1407,
                 reg1406,
                 forvar1405,
                 reg1404,
                 reg1403,
                 reg1402,
                 reg1401,
                 reg1400,
                 reg1399,
                 forvar1398,
                 reg1397,
                 reg1396,
                 reg1395,
                 forvar1394,
                 reg1393,
                 reg1392,
                 reg1391,
                 forvar1390,
                 forvar1389,
                 reg1388,
                 reg1387,
                 forvar1386,
                 wire1385,
                 reg1384,
                 reg1383,
                 reg1382,
                 reg1381,
                 reg1380,
                 reg1379,
                 forvar1378,
                 reg1377,
                 reg1376,
                 forvar1375,
                 reg1374,
                 reg1373,
                 forvar1372,
                 reg1371,
                 reg1370,
                 reg1369,
                 reg1368,
                 reg1367,
                 reg1366,
                 reg1365,
                 reg1364,
                 reg1363,
                 reg1362,
                 reg1361,
                 reg1360,
                 reg1359,
                 forvar1358,
                 forvar1357,
                 forvar1356,
                 reg1355,
                 reg1354,
                 reg1353,
                 reg1352,
                 reg1351,
                 reg1350,
                 reg1349,
                 reg1348,
                 forvar1347,
                 reg1346,
                 reg1345,
                 forvar1344,
                 reg1343,
                 reg1342,
                 reg1341,
                 reg1340,
                 forvar1339,
                 reg1338,
                 forvar1337,
                 forvar1336,
                 reg1335,
                 reg1334,
                 reg1333,
                 reg1332,
                 forvar1331,
                 reg1330,
                 reg1329,
                 reg1328,
                 reg1327,
                 reg1326,
                 forvar1325,
                 reg1324,
                 reg1323,
                 forvar1322,
                 reg1321,
                 reg1320,
                 reg1319,
                 reg1318,
                 reg1317,
                 reg1316,
                 wire1315,
                 reg1314,
                 reg1313,
                 reg1312,
                 reg1311,
                 reg1310,
                 forvar1309,
                 reg1308,
                 reg1307,
                 reg1306,
                 reg1305,
                 reg1304,
                 forvar1303,
                 reg1302,
                 reg1301,
                 reg1300,
                 reg1299,
                 reg1298,
                 reg1297,
                 reg1296,
                 reg1295,
                 forvar1294,
                 reg1293,
                 forvar1292,
                 reg1291,
                 reg1290,
                 reg1289,
                 reg1288,
                 reg1287,
                 reg1286,
                 reg1285,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1281,
                 reg1280,
                 reg1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 reg1275,
                 reg1274,
                 reg1273,
                 reg1272,
                 reg1271,
                 forvar1270,
                 reg1269,
                 reg1268,
                 reg1267,
                 forvar1266,
                 reg1265,
                 reg1264,
                 reg1263,
                 reg1262,
                 reg1261,
                 reg1260,
                 reg1259,
                 forvar1258,
                 reg1257,
                 reg1256,
                 wire1255,
                 (1'h0)};
  assign wire1255 = (~|$unsigned((8'ha9)));
  always
    @(posedge clk) begin
      reg1256 <= $signed(($unsigned(wire1251) ?
          $signed(({wire1252,
              wire1253} - $signed(wire1251))) : wire1254[(1'h1):(1'h0)]));
      reg1257 <= (wire1254[(4'h8):(2'h2)] ?
          $unsigned($unsigned((^wire1253))) : {"ivLk",
              $signed(((wire1254 ?
                  (7'h48) : wire1254) + reg1256[(3'h6):(2'h3)]))});
      for (forvar1258 = (1'h0); (forvar1258 < (1'h0)); forvar1258 = (forvar1258 + (1'h1)))
        begin
          reg1259 <= "vwVyMAhbXNOFoCM41seRv";
          reg1260 <= ("GCcWfrxGJ5NK9AL" ?
              (&(|wire1253[(5'h13):(5'h13)])) : (($unsigned((8'haf)) ?
                      (+(&wire1253)) : $signed((wire1251 ?
                          reg1257 : (8'hb7)))) ?
                  reg1257 : $unsigned(reg1259)));
        end
      reg1261 <= $unsigned(($signed(((wire1251 ?
          wire1251 : reg1259) << (reg1256 ?
          wire1253 : reg1260))) < $signed("xHsIs")));
      reg1262 <= reg1257[(4'hb):(3'h7)];
      reg1263 <= (({{"9cYLWermxZl5O6fALX5Td7g"}, reg1262} ?
          wire1252[(4'hc):(4'h9)] : "pwK0UUWiCwFt7fx") >> (^~(8'h9d)));
    end
  always
    @(posedge clk) begin
      reg1264 <= reg1262;
      reg1265 <= $unsigned($unsigned((!wire1254)));
      for (forvar1266 = (1'h0); (forvar1266 < (3'h4)); forvar1266 = (forvar1266 + (1'h1)))
        begin
          reg1267 <= (~&(forvar1258[(3'h7):(2'h2)] ?
              $unsigned("vLHGBQ6h1ZQoyU20I") : (~&$unsigned({reg1264}))));
          reg1268 <= wire1252;
          reg1269 = (!$unsigned($signed((^$unsigned(reg1267)))));
          for (forvar1270 = (1'h0); (forvar1270 < (1'h1)); forvar1270 = (forvar1270 + (1'h1)))
            begin
              reg1271 <= {"SBg3e2gpZ8v"};
              reg1272 <= ($signed("sBeK6AUp") ?
                  (("nPILc" <<< ({wire1251,
                      reg1265} & reg1264)) >>> (($unsigned(wire1253) ?
                          (wire1252 || (8'hac)) : (forvar1270 < wire1255)) ?
                      "PEvVNMQWITqIIXyTqf4NqMO" : reg1269)) : $unsigned(reg1265));
            end
          reg1273 <= {"buZ2EmVa", $unsigned(("LZvD0" <<< $signed(reg1264)))};
          reg1274 <= "II61";
        end
      reg1275 <= (-(forvar1258[(3'h6):(1'h0)] >>> $unsigned(("nsfQ" + reg1265))));
      reg1276 = (forvar1270 >> "8cyAfwyyrEzOqPLF");
      reg1277 <= "sG5Ip3lAegX";
    end
  always
    @(posedge clk) begin
      reg1278 <= $unsigned($signed(reg1275));
      reg1279 = reg1273[(3'h4):(2'h3)];
      reg1280 <= $signed("zE5o8ehfXswP53");
      reg1281 = $signed((&reg1278[(3'h7):(1'h0)]));
      reg1282 = (~^$signed(reg1260));
      reg1283 <= ((reg1275 ?
          $unsigned((&$unsigned(reg1274))) : $signed(((~reg1274) ?
              $unsigned((8'hac)) : $unsigned(reg1278)))) ^ $unsigned(((~&reg1276[(5'h13):(4'hb)]) ?
          ($signed(reg1273) > $unsigned((7'h42))) : $unsigned(reg1260[(5'h14):(1'h0)]))));
    end
  always
    @(posedge clk) begin
      reg1284 <= $unsigned("2k6U");
      reg1285 <= (!(($unsigned($signed(reg1267)) ?
          (reg1259[(5'h11):(1'h0)] ?
              "aPmHU3k5zPLzsXUkiQ2Ea6" : (reg1268 ?
                  reg1284 : forvar1270)) : $unsigned("a1sBk9Nod2TA8Y")) == "Dfr"));
      reg1286 <= (^~$unsigned((7'h47)));
      reg1287 <= $signed($signed(reg1286[(4'hf):(4'hf)]));
    end
  always
    @(posedge clk) begin
      reg1288 = "hxZ";
      reg1289 <= ($signed((7'h4a)) != (~({$unsigned(reg1283),
          "gy1UeEf7"} > "qIKyQqfD3BYir")));
      reg1290 <= "zR5Gl3kDaCk";
      reg1291 <= $unsigned((($signed($signed(reg1274)) && ((reg1259 * reg1277) - $unsigned((7'h43)))) * $signed($signed(reg1279[(3'h7):(3'h6)]))));
      for (forvar1292 = (1'h0); (forvar1292 < (2'h3)); forvar1292 = (forvar1292 + (1'h1)))
        begin
          reg1293 <= "wNyDRM2lycihQD0LAR";
        end
    end
  always
    @(posedge clk) begin
      for (forvar1294 = (1'h0); (forvar1294 < (2'h2)); forvar1294 = (forvar1294 + (1'h1)))
        begin
          reg1295 <= (&$unsigned((~|($unsigned(reg1291) ?
              $signed(reg1271) : (reg1267 ? (8'ha5) : reg1257)))));
          reg1296 = (("0DeTWmxfR9" ^~ reg1293) ? reg1279 : reg1293);
          reg1297 = $unsigned(reg1274[(1'h1):(1'h1)]);
          reg1298 <= (~|$unsigned({((reg1273 << reg1273) ?
                  (forvar1292 ?
                      reg1297 : reg1281) : wire1252[(4'hf):(1'h1)])}));
        end
      reg1299 <= (+$unsigned(reg1296[(3'h7):(1'h1)]));
      reg1300 <= ($unsigned("6V9nCBsDcUpsZMh3t8p7") * (($unsigned({reg1299}) ?
              ($signed((8'hbd)) ?
                  reg1285 : (-reg1259)) : "zlBqr4e9FotW4hsxGJ") ?
          reg1290[(4'h8):(4'h8)] : ({{reg1260, reg1286},
              (reg1282 && reg1282)} ^~ $unsigned(reg1291[(2'h2):(1'h1)]))));
      reg1301 <= (8'hab);
      reg1302 = reg1300[(5'h15):(5'h14)];
    end
  always
    @(posedge clk) begin
      for (forvar1303 = (1'h0); (forvar1303 < (3'h4)); forvar1303 = (forvar1303 + (1'h1)))
        begin
          reg1304 <= ((&"RtoHrSy5nDFnLhnLqKosZrP") << ((^{$unsigned((8'ha7))}) >= $signed((!forvar1266[(5'h10):(4'he)]))));
          reg1305 <= (($unsigned(reg1286) && $signed(((reg1287 <<< (8'h9c)) ?
              ((8'ha5) ?
                  reg1265 : reg1261) : $unsigned(reg1297)))) >= $signed("IWy13Ez3rcun5l0PmYcm6yt"));
          reg1306 <= (("n" ?
              $unsigned($signed("WMNKMCUdCG3K")) : {((reg1300 ?
                      (8'had) : reg1281) != $unsigned((8'ha0))),
                  reg1293}) - (^$unsigned($signed("BIv1f25IG"))));
        end
      reg1307 <= $signed((8'hba));
      reg1308 <= ((($signed($unsigned(reg1256)) ?
              reg1282 : reg1256) ^~ (~^reg1272)) ?
          $unsigned({"3GFdUA3JJsWVhudTS3"}) : reg1283);
      for (forvar1309 = (1'h0); (forvar1309 < (1'h0)); forvar1309 = (forvar1309 + (1'h1)))
        begin
          reg1310 <= ({reg1262[(1'h1):(1'h0)]} <= ((^$signed((^reg1271))) == ({(reg1288 <= (8'hb4))} ?
              reg1300 : wire1253)));
          reg1311 <= $unsigned(reg1265);
          reg1312 <= $signed(wire1254[(4'he):(3'h7)]);
          reg1313 <= $unsigned(($unsigned((reg1265[(2'h3):(2'h3)] ?
                  $unsigned((7'h47)) : {reg1278, reg1296})) ?
              "TLQhZY" : "a5VlRL4TDoIOEZDm7bD2HRXAb"));
        end
      reg1314 <= ("vZfUqWmJl3Rowl7LBiaa" <= (^(((reg1293 ?
          reg1279 : forvar1292) > ((8'ha3) ?
          reg1312 : reg1312)) && (^$signed((8'had))))));
    end
  assign wire1315 = $unsigned(reg1305);
  always
    @(posedge clk) begin
      reg1316 = $unsigned((wire1255[(2'h3):(1'h1)] ?
          reg1281[(4'h9):(4'h8)] : (~&(!wire1252[(3'h4):(2'h3)]))));
      reg1317 <= forvar1258[(1'h0):(1'h0)];
      reg1318 <= ((8'ha9) ?
          {reg1284[(3'h6):(3'h4)],
              (~((&reg1286) ?
                  ((7'h43) ? reg1261 : wire1254) : (8'h9c)))} : (+reg1272));
      reg1319 = ((^~reg1269) ?
          ($unsigned($signed(((7'h4d) | forvar1258))) ?
              reg1302 : ($signed($signed(reg1296)) <= (((7'h45) <= reg1259) <<< $signed(reg1282)))) : "Oiq6hs2Ym5FgSoX");
      reg1320 <= reg1313;
      reg1321 = "qTxGl0Lr";
    end
  always
    @(posedge clk) begin
      for (forvar1322 = (1'h0); (forvar1322 < (2'h3)); forvar1322 = (forvar1322 + (1'h1)))
        begin
          reg1323 <= $unsigned($unsigned($unsigned($unsigned($signed(reg1312)))));
          reg1324 = forvar1303;
          for (forvar1325 = (1'h0); (forvar1325 < (2'h2)); forvar1325 = (forvar1325 + (1'h1)))
            begin
              reg1326 <= (reg1277 ?
                  ("z6T" ?
                      "vKNgFPlY3CGolwtaY" : $signed($unsigned(reg1264))) : "2QYF5OoXwWXNYaZCOsL7ivfs");
              reg1327 = ($signed(($unsigned((^reg1295)) & ({reg1256} ?
                  reg1265[(4'h8):(3'h5)] : $unsigned(forvar1270)))) - $unsigned($unsigned({(forvar1322 ?
                      reg1323 : reg1297),
                  reg1280[(1'h1):(1'h0)]})));
              reg1328 <= {(~((~^$unsigned((7'h40))) ?
                      {forvar1325, {reg1259}} : ((reg1301 <<< (8'ha0)) ?
                          {reg1296} : (reg1321 != (8'hb6))))),
                  reg1327[(5'h10):(4'h9)]};
              reg1329 <= $signed(($signed(reg1308) == ((wire1254 || (~&(8'ha7))) ?
                  "Mg4gyb7Qnpfxsm9NO90JeQ" : ("1fNeXgG3o1SbFBQ1sb" ~^ $unsigned(reg1310)))));
              reg1330 <= wire1252;
              for (forvar1331 = (1'h0); (forvar1331 < (2'h2)); forvar1331 = (forvar1331 + (1'h1)))
                begin
                  reg1332 <= ((7'h43) != (reg1310 ?
                      (reg1307 ? "vo49cmIZnU4m" : (^~(-(8'hb9)))) : reg1307));
                  reg1333 <= $unsigned((+("AmfwI9VvzOLodHnhqe" ?
                      $unsigned({reg1319, reg1271}) : ($signed(reg1308) ?
                          (!reg1310) : {(8'hac)}))));
                end
            end
        end
      reg1334 <= (~&$unsigned(($unsigned((reg1332 + wire1254)) - reg1330)));
    end
  always
    @(posedge clk) begin
      reg1335 <= reg1286[(3'h6):(2'h2)];
      for (forvar1336 = (1'h0); (forvar1336 < (3'h5)); forvar1336 = (forvar1336 + (1'h1)))
        begin
          for (forvar1337 = (1'h0); (forvar1337 < (3'h5)); forvar1337 = (forvar1337 + (1'h1)))
            begin
              reg1338 <= $signed({reg1282[(4'hc):(3'h6)]});
              for (forvar1339 = (1'h0); (forvar1339 < (1'h1)); forvar1339 = (forvar1339 + (1'h1)))
                begin
                  reg1340 = $signed(reg1281[(5'h10):(1'h1)]);
                end
              reg1341 <= ("799uFGFYxBc1DI" ?
                  (+$signed(($signed(reg1268) ?
                      (reg1304 ?
                          wire1253 : reg1340) : (^forvar1339)))) : reg1304);
              reg1342 <= (~&((+"cLLHEhN3BXLy9wV1Q5JW2") > ((^~reg1295[(1'h0):(1'h0)]) ?
                  reg1317 : reg1256)));
              reg1343 <= (~{"7K1c3z4Yas5t0agq", $signed(reg1291)});
            end
          for (forvar1344 = (1'h0); (forvar1344 < (2'h2)); forvar1344 = (forvar1344 + (1'h1)))
            begin
              reg1345 <= forvar1309;
              reg1346 <= "ku304skqsNv";
              for (forvar1347 = (1'h0); (forvar1347 < (3'h4)); forvar1347 = (forvar1347 + (1'h1)))
                begin
                  reg1348 <= "hxA3X2uUBACZzlTeBmuiM2";
                  reg1349 <= reg1346;
                end
            end
          reg1350 <= {(+$signed({(reg1296 ? reg1264 : reg1289),
                  (reg1300 != (8'h9d))}))};
        end
      reg1351 = (reg1332[(3'h6):(1'h0)] ?
          $signed((($signed(reg1341) <<< $signed(reg1343)) ?
              ($unsigned(forvar1322) | {reg1314, reg1280}) : ((reg1274 ?
                  (8'hbf) : (8'hb9)) ~^ $unsigned(reg1313)))) : wire1254[(4'hd):(1'h0)]);
      reg1352 <= (|wire1253);
    end
  always
    @(posedge clk) begin
      reg1353 = (7'h46);
      reg1354 = ($signed($signed($signed((reg1304 ~^ reg1352)))) ?
          ("X3ir" + $signed($unsigned({(8'hbc)}))) : $signed({(~reg1297)}));
      reg1355 <= (~reg1345[(3'h5):(1'h1)]);
    end
  always
    @(posedge clk) begin
      for (forvar1356 = (1'h0); (forvar1356 < (1'h1)); forvar1356 = (forvar1356 + (1'h1)))
        begin
          for (forvar1357 = (1'h0); (forvar1357 < (2'h3)); forvar1357 = (forvar1357 + (1'h1)))
            begin
              for (forvar1358 = (1'h0); (forvar1358 < (1'h0)); forvar1358 = (forvar1358 + (1'h1)))
                begin
                  reg1359 <= "ZwbuvSQiSCR6YMuGbk";
                  reg1360 <= "VsBosU";
                  reg1361 <= ($unsigned("8JbWvzaQRgONr1VEnqyoUWHyA") ?
                      reg1293 : ((reg1290 ?
                          (reg1284[(4'h8):(4'h8)] & "nVE") : reg1291) && (forvar1344 ?
                          (reg1334 ^~ (~&(7'h49))) : $signed({reg1260}))));
                  reg1362 <= reg1300;
                  reg1363 <= reg1262;
                  reg1364 <= (~^reg1340[(4'he):(1'h1)]);
                end
              reg1365 <= (~&((-(^forvar1331)) >> ("4D4LZLOO" ?
                  reg1338 : $unsigned(reg1262))));
              reg1366 = reg1338[(1'h1):(1'h1)];
              reg1367 <= ($unsigned("UEychbHuHru6ieDGKxqYTx") ?
                  "5KXTFmmsOtJYtc" : {$unsigned((^reg1311[(3'h5):(1'h1)]))});
              reg1368 <= $signed($signed(((+"yDn") ? (8'hab) : forvar1266)));
            end
          reg1369 <= (+(8'hab));
          reg1370 <= reg1295[(3'h4):(2'h2)];
          reg1371 <= (8'ha7);
        end
      for (forvar1372 = (1'h0); (forvar1372 < (2'h2)); forvar1372 = (forvar1372 + (1'h1)))
        begin
          reg1373 <= (8'hae);
          reg1374 <= (forvar1292 ? forvar1331[(5'h10):(1'h0)] : "J1JwntWghOyI");
          for (forvar1375 = (1'h0); (forvar1375 < (1'h1)); forvar1375 = (forvar1375 + (1'h1)))
            begin
              reg1376 <= "OuWOsaaS4HQbv";
              reg1377 <= $unsigned(reg1316);
              for (forvar1378 = (1'h0); (forvar1378 < (2'h3)); forvar1378 = (forvar1378 + (1'h1)))
                begin
                  reg1379 = reg1278[(3'h7):(3'h5)];
                  reg1380 <= $signed(($signed((reg1340 ?
                      (|forvar1258) : (~|wire1252))) >>> $unsigned("lYz5H")));
                  reg1381 <= (~^reg1297);
                  reg1382 <= "yaVncuwKOlnuvYFgGuyKM7";
                end
              reg1383 <= (|$signed($signed(($unsigned((8'hb4)) ?
                  (reg1312 ? (8'ha1) : reg1305) : "oKW2KD29IHcP8b"))));
              reg1384 <= reg1304;
            end
        end
    end
  assign wire1385 = (~{"bTz9gH473ExTUvbl7EKgKV",
                        $unsigned((reg1285 ?
                            (^~reg1257) : (reg1316 * reg1276)))});
  always
    @(posedge clk) begin
      for (forvar1386 = (1'h0); (forvar1386 < (2'h2)); forvar1386 = (forvar1386 + (1'h1)))
        begin
          reg1387 = {(($unsigned(reg1313[(2'h3):(2'h2)]) ?
                      ((forvar1322 == reg1308) ?
                          reg1306[(3'h7):(1'h1)] : $unsigned(reg1288)) : (~|(~^reg1261))) ?
                  (+$signed($unsigned(reg1341))) : reg1348[(4'h9):(3'h7)])};
          reg1388 <= ((reg1286 ^ {reg1354[(3'h5):(1'h0)]}) == reg1376);
          for (forvar1389 = (1'h0); (forvar1389 < (1'h1)); forvar1389 = (forvar1389 + (1'h1)))
            begin
              for (forvar1390 = (1'h0); (forvar1390 < (3'h5)); forvar1390 = (forvar1390 + (1'h1)))
                begin
                  reg1391 <= {($signed(((-forvar1390) < (!reg1374))) ?
                          (7'h49) : "HGgb7qtThSFSNyDmXx7oo2p")};
                  reg1392 <= (^~"AfU7NKwuHTYatk");
                  reg1393 <= ((!reg1345) >>> ((reg1296[(3'h7):(3'h4)] ?
                      reg1329[(4'hb):(1'h1)] : (8'hbf)) == reg1272[(1'h1):(1'h0)]));
                end
              for (forvar1394 = (1'h0); (forvar1394 < (3'h5)); forvar1394 = (forvar1394 + (1'h1)))
                begin
                  reg1395 <= (reg1371[(1'h1):(1'h0)] ?
                      forvar1258[(3'h4):(2'h3)] : forvar1347[(3'h6):(3'h6)]);
                  reg1396 = $signed((("FivcxRdpRw0KTvpt9p" ?
                      $unsigned(reg1327[(4'he):(3'h5)]) : {$unsigned((7'h42)),
                          "BdTX7GNHi"}) << $signed(forvar1389)));
                  reg1397 <= $signed(((("" ?
                      {(8'hbb),
                          reg1330} : $signed(forvar1394)) >= $signed((reg1363 | reg1340))) ^ $unsigned($signed("eKTmmssUh8Hs7"))));
                end
            end
          for (forvar1398 = (1'h0); (forvar1398 < (3'h5)); forvar1398 = (forvar1398 + (1'h1)))
            begin
              reg1399 <= (reg1256[(4'h8):(2'h2)] ? $signed((8'ha3)) : wire1253);
            end
          reg1400 <= (forvar1394[(1'h1):(1'h1)] ?
              forvar1266[(5'h11):(4'hf)] : (^~reg1265[(2'h2):(1'h1)]));
        end
    end
  always
    @(posedge clk) begin
      reg1401 <= $signed(reg1272[(1'h0):(1'h0)]);
      reg1402 <= ($unsigned(reg1352) ?
          reg1329[(5'h14):(4'ha)] : reg1392[(4'h8):(3'h5)]);
      reg1403 <= $unsigned($signed(({$unsigned(reg1379),
              "T8UBuzZkGRTdfeSavOpwC2qhk"} ?
          ("f8scAsw5CyI4bQvNEluGqD1S" < (~&reg1299)) : {(~reg1323),
              $signed(reg1361)})));
      reg1404 <= ("lJnJrw5k2SbA0iH4Lw" ?
          ($unsigned(((~|reg1333) ?
              ((8'ha8) ?
                  reg1320 : reg1289) : reg1360[(4'hd):(4'ha)])) == forvar1270[(2'h2):(1'h0)]) : "9Op");
      for (forvar1405 = (1'h0); (forvar1405 < (3'h4)); forvar1405 = (forvar1405 + (1'h1)))
        begin
          reg1406 <= (|{{("xCBqV44hz" ?
                      (forvar1292 && forvar1266) : (forvar1294 ?
                          forvar1389 : reg1312)),
                  reg1402[(5'h15):(3'h6)]},
              "Nbh1oJ8HIzrvn183"});
        end
      for (forvar1407 = (1'h0); (forvar1407 < (3'h5)); forvar1407 = (forvar1407 + (1'h1)))
        begin
          reg1408 = reg1342;
          reg1409 <= {((^(&$unsigned(reg1374))) <= reg1399[(3'h4):(2'h2)])};
          reg1410 <= (|reg1301[(2'h2):(1'h0)]);
          reg1411 <= ((^"Z") >> reg1285);
          reg1412 = wire1252;
        end
    end
  always
    @(posedge clk) begin
      reg1413 <= "cL4U2NF";
      reg1414 <= (8'ha7);
      reg1415 = (!(!reg1280[(3'h6):(1'h1)]));
      for (forvar1416 = (1'h0); (forvar1416 < (1'h0)); forvar1416 = (forvar1416 + (1'h1)))
        begin
          reg1417 <= {$unsigned((({(7'h42), reg1410} ?
                  $signed((8'hbb)) : $signed(forvar1292)) ^~ forvar1294))};
          reg1418 = reg1313[(1'h1):(1'h0)];
          reg1419 = forvar1358;
          for (forvar1420 = (1'h0); (forvar1420 < (3'h4)); forvar1420 = (forvar1420 + (1'h1)))
            begin
              reg1421 <= $unsigned(((~reg1318) ?
                  {(^~"vRFHWES06kZCPMVmg14GyS")} : ($unsigned($unsigned(reg1310)) ?
                      ($unsigned(reg1296) ?
                          (reg1318 && reg1256) : (reg1369 ~^ reg1363)) : reg1396)));
              reg1422 <= (!$signed("pzn6Rwl8A6AD7zXr"));
              reg1423 <= $unsigned((~forvar1358));
              reg1424 <= reg1289[(1'h0):(1'h0)];
              reg1425 <= forvar1390[(2'h3):(2'h3)];
              for (forvar1426 = (1'h0); (forvar1426 < (3'h4)); forvar1426 = (forvar1426 + (1'h1)))
                begin
                  reg1427 <= (+forvar1426[(3'h5):(1'h1)]);
                  reg1428 <= $unsigned(("mos0" ?
                      (($unsigned(forvar1336) ?
                          forvar1303[(3'h5):(1'h1)] : (~&reg1361)) != ($signed(reg1381) >> reg1417)) : "pX9PnO2vc6MVIBbO3"));
                  reg1429 = reg1307[(4'h9):(2'h3)];
                  reg1430 <= (8'hb6);
                  reg1431 <= (&reg1334);
                end
            end
          reg1432 <= $unsigned(reg1297[(1'h0):(1'h0)]);
        end
    end
  always
    @(posedge clk) begin
      reg1433 <= reg1380[(1'h0):(1'h0)];
      reg1434 <= reg1259[(3'h4):(3'h4)];
    end
  assign wire1435 = (!$signed({$signed((reg1340 ? forvar1322 : reg1329))}));
  always
    @(posedge clk) begin
      for (forvar1436 = (1'h0); (forvar1436 < (1'h1)); forvar1436 = (forvar1436 + (1'h1)))
        begin
          for (forvar1437 = (1'h0); (forvar1437 < (2'h2)); forvar1437 = (forvar1437 + (1'h1)))
            begin
              reg1438 = $signed(reg1300[(1'h1):(1'h0)]);
            end
          for (forvar1439 = (1'h0); (forvar1439 < (3'h4)); forvar1439 = (forvar1439 + (1'h1)))
            begin
              reg1440 <= (($unsigned($signed("7da5eRbuTz635UREPEzf")) ?
                      (reg1349[(2'h3):(1'h1)] ?
                          reg1256 : (reg1404[(4'hd):(2'h3)] <= $unsigned(wire1252))) : "I8W1e12cMpBktNcUkIl") ?
                  "Um" : forvar1270[(3'h7):(2'h3)]);
              reg1441 <= "qYDJW8CYT0TnNoBQyy";
            end
        end
      reg1442 <= forvar1331;
      for (forvar1443 = (1'h0); (forvar1443 < (3'h4)); forvar1443 = (forvar1443 + (1'h1)))
        begin
          reg1444 <= (reg1296[(2'h3):(1'h0)] ^~ "Iix");
          reg1445 <= reg1257;
          reg1446 <= reg1256;
          reg1447 <= $unsigned($signed(($signed((8'hb4)) || {forvar1394,
              reg1335[(3'h5):(1'h0)]})));
          reg1448 <= ((~^($unsigned((&reg1396)) <<< $signed($unsigned(reg1441)))) && (+reg1400[(2'h3):(2'h2)]));
        end
    end
  always
    @(posedge clk) begin
      reg1449 <= reg1291;
      reg1450 <= "BC6OzbEs0MhAKgZVJFlR";
      reg1451 = reg1302[(1'h0):(1'h0)];
      for (forvar1452 = (1'h0); (forvar1452 < (3'h5)); forvar1452 = (forvar1452 + (1'h1)))
        begin
          reg1453 <= reg1293;
          reg1454 = "1HE7HgyqH";
          reg1455 <= $signed((-{((reg1442 <= reg1319) != (~^(8'hb8)))}));
          reg1456 <= (forvar1437[(5'h11):(3'h7)] ?
              (&reg1271) : (~(~$unsigned(reg1421))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar1457 = (1'h0); (forvar1457 < (2'h2)); forvar1457 = (forvar1457 + (1'h1)))
        begin
          reg1458 <= (reg1446 ~^ (({(reg1327 ? forvar1336 : reg1305),
              $unsigned(reg1275)} * ((forvar1437 ? reg1332 : reg1366) ?
              reg1273[(4'h9):(2'h3)] : reg1304)) <= (~|(reg1308[(1'h1):(1'h0)] ~^ $unsigned(reg1350)))));
          reg1459 <= {$signed({$signed((|reg1277))}),
              (("WJCgw7t" ? $signed("kEGzR5kuqew6kk") : $unsigned({reg1374})) ?
                  (|($unsigned(wire1251) != "W8IiaBo8tA")) : (reg1404[(2'h3):(2'h3)] & $signed(reg1430[(4'hb):(3'h7)])))};
          for (forvar1460 = (1'h0); (forvar1460 < (1'h0)); forvar1460 = (forvar1460 + (1'h1)))
            begin
              reg1461 <= $signed((reg1381[(3'h5):(2'h2)] ?
                  forvar1325 : reg1397[(2'h3):(2'h2)]));
              for (forvar1462 = (1'h0); (forvar1462 < (1'h0)); forvar1462 = (forvar1462 + (1'h1)))
                begin
                  reg1463 <= (reg1361 ? (8'hb3) : {(-$unsigned((+reg1444)))});
                  reg1464 <= forvar1462[(2'h3):(1'h0)];
                  reg1465 <= (forvar1394 > "RFx6oNsJc2");
                  reg1466 = forvar1398[(1'h1):(1'h0)];
                  reg1467 <= (($unsigned($signed((reg1334 ?
                              forvar1344 : reg1295))) ?
                          (reg1465 >> (|reg1296)) : (!forvar1292)) ?
                      wire1435[(1'h0):(1'h0)] : (^(^~(reg1401[(5'h12):(4'ha)] ?
                          (reg1430 ? reg1327 : forvar1378) : (reg1271 ?
                              (8'ha7) : reg1323)))));
                end
              reg1468 <= $signed($signed({"tkz6Ztbdm29nNcEkSNydW"}));
            end
          reg1469 = $signed(((($signed(reg1293) ?
              (~^forvar1266) : (|reg1277)) == $unsigned((reg1448 * forvar1270))) * ($unsigned((reg1366 >> reg1414)) == ("0MEqztezGLzluR5Iivde" ?
              (~&reg1466) : $unsigned(reg1412)))));
          reg1470 <= $unsigned(($unsigned((~&(reg1268 ?
              reg1281 : (8'ha7)))) != ("BsIO1u7mwLbKwWEvdq" ?
              $signed(forvar1443) : ("bT69rwkre7PxG" ^~ reg1413[(1'h0):(1'h0)]))));
          reg1471 <= forvar1457;
        end
    end
  assign wire1472 = "zPWab4nPGk";
  always
    @(posedge clk) begin
      reg1473 <= $unsigned(forvar1436[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg1474 = $signed((forvar1390 ?
          ($unsigned("6ifIXIhmdvgr") <= (8'hb1)) : {$signed($unsigned(reg1271)),
              $unsigned(reg1396[(4'h9):(3'h6)])}));
      reg1475 = reg1440[(4'h8):(2'h3)];
      reg1476 = (forvar1439 ?
          reg1427[(3'h6):(2'h3)] : (("vVIfkJUBKWX0ZaRmOvgLSMa" * $signed(forvar1439)) ?
              (+(reg1393 - (-(8'hb7)))) : (((reg1312 ?
                  reg1362 : reg1384) - (~&reg1362)) < (^~reg1311))));
      reg1477 <= reg1471;
      reg1478 <= $unsigned("7");
    end
  assign wire1479 = $signed((8'hab));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1210
#( parameter param1246 = (!(7'h4e))
, parameter param1247 = ((^param1246) ? param1246 : ((param1246 ~^ (^(~param1246))) + ((7'h42) ? ((param1246 ? param1246 : param1246) ? (param1246 ^ param1246) : (8'hb3)) : param1246))) )
(y, clk, wire1214, wire1213, wire1212, wire1211);
  output wire [(32'h1b0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire1214;
  input wire [(3'h5):(1'h0)] wire1213;
  input wire [(3'h7):(1'h0)] wire1212;
  input wire signed [(5'h12):(1'h0)] wire1211;
  wire signed [(3'h5):(1'h0)] wire1245;
  reg signed [(3'h4):(1'h0)] reg1244 = (1'h0);
  reg [(4'he):(1'h0)] reg1243 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1242 = (1'h0);
  reg [(5'h17):(1'h0)] reg1241 = (1'h0);
  wire signed [(5'h16):(1'h0)] wire1240;
  wire [(3'h4):(1'h0)] wire1239;
  reg [(4'hb):(1'h0)] reg1238 = (1'h0);
  reg [(5'h10):(1'h0)] reg1237 = (1'h0);
  reg [(4'ha):(1'h0)] reg1236 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1235 = (1'h0);
  reg [(5'h10):(1'h0)] reg1234 = (1'h0);
  reg [(4'hb):(1'h0)] reg1233 = (1'h0);
  reg [(5'h14):(1'h0)] reg1232 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1231 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1230 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1229 = (1'h0);
  reg [(5'h16):(1'h0)] reg1228 = (1'h0);
  reg [(4'hc):(1'h0)] reg1227 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1226 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1225 = (1'h0);
  reg [(3'h4):(1'h0)] reg1224 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1223 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1222 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1221 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1220 = (1'h0);
  reg [(3'h6):(1'h0)] reg1219 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1218 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1217 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1216 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1215 = (1'h0);
  assign y = {wire1245,
                 reg1244,
                 reg1243,
                 reg1242,
                 reg1241,
                 wire1240,
                 wire1239,
                 reg1238,
                 reg1237,
                 reg1236,
                 reg1235,
                 reg1234,
                 reg1233,
                 reg1232,
                 reg1231,
                 reg1230,
                 forvar1229,
                 reg1228,
                 reg1227,
                 reg1226,
                 reg1225,
                 reg1224,
                 forvar1223,
                 reg1222,
                 reg1221,
                 forvar1220,
                 reg1219,
                 reg1218,
                 reg1217,
                 reg1216,
                 reg1215,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1215 <= {"Rf",
          ((+((wire1213 != wire1213) - wire1211)) ?
              "fhF14R" : ({$signed(wire1211),
                  $unsigned(wire1214)} ^ (&wire1214)))};
      reg1216 = $signed("CyaxyhhEUQxymMatwlvefGxC");
      reg1217 = wire1214[(4'h9):(1'h1)];
      reg1218 = $unsigned($unsigned(wire1212[(3'h5):(3'h5)]));
    end
  always
    @(posedge clk) begin
      reg1219 <= "h10PoWk1lmeHGTFJFLa2WnBG";
      for (forvar1220 = (1'h0); (forvar1220 < (1'h0)); forvar1220 = (forvar1220 + (1'h1)))
        begin
          reg1221 <= ((-$signed((+$signed(reg1219)))) ?
              reg1217 : (reg1216 ? forvar1220 : reg1219[(2'h2):(1'h0)]));
          reg1222 <= ($signed("Xtx1PRqkcCUk") ?
              wire1212[(1'h0):(1'h0)] : "mwkplc");
          for (forvar1223 = (1'h0); (forvar1223 < (2'h2)); forvar1223 = (forvar1223 + (1'h1)))
            begin
              reg1224 <= ("pLpKnbkcZfLFNzAxII8" ?
                  $unsigned($unsigned((-$signed(reg1215)))) : ($unsigned("2fOw7") ?
                      "" : ($unsigned((reg1219 >>> reg1221)) ?
                          "0Y" : (~^$signed((8'hae))))));
              reg1225 <= (("CLWZFcUJzKTOsRyqRGyX" < "WfLJZKYpBvhCZvBJhahMGD") ?
                  (reg1218 ?
                      $signed(((forvar1223 >> wire1212) ?
                          (reg1219 < forvar1220) : {reg1216})) : (!reg1219)) : reg1218[(2'h3):(1'h0)]);
            end
          reg1226 <= forvar1223;
          reg1227 <= ($signed(($unsigned({forvar1223, (8'hbb)}) ?
              $signed($unsigned(reg1217)) : "RLGDhyRCdznPHsb")) ^ wire1212[(3'h4):(1'h1)]);
        end
      reg1228 <= {wire1212, reg1217};
      for (forvar1229 = (1'h0); (forvar1229 < (1'h0)); forvar1229 = (forvar1229 + (1'h1)))
        begin
          reg1230 = reg1216;
          reg1231 = ((~|$unsigned($unsigned(reg1228[(3'h7):(1'h0)]))) ?
              (forvar1223 != (({wire1214} ?
                      (reg1221 + wire1211) : reg1227[(4'h9):(4'h9)]) ?
                  $unsigned({reg1218}) : $signed(reg1227[(4'h8):(3'h4)]))) : reg1222[(2'h2):(1'h0)]);
          reg1232 <= ((~(|"JnkFunyX")) ?
              $unsigned((-((!wire1213) ?
                  $unsigned(reg1226) : $unsigned(forvar1220)))) : $signed({$signed(forvar1220)}));
        end
      reg1233 <= $signed((((~&(wire1213 ? reg1215 : forvar1220)) ?
              {$signed(reg1226)} : forvar1223[(2'h3):(2'h2)]) ?
          reg1222[(2'h2):(1'h1)] : reg1221));
      reg1234 <= "7hGw84f";
    end
  always
    @(posedge clk) begin
      reg1235 <= $unsigned(reg1230[(5'h12):(4'hf)]);
      reg1236 <= {$signed($signed(("AnZcHnmSUJzJgYnKY" ^~ (reg1221 ?
              (7'h4c) : reg1219))))};
      reg1237 <= $signed("J6");
      reg1238 <= $unsigned(wire1214);
    end
  assign wire1239 = forvar1223;
  assign wire1240 = ((~&$unsigned(reg1218)) >= (($unsigned($signed(reg1228)) ?
                            ((!reg1238) >= (forvar1220 * wire1214)) : reg1219[(3'h5):(3'h4)]) ?
                        (reg1234 ?
                            ($signed(wire1211) ?
                                reg1222 : (reg1222 ?
                                    forvar1220 : reg1218)) : "r2WQDJ") : ("0cN5oQppDGE1X0JiHyw" ^ ($signed(reg1238) >>> (|forvar1223)))));
  always
    @(posedge clk) begin
      reg1241 <= $signed($unsigned(({wire1212[(1'h1):(1'h1)]} <<< reg1232[(2'h2):(2'h2)])));
      reg1242 <= $unsigned((8'ha3));
      reg1243 <= (("Vd0JLeR4aFshIok" ?
          $unsigned({"VzWxBStBk0LdHmMK1",
              reg1216}) : wire1211) == $signed({reg1233[(3'h7):(2'h3)],
          {$unsigned(reg1217)}}));
      reg1244 <= $unsigned($unsigned(("yiMd3f0" ? "zJ9LOf49" : "")));
    end
  assign wire1245 = {(~^"KoRzgbdN2QPn3RAMV1Z"), $signed("")};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1013
#(parameter param1207 = (8'hb4))
(y, clk, wire1017, wire1016, wire1015, wire1014);
  output wire [(32'haac):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire1017;
  input wire signed [(5'h1a):(1'h0)] wire1016;
  input wire signed [(5'h15):(1'h0)] wire1015;
  input wire [(5'h12):(1'h0)] wire1014;
  reg signed [(3'h4):(1'h0)] reg1206 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1205 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1204 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1203 = (1'h0);
  reg [(5'h17):(1'h0)] reg1202 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1201 = (1'h0);
  reg [(4'hf):(1'h0)] reg1200 = (1'h0);
  reg [(3'h6):(1'h0)] reg1199 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1198 = (1'h0);
  reg [(4'hb):(1'h0)] reg1197 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1196 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1195 = (1'h0);
  reg [(3'h4):(1'h0)] reg1194 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1193 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1192 = (1'h0);
  reg [(3'h5):(1'h0)] reg1191 = (1'h0);
  reg [(4'he):(1'h0)] forvar1189 = (1'h0);
  reg [(5'h17):(1'h0)] reg1190 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1189 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1188 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1187 = (1'h0);
  reg [(5'h16):(1'h0)] reg1186 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1185 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1184 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1183 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1182 = (1'h0);
  reg [(4'h8):(1'h0)] reg1181 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire1180;
  reg signed [(4'hb):(1'h0)] reg1179 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1178 = (1'h0);
  reg [(5'h10):(1'h0)] reg1177 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1176 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1175 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1174 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1173 = (1'h0);
  reg [(3'h7):(1'h0)] reg1172 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1171 = (1'h0);
  reg [(5'h17):(1'h0)] reg1170 = (1'h0);
  reg [(5'h13):(1'h0)] reg1169 = (1'h0);
  reg [(2'h2):(1'h0)] reg1168 = (1'h0);
  wire [(4'hf):(1'h0)] wire1167;
  wire [(5'h10):(1'h0)] wire1166;
  reg signed [(5'h12):(1'h0)] reg1165 = (1'h0);
  reg [(5'h11):(1'h0)] reg1164 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1163 = (1'h0);
  reg [(5'h15):(1'h0)] reg1162 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1161 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1160 = (1'h0);
  reg [(4'hb):(1'h0)] reg1159 = (1'h0);
  reg [(5'h17):(1'h0)] reg1158 = (1'h0);
  reg [(4'he):(1'h0)] reg1157 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1156 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1155 = (1'h0);
  reg [(5'h10):(1'h0)] reg1154 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1153 = (1'h0);
  reg [(3'h6):(1'h0)] reg1152 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1151 = (1'h0);
  reg [(5'h17):(1'h0)] reg1150 = (1'h0);
  reg [(5'h17):(1'h0)] reg1149 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1148 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1147 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1146 = (1'h0);
  reg [(4'h8):(1'h0)] reg1145 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1144 = (1'h0);
  reg [(4'hb):(1'h0)] reg1143 = (1'h0);
  reg [(4'hb):(1'h0)] reg1142 = (1'h0);
  reg [(4'ha):(1'h0)] reg1141 = (1'h0);
  reg [(4'hb):(1'h0)] reg1140 = (1'h0);
  reg [(5'h16):(1'h0)] reg1139 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1138 = (1'h0);
  reg [(5'h18):(1'h0)] reg1137 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1136 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1135 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1134 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1133 = (1'h0);
  reg [(4'hc):(1'h0)] reg1132 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1131 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1130 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1129 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1128 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1127 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1126 = (1'h0);
  reg [(3'h6):(1'h0)] reg1125 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1124 = (1'h0);
  reg [(5'h17):(1'h0)] reg1123 = (1'h0);
  reg [(5'h12):(1'h0)] reg1122 = (1'h0);
  reg [(4'he):(1'h0)] reg1121 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1120 = (1'h0);
  reg [(3'h6):(1'h0)] reg1119 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1118 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1117 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1116 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1115 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1114 = (1'h0);
  reg [(4'hf):(1'h0)] reg1113 = (1'h0);
  reg [(5'h16):(1'h0)] reg1112 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1111 = (1'h0);
  reg [(3'h4):(1'h0)] reg1110 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1109 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1108 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1107 = (1'h0);
  reg [(2'h3):(1'h0)] reg1106 = (1'h0);
  reg [(4'he):(1'h0)] forvar1105 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1104 = (1'h0);
  reg [(4'ha):(1'h0)] reg1103 = (1'h0);
  reg [(5'h19):(1'h0)] reg1102 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1101 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1100 = (1'h0);
  reg [(4'hb):(1'h0)] reg1099 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1098 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1097 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1096 = (1'h0);
  reg [(4'he):(1'h0)] reg1095 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1094 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1093 = (1'h0);
  reg [(4'hb):(1'h0)] reg1092 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1091 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1090 = (1'h0);
  reg [(4'hf):(1'h0)] reg1089 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire1088;
  wire [(3'h6):(1'h0)] wire1087;
  reg [(5'h12):(1'h0)] reg1086 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1085 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1084 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1083 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1082 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1081 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1080 = (1'h0);
  reg [(2'h2):(1'h0)] reg1079 = (1'h0);
  reg [(5'h13):(1'h0)] reg1078 = (1'h0);
  reg [(4'hc):(1'h0)] reg1077 = (1'h0);
  reg [(4'ha):(1'h0)] reg1076 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1075 = (1'h0);
  reg [(5'h16):(1'h0)] reg1074 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1073 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1072 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1071 = (1'h0);
  reg [(4'he):(1'h0)] reg1070 = (1'h0);
  reg [(4'hc):(1'h0)] reg1069 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1068 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1067 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1066 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1065 = (1'h0);
  reg [(5'h15):(1'h0)] reg1064 = (1'h0);
  reg [(4'h9):(1'h0)] reg1063 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1062 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1061 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1060 = (1'h0);
  reg [(4'ha):(1'h0)] reg1059 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1058 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1057 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1056 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1055 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1054 = (1'h0);
  reg [(2'h3):(1'h0)] reg1053 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1052 = (1'h0);
  reg [(3'h6):(1'h0)] reg1051 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1050 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1049 = (1'h0);
  reg [(3'h7):(1'h0)] reg1048 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1047 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1046 = (1'h0);
  reg [(4'h9):(1'h0)] reg1045 = (1'h0);
  reg [(4'he):(1'h0)] reg1044 = (1'h0);
  reg [(5'h15):(1'h0)] reg1043 = (1'h0);
  reg [(2'h3):(1'h0)] reg1042 = (1'h0);
  reg [(4'hd):(1'h0)] reg1041 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1040 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1039 = (1'h0);
  reg [(4'he):(1'h0)] reg1038 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1037 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1036 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1035 = (1'h0);
  reg [(4'hc):(1'h0)] reg1034 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1033 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1032 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1031 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1030 = (1'h0);
  reg [(5'h11):(1'h0)] reg1029 = (1'h0);
  reg [(4'h8):(1'h0)] reg1028 = (1'h0);
  reg [(3'h7):(1'h0)] reg1027 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1026 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1025 = (1'h0);
  reg [(5'h18):(1'h0)] reg1024 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1023 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1022 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1021 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1020 = (1'h0);
  reg [(5'h19):(1'h0)] reg1019 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire1018;
  assign y = {reg1206,
                 reg1205,
                 reg1204,
                 reg1203,
                 reg1202,
                 reg1201,
                 reg1200,
                 reg1199,
                 forvar1198,
                 reg1197,
                 reg1196,
                 forvar1195,
                 reg1194,
                 reg1193,
                 reg1192,
                 reg1191,
                 forvar1189,
                 reg1190,
                 reg1189,
                 reg1188,
                 reg1187,
                 reg1186,
                 reg1185,
                 forvar1184,
                 forvar1183,
                 reg1182,
                 reg1181,
                 wire1180,
                 reg1179,
                 reg1178,
                 reg1177,
                 reg1176,
                 reg1175,
                 reg1174,
                 reg1173,
                 reg1172,
                 forvar1171,
                 reg1170,
                 reg1169,
                 reg1168,
                 wire1167,
                 wire1166,
                 reg1165,
                 reg1164,
                 reg1163,
                 reg1162,
                 reg1161,
                 forvar1160,
                 reg1159,
                 reg1158,
                 reg1157,
                 forvar1156,
                 reg1155,
                 reg1154,
                 forvar1153,
                 reg1152,
                 reg1151,
                 reg1150,
                 reg1149,
                 forvar1148,
                 reg1147,
                 reg1146,
                 reg1145,
                 reg1144,
                 reg1143,
                 reg1142,
                 reg1141,
                 reg1140,
                 reg1139,
                 reg1138,
                 reg1137,
                 reg1136,
                 reg1135,
                 reg1134,
                 forvar1133,
                 reg1132,
                 forvar1131,
                 forvar1130,
                 reg1129,
                 reg1128,
                 reg1127,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1123,
                 reg1122,
                 reg1121,
                 forvar1120,
                 reg1119,
                 forvar1118,
                 reg1117,
                 forvar1116,
                 forvar1115,
                 reg1114,
                 reg1113,
                 reg1112,
                 reg1111,
                 reg1110,
                 reg1109,
                 reg1108,
                 reg1107,
                 reg1106,
                 forvar1105,
                 reg1104,
                 reg1103,
                 reg1102,
                 reg1101,
                 reg1100,
                 reg1099,
                 forvar1098,
                 forvar1097,
                 forvar1096,
                 reg1095,
                 reg1094,
                 reg1093,
                 reg1092,
                 reg1091,
                 reg1090,
                 reg1089,
                 wire1088,
                 wire1087,
                 reg1086,
                 reg1085,
                 reg1084,
                 reg1083,
                 reg1082,
                 reg1081,
                 reg1080,
                 reg1079,
                 reg1078,
                 reg1077,
                 reg1076,
                 reg1075,
                 reg1074,
                 reg1073,
                 reg1072,
                 reg1071,
                 reg1070,
                 reg1069,
                 forvar1068,
                 forvar1067,
                 forvar1066,
                 reg1065,
                 reg1064,
                 reg1063,
                 reg1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 forvar1058,
                 forvar1057,
                 reg1056,
                 reg1055,
                 reg1054,
                 reg1053,
                 forvar1052,
                 reg1051,
                 reg1050,
                 forvar1049,
                 reg1048,
                 forvar1047,
                 reg1046,
                 reg1045,
                 reg1044,
                 reg1043,
                 reg1042,
                 reg1041,
                 reg1040,
                 reg1039,
                 reg1038,
                 reg1037,
                 forvar1036,
                 reg1035,
                 reg1034,
                 forvar1033,
                 reg1032,
                 forvar1031,
                 forvar1030,
                 reg1029,
                 reg1028,
                 reg1027,
                 reg1026,
                 reg1025,
                 reg1024,
                 reg1023,
                 reg1022,
                 reg1021,
                 forvar1020,
                 reg1019,
                 wire1018,
                 (1'h0)};
  assign wire1018 = wire1014[(5'h11):(4'ha)];
  always
    @(posedge clk) begin
      reg1019 <= $signed($unsigned(wire1015[(4'hd):(4'ha)]));
    end
  always
    @(posedge clk) begin
      for (forvar1020 = (1'h0); (forvar1020 < (3'h5)); forvar1020 = (forvar1020 + (1'h1)))
        begin
          reg1021 <= wire1017;
          reg1022 = (~&reg1019);
          reg1023 <= (wire1014 ^ ("bp10CrPCgT0bp" ?
              (($unsigned(reg1019) ? (~&wire1014) : (-(8'hba))) ?
                  ((~reg1019) ?
                      (forvar1020 ? reg1021 : wire1014) : (reg1021 ?
                          forvar1020 : wire1017)) : $signed(wire1014)) : wire1015[(4'hf):(3'h5)]));
          reg1024 <= wire1014;
        end
      reg1025 <= (reg1019 ^ (wire1018 ^~ ($signed((reg1022 ~^ wire1015)) ?
          (reg1019 ? $unsigned(reg1022) : wire1014[(3'h7):(2'h2)]) : ((8'hb1) ?
              (+wire1015) : "0a"))));
      reg1026 <= "xKeox";
      reg1027 <= (8'hb9);
      reg1028 <= wire1018;
      reg1029 <= reg1023;
    end
  always
    @(posedge clk) begin
      for (forvar1030 = (1'h0); (forvar1030 < (1'h0)); forvar1030 = (forvar1030 + (1'h1)))
        begin
          for (forvar1031 = (1'h0); (forvar1031 < (3'h4)); forvar1031 = (forvar1031 + (1'h1)))
            begin
              reg1032 <= (~&$signed((wire1018 > $unsigned((forvar1030 ?
                  reg1026 : wire1015)))));
            end
          for (forvar1033 = (1'h0); (forvar1033 < (2'h3)); forvar1033 = (forvar1033 + (1'h1)))
            begin
              reg1034 = (("RV5YfFGDPFhZD1N0YK7K3c" ?
                  {("hBaXZ9LVNWpHFPULlQVftwlQ" ?
                          (reg1026 << reg1032) : (^wire1018)),
                      $signed($unsigned(reg1023))} : $unsigned((forvar1033 == (reg1021 ^ wire1017)))) >>> forvar1030);
              reg1035 <= $signed(reg1026);
            end
          for (forvar1036 = (1'h0); (forvar1036 < (2'h2)); forvar1036 = (forvar1036 + (1'h1)))
            begin
              reg1037 <= reg1025;
              reg1038 <= wire1017;
              reg1039 <= wire1016;
              if (((!$unsigned("rh5MroIu4QFUB0Rg")) >> $signed(wire1018)))
                begin
                  reg1040 <= (~({$unsigned((~|forvar1033))} - {$unsigned({reg1027,
                          reg1028}),
                      ({reg1038, (7'h48)} ?
                          (wire1016 & (7'h45)) : "YLT2qiP5GmsdXoUPn")}));
                  reg1041 <= {$signed({reg1027, "ZGi8hPMHKfI0QUZI"}), (7'h45)};
                  reg1042 <= $signed(("" ? "ygRw" : reg1039[(4'he):(3'h7)]));
                end
              else
                begin
                  reg1040 <= "3";
                  reg1041 = (wire1018 == (|{(~^(reg1024 << reg1037)),
                      reg1023[(5'h12):(4'ha)]}));
                  reg1042 <= (+reg1041[(2'h2):(2'h2)]);
                  reg1043 = ($unsigned(reg1028) || forvar1030);
                  reg1044 <= ($signed($unsigned("")) ?
                      forvar1030[(4'hc):(4'h9)] : (("MRfID6ivZZ92MGwWAT" || reg1032[(1'h1):(1'h0)]) && ((~|$unsigned(reg1032)) ?
                          (8'hb2) : (&reg1029[(3'h5):(2'h2)]))));
                  reg1045 <= forvar1036;
                end
            end
          reg1046 <= $unsigned($unsigned((8'hb7)));
          for (forvar1047 = (1'h0); (forvar1047 < (2'h3)); forvar1047 = (forvar1047 + (1'h1)))
            begin
              reg1048 <= ($signed(forvar1047[(4'h9):(4'h9)]) << $signed((+({reg1042} ?
                  ((7'h44) ? reg1043 : reg1035) : "8IJ801sr"))));
              for (forvar1049 = (1'h0); (forvar1049 < (3'h5)); forvar1049 = (forvar1049 + (1'h1)))
                begin
                  reg1050 <= $unsigned("LD");
                end
              reg1051 <= wire1018[(2'h3):(1'h1)];
            end
          for (forvar1052 = (1'h0); (forvar1052 < (3'h4)); forvar1052 = (forvar1052 + (1'h1)))
            begin
              reg1053 <= $signed((reg1048 ?
                  (("KguYhk5MNydanxtwKVm" ?
                      "U9oWGEk" : (wire1018 ?
                          reg1038 : reg1028)) > $unsigned($unsigned(reg1048))) : forvar1020[(3'h4):(2'h2)]));
            end
        end
    end
  always
    @(posedge clk) begin
      reg1054 = reg1023;
      reg1055 <= reg1037[(3'h4):(3'h4)];
      reg1056 <= reg1019[(4'hc):(4'h8)];
    end
  always
    @(posedge clk) begin
      for (forvar1057 = (1'h0); (forvar1057 < (1'h1)); forvar1057 = (forvar1057 + (1'h1)))
        begin
          for (forvar1058 = (1'h0); (forvar1058 < (3'h5)); forvar1058 = (forvar1058 + (1'h1)))
            begin
              reg1059 <= "aufSFgT1";
              reg1060 <= $unsigned({((reg1041[(3'h4):(1'h1)] | {reg1021}) ?
                      ((+reg1034) ?
                          (reg1032 ?
                              reg1044 : reg1053) : (~|wire1018)) : reg1046[(1'h1):(1'h0)]),
                  (8'ha1)});
            end
          reg1061 <= "xe";
          if ("")
            begin
              reg1062 = (^forvar1049);
              reg1063 <= $signed({(reg1053[(2'h2):(2'h2)] >>> {"3cpwep2AsBPmbdLPNSN",
                      "m5CXL6A0yOC"}),
                  "ifHalmxf3cGNxe"});
              reg1064 <= {$unsigned((forvar1030[(1'h0):(1'h0)] ?
                      (7'h48) : ({reg1053} != ((7'h4c) ? reg1042 : reg1061)))),
                  $signed($signed((!((7'h42) ~^ forvar1033))))};
              reg1065 <= reg1021[(4'ha):(3'h4)];
            end
          else
            begin
              reg1062 = reg1041[(3'h6):(3'h4)];
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1066 = (1'h0); (forvar1066 < (3'h5)); forvar1066 = (forvar1066 + (1'h1)))
        begin
          for (forvar1067 = (1'h0); (forvar1067 < (3'h5)); forvar1067 = (forvar1067 + (1'h1)))
            begin
              for (forvar1068 = (1'h0); (forvar1068 < (1'h0)); forvar1068 = (forvar1068 + (1'h1)))
                begin
                  reg1069 = (&reg1028[(3'h6):(2'h2)]);
                  reg1070 <= ({($unsigned((reg1025 >>> (8'ha0))) ~^ reg1035)} && wire1018[(2'h3):(2'h3)]);
                  reg1071 <= ((reg1063 ?
                          "T8" : (reg1046[(2'h2):(1'h0)] ?
                              ((forvar1068 & forvar1068) ?
                                  $unsigned(reg1021) : (reg1026 ?
                                      reg1029 : reg1042)) : "H1CpXIpyqiZbApdlA5QR")) ?
                      ((7'h49) ?
                          {reg1035[(4'hf):(4'h9)],
                              ((reg1069 >> (8'hba)) <<< (8'ha9))} : "J4rVt90KzC6pVY9Ab9E9lL") : $unsigned((7'h41)));
                  reg1072 = ("vYf" + (~$unsigned(reg1023[(4'hb):(3'h6)])));
                end
              reg1073 <= reg1060[(4'hb):(2'h3)];
              reg1074 <= "NZEu6P4fkAmAuOHsplfAPA";
            end
          reg1075 <= $signed((^~reg1065[(2'h3):(1'h1)]));
          reg1076 <= "bFJbdmUqd3EyUbYfVK";
          reg1077 <= (+$unsigned(reg1054));
          reg1078 <= $unsigned(forvar1047[(4'hb):(1'h0)]);
        end
      reg1079 <= reg1064[(5'h15):(5'h12)];
      reg1080 = {"0gQW0vBYKuwXF"};
      reg1081 <= $unsigned($unsigned(($unsigned((&reg1019)) + "gIuV8KKdw4")));
      reg1082 <= ((((^((8'hbd) > reg1060)) ?
              {$unsigned(reg1040)} : (&"UGiyWk2xy")) << reg1050[(2'h3):(2'h3)]) ?
          "" : $unsigned((7'h4d)));
      reg1083 <= "vlAqLXFn";
    end
  always
    @(posedge clk) begin
      reg1084 <= $unsigned({"SgyzsywpbGnE0gXpKFXnbl"});
      reg1085 <= "s";
      reg1086 <= (^{"Hd"});
    end
  assign wire1087 = (reg1080 ? "gWgH" : (reg1046 <= forvar1058[(4'ha):(4'ha)]));
  assign wire1088 = $signed(reg1024);
  always
    @(posedge clk) begin
      reg1089 <= $unsigned($signed($unsigned($signed((reg1029 ?
          reg1048 : (8'ha0))))));
      reg1090 <= $unsigned($unsigned("bb3UiBudi"));
      reg1091 <= reg1056;
      reg1092 <= "WYnJwBAS1";
      reg1093 = (reg1023 ^ "5SsCILEAtv2EZN");
      reg1094 = $signed($unsigned((((reg1077 | (8'hba)) ?
              (~|reg1085) : (wire1014 < forvar1058)) ?
          $signed((8'ha1)) : wire1088[(4'h9):(2'h3)])));
    end
  always
    @(posedge clk) begin
      reg1095 <= ((forvar1049[(2'h2):(2'h2)] ?
          (({forvar1058, reg1093} && (forvar1066 <= reg1028)) > (~&(reg1086 ?
              wire1017 : reg1074))) : $unsigned(((reg1034 * forvar1052) <<< {(7'h41),
              reg1093}))) && "5yuwWBd");
      for (forvar1096 = (1'h0); (forvar1096 < (1'h1)); forvar1096 = (forvar1096 + (1'h1)))
        begin
          for (forvar1097 = (1'h0); (forvar1097 < (1'h1)); forvar1097 = (forvar1097 + (1'h1)))
            begin
              for (forvar1098 = (1'h0); (forvar1098 < (1'h0)); forvar1098 = (forvar1098 + (1'h1)))
                begin
                  reg1099 = $unsigned(forvar1057[(3'h4):(3'h4)]);
                  reg1100 = (({(|$signed(reg1043)), $unsigned("esOY0fJVF5")} ?
                      (8'hbf) : ((~&reg1061[(3'h7):(3'h4)]) ?
                          ({reg1028,
                              reg1095} ^ $unsigned(wire1088)) : $signed((~reg1090)))) ^~ forvar1098);
                  reg1101 <= $unsigned(((8'hbf) < reg1094));
                end
              reg1102 <= $signed($unsigned((forvar1067[(3'h4):(1'h1)] ?
                  forvar1057 : (~&(reg1069 * forvar1049)))));
              reg1103 <= (^$signed("zxeJuoQ5DCOVmHrPOhbNuu"));
              reg1104 <= wire1015[(4'hd):(4'hd)];
              for (forvar1105 = (1'h0); (forvar1105 < (1'h0)); forvar1105 = (forvar1105 + (1'h1)))
                begin
                  reg1106 <= ($unsigned(("AoboT" & {(8'hab)})) ?
                      {"wy7pnGrpsoTfFVyoDI",
                          reg1079} : reg1029[(5'h10):(3'h4)]);
                  reg1107 = (^$unsigned(({((8'ha3) <<< reg1083)} - (wire1014 ?
                      $signed(reg1092) : reg1054[(1'h0):(1'h0)]))));
                  reg1108 <= reg1084;
                end
            end
          reg1109 <= reg1045;
          reg1110 <= (~^((reg1042 >= reg1091[(1'h1):(1'h1)]) ~^ reg1085[(3'h5):(1'h1)]));
        end
      reg1111 <= reg1101[(1'h0):(1'h0)];
      reg1112 <= (~^$unsigned(reg1082));
      reg1113 = (~reg1043);
    end
  always
    @(posedge clk) begin
      reg1114 = $signed($unsigned({{wire1016[(4'h9):(2'h3)],
              (reg1078 ? (7'h4e) : forvar1097)},
          ({reg1069, reg1104} && {reg1027})}));
      for (forvar1115 = (1'h0); (forvar1115 < (1'h1)); forvar1115 = (forvar1115 + (1'h1)))
        begin
          for (forvar1116 = (1'h0); (forvar1116 < (1'h0)); forvar1116 = (forvar1116 + (1'h1)))
            begin
              reg1117 = forvar1066[(2'h2):(1'h1)];
              for (forvar1118 = (1'h0); (forvar1118 < (1'h1)); forvar1118 = (forvar1118 + (1'h1)))
                begin
                  reg1119 <= ($unsigned($unsigned("DK")) ?
                      "h4ECdJUGLEgbpOETp6" : $signed({(~|((8'ha5) >> reg1100)),
                          {(^~forvar1067), {reg1101}}}));
                end
              for (forvar1120 = (1'h0); (forvar1120 < (1'h0)); forvar1120 = (forvar1120 + (1'h1)))
                begin
                  reg1121 = ("1msOos8ugDDsY" ?
                      ($signed($unsigned((~|reg1077))) + "c2Q") : "o4PRmUevFIdvHP49");
                  reg1122 = (($signed((8'hb0)) ?
                      $unsigned($unsigned("NruysXFfaI")) : ($unsigned("O04nCJ50CKaq8D8aGWocuVov") ^ ((forvar1105 ^ reg1091) <= "J9TtS72ff2BP8OqML0Q43rtii"))) & reg1064);
                  reg1123 <= {forvar1105, {"Cmect", (^reg1082[(3'h4):(3'h4)])}};
                  reg1124 <= (-{$unsigned(((8'ha8) ? (&reg1061) : (8'hbc))),
                      "OY"});
                end
              reg1125 <= (~^(reg1034 ? (+$unsigned((~|forvar1116))) : (8'hb2)));
              reg1126 <= reg1065[(2'h3):(1'h1)];
            end
        end
      reg1127 <= reg1026[(2'h2):(2'h2)];
      reg1128 <= $unsigned((($unsigned($signed(reg1027)) + "maSaMkhuZ0w7SnXTAR4b3BADW") <= $signed($signed({reg1032,
          reg1038}))));
    end
  always
    @(posedge clk) begin
      reg1129 <= ($signed({$unsigned(((8'hba) <<< reg1084))}) - {($unsigned($signed(reg1111)) ?
              forvar1049 : (^(reg1045 ? reg1032 : reg1100)))});
      for (forvar1130 = (1'h0); (forvar1130 < (2'h2)); forvar1130 = (forvar1130 + (1'h1)))
        begin
          for (forvar1131 = (1'h0); (forvar1131 < (2'h2)); forvar1131 = (forvar1131 + (1'h1)))
            begin
              reg1132 <= reg1061;
              for (forvar1133 = (1'h0); (forvar1133 < (2'h2)); forvar1133 = (forvar1133 + (1'h1)))
                begin
                  reg1134 <= $unsigned(reg1092);
                  reg1135 <= ((($signed({reg1078}) <<< $signed($unsigned((8'hbc)))) ?
                      (reg1023 ?
                          reg1021 : reg1060) : $signed(reg1134[(1'h1):(1'h0)])) >>> $signed(reg1132));
                end
              reg1136 <= reg1079;
              if ("Mq1TWldH9xJgQKU8lTom5XlFG")
                begin
                  reg1137 <= reg1028[(4'h8):(4'h8)];
                  reg1138 <= (-{$signed(reg1085)});
                  reg1139 <= reg1048;
                  reg1140 <= ($signed(reg1137) && "8ow");
                  reg1141 <= ($unsigned(reg1083) ~^ $unsigned(((reg1051 ?
                          "n2CZcipqsJRfh" : reg1043[(1'h1):(1'h0)]) ?
                      reg1128[(3'h5):(2'h2)] : forvar1105[(4'hb):(3'h6)])));
                  reg1142 <= reg1055;
                end
              else
                begin
                  reg1137 <= {(~^"Prwm9HRdzAa3SFe2dU1Ov"),
                      wire1015[(4'hf):(4'h9)]};
                  reg1138 <= (reg1053[(1'h0):(1'h0)] ~^ $signed((((|reg1028) ?
                      ((8'hb5) & reg1021) : {(7'h41)}) & reg1107)));
                  reg1139 <= reg1061;
                  reg1140 <= (^"l63p8DnF3L2");
                  reg1141 = $signed($signed($unsigned($unsigned((^reg1137)))));
                end
              reg1143 <= "HdZdp8TCFqzTtwHII";
              reg1144 <= $unsigned($unsigned((reg1069[(2'h3):(1'h1)] ?
                  ($signed(forvar1097) ~^ (reg1029 * forvar1057)) : (reg1046 > {reg1054}))));
            end
          reg1145 <= $signed(reg1106[(2'h2):(2'h2)]);
          reg1146 = (^reg1056);
          reg1147 <= (^~{reg1048});
          for (forvar1148 = (1'h0); (forvar1148 < (3'h5)); forvar1148 = (forvar1148 + (1'h1)))
            begin
              reg1149 = {forvar1130, $unsigned((~|$signed("wpU9IJXhfB")))};
            end
          reg1150 <= forvar1058[(4'ha):(2'h3)];
        end
      reg1151 <= {forvar1148};
      reg1152 <= reg1126;
      for (forvar1153 = (1'h0); (forvar1153 < (2'h2)); forvar1153 = (forvar1153 + (1'h1)))
        begin
          reg1154 <= $signed(($signed({$unsigned(reg1041),
              reg1127[(1'h1):(1'h1)]}) << (~^{(reg1064 ? forvar1068 : reg1145),
              ((8'haa) || (8'hb0))})));
        end
      reg1155 <= ("57g5zRulN1" >= $unsigned(reg1109));
    end
  always
    @(posedge clk) begin
      for (forvar1156 = (1'h0); (forvar1156 < (1'h0)); forvar1156 = (forvar1156 + (1'h1)))
        begin
          reg1157 <= (("ncQ5oRbx5UTERMJAHs7IqGi" ?
                  $unsigned((~(reg1046 ?
                      (8'hb9) : (8'hb5)))) : wire1087[(1'h0):(1'h0)]) ?
              (|reg1135[(2'h2):(2'h2)]) : $unsigned(($signed((~&wire1015)) ?
                  reg1154 : reg1078)));
          reg1158 = (8'hb8);
          reg1159 = reg1104[(1'h0):(1'h0)];
          for (forvar1160 = (1'h0); (forvar1160 < (3'h4)); forvar1160 = (forvar1160 + (1'h1)))
            begin
              reg1161 <= (~&"II0fbdxh7HaAtlkuC");
            end
        end
      reg1162 <= {$unsigned(("cRMW6oniH2462" ?
              {{reg1157, wire1014},
                  "MShZcX"} : $unsigned("390uuXGWtxWC3aHVrFB"))),
          (!($unsigned((forvar1096 ? reg1117 : reg1151)) ?
              $unsigned(forvar1033[(2'h3):(1'h1)]) : reg1129))};
      reg1163 <= wire1088[(5'h11):(4'h9)];
      reg1164 <= reg1076[(3'h6):(2'h2)];
      reg1165 <= reg1142[(4'h9):(2'h2)];
    end
  assign wire1166 = "RrtM9p2D7PWBHaUeHNfMtPDJ";
  assign wire1167 = (((~&$signed((reg1056 != wire1166))) ^ "AivbOeuGt80Z1opRYf") ?
                        ({$signed({reg1038, reg1126}),
                            (~&$unsigned(reg1117))} + forvar1153[(4'hd):(3'h7)]) : forvar1058);
  always
    @(posedge clk) begin
      reg1168 <= reg1037;
      reg1169 <= "HssOOP3Crf";
    end
  always
    @(posedge clk) begin
      reg1170 <= (((~^(!(forvar1068 | reg1064))) <<< "17aYznawrLIs0ayL3wTv") ?
          {reg1076, reg1137} : ((({reg1126, reg1150} ?
                      {reg1110, reg1141} : forvar1116[(4'he):(4'hc)]) ?
                  "m1WV0hIOJF" : $unsigned(reg1107[(3'h4):(2'h2)])) ?
              (+(!{reg1101, forvar1105})) : ({"OhbtTmk3O4"} ?
                  (^~reg1159) : reg1094)));
    end
  always
    @(posedge clk) begin
      for (forvar1171 = (1'h0); (forvar1171 < (2'h2)); forvar1171 = (forvar1171 + (1'h1)))
        begin
          reg1172 <= (7'h41);
          reg1173 <= reg1086[(4'hb):(2'h2)];
        end
    end
  always
    @(posedge clk) begin
      reg1174 <= reg1106[(1'h0):(1'h0)];
      reg1175 <= "SMo";
      reg1176 = $unsigned(reg1102[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg1177 = $signed((forvar1057[(1'h0):(1'h0)] ? "Uh" : "RM"));
      reg1178 <= {$signed(reg1029[(3'h4):(2'h2)]),
          $unsigned(("WnP" > $unsigned((reg1145 ? reg1176 : reg1150))))};
      reg1179 <= $signed(reg1041);
    end
  assign wire1180 = $unsigned("nhSoqDfBmBykP3BMEtG");
  always
    @(posedge clk) begin
      reg1181 <= reg1073[(2'h3):(2'h3)];
      reg1182 <= (~((&(reg1078 >>> reg1119)) ?
          forvar1160[(3'h4):(1'h0)] : reg1042));
      for (forvar1183 = (1'h0); (forvar1183 < (1'h0)); forvar1183 = (forvar1183 + (1'h1)))
        begin
          if ({reg1044})
            begin
              for (forvar1184 = (1'h0); (forvar1184 < (3'h5)); forvar1184 = (forvar1184 + (1'h1)))
                begin
                  reg1185 <= (+"44H17ALbLd");
                  reg1186 <= reg1143[(3'h7):(3'h5)];
                end
              reg1187 <= ("WwqqPzRK2PwFwbHnh" + $signed("FH0Y5tb"));
              reg1188 <= $unsigned((~&($unsigned("dxLvXrv32ACs") ?
                  reg1056 : (8'ha2))));
              reg1189 = (&(~reg1050));
              reg1190 <= (reg1070[(1'h0):(1'h0)] ?
                  forvar1148[(4'h8):(3'h7)] : (~reg1095[(2'h3):(2'h3)]));
            end
          else
            begin
              for (forvar1184 = (1'h0); (forvar1184 < (2'h2)); forvar1184 = (forvar1184 + (1'h1)))
                begin
                  reg1185 = reg1124;
                  reg1186 = ("kHwKPBtnW5ffzgJwZ" ?
                      $unsigned("iuDD8d3rB3aQ05PTQ1") : reg1150[(1'h1):(1'h1)]);
                  reg1187 = $signed((-{((reg1158 < reg1128) - (7'h4a)),
                      forvar1130[(2'h2):(1'h0)]}));
                  reg1188 <= ((+(|($signed(reg1146) << "W2rZHxwcrWHIHCqz7Y"))) ?
                      $signed({($unsigned(reg1059) ?
                              reg1048[(1'h1):(1'h0)] : (reg1186 ?
                                  reg1140 : reg1102)),
                          $signed(forvar1057[(3'h5):(2'h3)])}) : (~^{{reg1123}}));
                end
              for (forvar1189 = (1'h0); (forvar1189 < (2'h3)); forvar1189 = (forvar1189 + (1'h1)))
                begin
                  reg1190 <= (~|forvar1183[(2'h3):(2'h2)]);
                  reg1191 <= "y";
                  reg1192 <= "DGi0";
                end
              reg1193 = "31r";
              reg1194 <= ((8'h9e) ?
                  (!$unsigned({(reg1034 - (7'h40)),
                      reg1084[(5'h14):(4'hf)]})) : "wXb3LDyItO1hHJb7lw88sd");
              for (forvar1195 = (1'h0); (forvar1195 < (3'h4)); forvar1195 = (forvar1195 + (1'h1)))
                begin
                  reg1196 <= (~^(|$unsigned((&forvar1098[(5'h14):(4'hf)]))));
                end
            end
          reg1197 <= (~"4ufTuG");
          for (forvar1198 = (1'h0); (forvar1198 < (2'h3)); forvar1198 = (forvar1198 + (1'h1)))
            begin
              reg1199 <= $unsigned("pgYZOXGF");
              reg1200 <= ((^"0rrTCo4iuvoN5TKBdp") <= reg1145[(3'h5):(1'h0)]);
              reg1201 <= ($signed(("Gl5WHAl8iPNlX3h0S" ?
                      $signed($signed(reg1158)) : $signed((reg1135 <= forvar1116)))) ?
                  "7" : ($unsigned("KplJVMpn54gMFO") ?
                      $unsigned("LxIHFZbOByvWRPch") : reg1172));
              reg1202 <= ($signed($unsigned((~&(7'h48)))) >> ($signed($unsigned((reg1114 == reg1168))) ?
                  $unsigned(reg1178) : ("48m4TfxnN" ~^ {((8'haa) ?
                          reg1174 : reg1112)})));
              reg1203 <= "CrrQu2k";
            end
          reg1204 <= (-$signed(reg1145));
        end
      reg1205 = (reg1145 < (!("" ?
          $unsigned((+reg1185)) : $signed("DNwamxAszV7yabdY75TWsPQxr"))));
      reg1206 = $signed(($unsigned((^~(reg1078 ? reg1040 : (7'h42)))) ?
          (-({reg1073} ?
              {reg1126, reg1032} : (reg1147 ?
                  reg1109 : (8'ha7)))) : {({reg1128} >= reg1161[(4'hf):(3'h7)])}));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module984
#( parameter param1010 = ((!((((7'h45) ? (7'h40) : (8'h9c)) >>> (8'ha6)) ? {((8'hae) + (8'ha0)), (|(7'h4b))} : ({(8'hbc), (7'h44)} ? ((7'h41) >>> (7'h4b)) : ((7'h48) ? (8'h9d) : (7'h48))))) ~^ (^((((8'hbe) ? (8'had) : (7'h48)) ? (8'ha6) : {(8'ha7), (7'h41)}) ? (((8'ha6) != (8'hb4)) != ((8'h9f) ? (8'hb7) : (8'h9f))) : (!((8'hb8) ? (8'ha5) : (8'h9e)))))) )
(y, clk, wire988, wire987, wire986, wire985);
  output wire [(32'h146):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire988;
  input wire [(3'h5):(1'h0)] wire987;
  input wire signed [(5'h12):(1'h0)] wire986;
  input wire signed [(5'h18):(1'h0)] wire985;
  wire signed [(5'h1a):(1'h0)] wire1009;
  reg [(5'h17):(1'h0)] reg1008 = (1'h0);
  reg [(4'he):(1'h0)] reg1007 = (1'h0);
  reg [(5'h11):(1'h0)] reg1006 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1005 = (1'h0);
  reg [(5'h17):(1'h0)] reg1004 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1003 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1002 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1001 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1000 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg999 = (1'h0);
  reg [(5'h16):(1'h0)] reg998 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg997 = (1'h0);
  reg [(4'hc):(1'h0)] reg996 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg995 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg994 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg993 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg992 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg991 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg990 = (1'h0);
  reg [(3'h4):(1'h0)] reg989 = (1'h0);
  assign y = {wire1009,
                 reg1008,
                 reg1007,
                 reg1006,
                 reg1005,
                 reg1004,
                 reg1003,
                 reg1002,
                 reg1001,
                 reg1000,
                 reg999,
                 reg998,
                 reg997,
                 reg996,
                 reg995,
                 reg994,
                 reg993,
                 reg992,
                 reg991,
                 reg990,
                 reg989,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg989 = ($signed({wire985, $signed((8'ha9))}) != wire986[(4'h8):(3'h4)]);
      reg990 <= wire985;
      reg991 <= $signed(((^$signed($signed(wire986))) ?
          "LyYzW5dBUaxc9q2Dhp1Z" : $unsigned($unsigned($unsigned(wire988)))));
      reg992 = {"rc"};
      reg993 <= wire986;
    end
  always
    @(posedge clk) begin
      reg994 <= reg991;
    end
  always
    @(posedge clk) begin
      reg995 <= (reg991[(1'h1):(1'h1)] & $signed({$unsigned((!reg989)),
          reg990}));
    end
  always
    @(posedge clk) begin
      reg996 <= $unsigned(($signed(("6YV6NPOVrqP3kWE5qi" ?
          $unsigned(reg989) : "UQhEX5uwGmM8i13Y8Ix3")) ^~ wire985[(3'h7):(3'h7)]));
      reg997 = $signed($signed({wire986[(5'h10):(1'h1)], reg991}));
      reg998 = "yYhtAwJly9N4VIQlyAWNad46b";
    end
  always
    @(posedge clk) begin
      reg999 <= (8'hb2);
      reg1000 <= ({reg995[(1'h0):(1'h0)]} != (($unsigned((~|reg990)) ?
              "GO4bmoouQEmDmd6upHqh" : (+(wire986 < reg995))) ?
          $signed($unsigned($unsigned(reg992))) : "prULfYmgIqtHLzZyl63w6"));
      reg1001 <= (-$unsigned("LBs3kpHR2dutnmVnA6MX"));
      reg1002 <= $unsigned($signed((7'h42)));
      reg1003 <= reg990;
      reg1004 <= (($signed($signed({reg990, (8'haa)})) ?
          {$signed((~^(8'hb6))),
              "zUReIYlge"} : $signed(reg1001)) <= $signed($signed($unsigned($signed(reg993)))));
    end
  always
    @(posedge clk) begin
      reg1005 = $signed($unsigned({(((8'h9d) ? wire987 : reg993) ?
              ((8'ha2) ? wire986 : reg990) : "oDg603hoYoszPvC0IJUAi")}));
      reg1006 <= (reg1002[(2'h2):(1'h1)] ?
          "J0YxB5ATv8LDXv" : $unsigned(($unsigned($signed(reg999)) ~^ $signed(wire986))));
      reg1007 = (reg993 ? "Lw0eqIeWHHZAY5u" : reg995[(2'h3):(2'h2)]);
      reg1008 = {reg1000};
    end
  assign wire1009 = $signed(((((reg1003 ? reg993 : (8'h9d)) ?
                            "hLsr74rwwWUBVJ" : $unsigned((8'hab))) ?
                        $unsigned((~|reg992)) : $unsigned((reg1004 >> reg994))) - "dMVP3WNmmUoCkTx4aYmFRCyOD"));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module779  (y, clk, wire783, wire782, wire781, wire780);
  output wire [(32'hb40):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire783;
  input wire signed [(4'h8):(1'h0)] wire782;
  input wire [(4'he):(1'h0)] wire781;
  input wire signed [(5'h1a):(1'h0)] wire780;
  reg signed [(5'h19):(1'h0)] reg981 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg980 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg979 = (1'h0);
  reg [(5'h19):(1'h0)] reg978 = (1'h0);
  reg [(3'h6):(1'h0)] reg977 = (1'h0);
  reg [(4'hd):(1'h0)] reg976 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg975 = (1'h0);
  reg [(5'h14):(1'h0)] reg974 = (1'h0);
  reg [(4'hf):(1'h0)] forvar973 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg972 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar971 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg970 = (1'h0);
  reg [(4'he):(1'h0)] forvar969 = (1'h0);
  reg [(5'h19):(1'h0)] reg968 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg967 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg966 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar965 = (1'h0);
  reg [(3'h6):(1'h0)] forvar964 = (1'h0);
  reg [(5'h17):(1'h0)] reg963 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg962 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg961 = (1'h0);
  reg [(4'hb):(1'h0)] reg960 = (1'h0);
  reg [(5'h18):(1'h0)] reg959 = (1'h0);
  reg [(2'h3):(1'h0)] reg958 = (1'h0);
  reg [(5'h16):(1'h0)] reg957 = (1'h0);
  reg [(5'h12):(1'h0)] reg956 = (1'h0);
  reg [(5'h19):(1'h0)] forvar955 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg954 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg953 = (1'h0);
  reg [(4'hd):(1'h0)] reg952 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg951 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg950 = (1'h0);
  reg [(5'h16):(1'h0)] reg949 = (1'h0);
  reg [(3'h5):(1'h0)] reg948 = (1'h0);
  reg [(5'h13):(1'h0)] reg947 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg946 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar945 = (1'h0);
  reg [(4'hb):(1'h0)] reg944 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg943 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar942 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg941 = (1'h0);
  reg [(5'h15):(1'h0)] reg940 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg939 = (1'h0);
  reg [(4'hd):(1'h0)] reg938 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg937 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar936 = (1'h0);
  reg [(5'h1a):(1'h0)] reg935 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg934 = (1'h0);
  reg [(5'h13):(1'h0)] reg933 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg932 = (1'h0);
  reg [(5'h19):(1'h0)] forvar931 = (1'h0);
  reg [(4'he):(1'h0)] reg930 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg929 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg928 = (1'h0);
  reg [(4'h9):(1'h0)] forvar927 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg926 = (1'h0);
  reg [(4'he):(1'h0)] reg925 = (1'h0);
  reg [(5'h13):(1'h0)] reg924 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg923 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar922 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg921 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg920 = (1'h0);
  reg [(5'h1a):(1'h0)] reg919 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg918 = (1'h0);
  reg [(3'h7):(1'h0)] reg917 = (1'h0);
  reg [(5'h13):(1'h0)] forvar916 = (1'h0);
  reg [(5'h18):(1'h0)] reg915 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar914 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg913 = (1'h0);
  reg [(4'hc):(1'h0)] reg912 = (1'h0);
  reg [(4'he):(1'h0)] reg911 = (1'h0);
  reg [(5'h15):(1'h0)] reg910 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg909 = (1'h0);
  reg [(4'he):(1'h0)] reg908 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar907 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar906 = (1'h0);
  reg [(2'h2):(1'h0)] reg905 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg904 = (1'h0);
  reg [(5'h12):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg902 = (1'h0);
  reg [(5'h14):(1'h0)] reg901 = (1'h0);
  reg [(4'h8):(1'h0)] reg900 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar899 = (1'h0);
  reg [(4'ha):(1'h0)] reg898 = (1'h0);
  reg [(5'h1a):(1'h0)] reg897 = (1'h0);
  reg [(5'h16):(1'h0)] forvar896 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg895 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg894 = (1'h0);
  reg [(4'h8):(1'h0)] reg893 = (1'h0);
  reg [(4'h8):(1'h0)] reg892 = (1'h0);
  reg [(5'h10):(1'h0)] reg891 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg890 = (1'h0);
  wire [(5'h13):(1'h0)] wire889;
  reg [(3'h6):(1'h0)] reg888 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg887 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg886 = (1'h0);
  reg [(5'h15):(1'h0)] reg885 = (1'h0);
  reg [(5'h12):(1'h0)] reg884 = (1'h0);
  reg [(5'h19):(1'h0)] reg883 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg882 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg881 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg880 = (1'h0);
  reg [(5'h15):(1'h0)] reg879 = (1'h0);
  reg [(3'h6):(1'h0)] forvar878 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg877 = (1'h0);
  reg [(5'h18):(1'h0)] reg876 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg875 = (1'h0);
  reg [(3'h7):(1'h0)] reg874 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar873 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg872 = (1'h0);
  reg [(5'h15):(1'h0)] forvar871 = (1'h0);
  reg [(4'h9):(1'h0)] forvar870 = (1'h0);
  reg [(4'ha):(1'h0)] reg869 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg868 = (1'h0);
  reg [(5'h16):(1'h0)] reg867 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg866 = (1'h0);
  reg [(5'h10):(1'h0)] reg865 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg864 = (1'h0);
  reg [(4'h8):(1'h0)] reg863 = (1'h0);
  reg [(4'h9):(1'h0)] reg862 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg861 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg860 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar859 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg858 = (1'h0);
  reg [(5'h1a):(1'h0)] reg857 = (1'h0);
  reg [(2'h2):(1'h0)] reg856 = (1'h0);
  reg [(4'h9):(1'h0)] reg855 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg854 = (1'h0);
  reg [(3'h5):(1'h0)] reg853 = (1'h0);
  reg [(5'h12):(1'h0)] reg852 = (1'h0);
  reg [(3'h4):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg850 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg849 = (1'h0);
  reg [(2'h2):(1'h0)] forvar848 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg847 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg846 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg845 = (1'h0);
  reg [(3'h6):(1'h0)] reg844 = (1'h0);
  reg [(4'hd):(1'h0)] forvar843 = (1'h0);
  reg [(4'hc):(1'h0)] forvar842 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg841 = (1'h0);
  reg [(5'h1a):(1'h0)] reg840 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire839;
  reg [(4'hf):(1'h0)] reg838 = (1'h0);
  reg [(3'h6):(1'h0)] reg837 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg836 = (1'h0);
  reg [(4'hd):(1'h0)] reg835 = (1'h0);
  reg [(4'hc):(1'h0)] reg834 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg833 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg832 = (1'h0);
  reg [(3'h4):(1'h0)] reg831 = (1'h0);
  reg [(5'h12):(1'h0)] reg830 = (1'h0);
  reg [(4'hd):(1'h0)] forvar829 = (1'h0);
  reg [(2'h2):(1'h0)] forvar828 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg827 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg826 = (1'h0);
  reg [(4'hb):(1'h0)] forvar825 = (1'h0);
  reg [(5'h18):(1'h0)] reg824 = (1'h0);
  reg [(5'h1a):(1'h0)] reg823 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg822 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar821 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg820 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar807 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg819 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg818 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar810 = (1'h0);
  reg [(5'h1a):(1'h0)] reg809 = (1'h0);
  reg [(5'h15):(1'h0)] reg817 = (1'h0);
  reg [(3'h4):(1'h0)] reg816 = (1'h0);
  reg [(4'ha):(1'h0)] reg815 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg814 = (1'h0);
  reg [(4'h9):(1'h0)] reg813 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg812 = (1'h0);
  reg [(5'h14):(1'h0)] reg811 = (1'h0);
  reg [(3'h7):(1'h0)] reg810 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar809 = (1'h0);
  reg [(4'ha):(1'h0)] reg808 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg807 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg806 = (1'h0);
  reg signed [(4'he):(1'h0)] reg805 = (1'h0);
  reg [(2'h3):(1'h0)] reg804 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg803 = (1'h0);
  reg [(4'hf):(1'h0)] reg802 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg801 = (1'h0);
  reg [(5'h16):(1'h0)] reg800 = (1'h0);
  reg [(5'h14):(1'h0)] reg799 = (1'h0);
  reg [(2'h3):(1'h0)] reg798 = (1'h0);
  reg [(2'h2):(1'h0)] reg797 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg796 = (1'h0);
  reg [(2'h3):(1'h0)] reg795 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg794 = (1'h0);
  wire [(5'h16):(1'h0)] wire793;
  wire [(4'he):(1'h0)] wire792;
  wire [(5'h14):(1'h0)] wire791;
  wire [(5'h14):(1'h0)] wire790;
  reg signed [(5'h19):(1'h0)] reg789 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg788 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg787 = (1'h0);
  reg [(3'h5):(1'h0)] reg786 = (1'h0);
  wire [(4'h8):(1'h0)] wire785;
  wire [(4'ha):(1'h0)] wire784;
  assign y = {reg981,
                 reg980,
                 reg979,
                 reg978,
                 reg977,
                 reg976,
                 reg975,
                 reg974,
                 forvar973,
                 reg972,
                 forvar971,
                 reg970,
                 forvar969,
                 reg968,
                 reg967,
                 reg966,
                 forvar965,
                 forvar964,
                 reg963,
                 reg962,
                 reg961,
                 reg960,
                 reg959,
                 reg958,
                 reg957,
                 reg956,
                 forvar955,
                 reg954,
                 reg953,
                 reg952,
                 reg951,
                 reg950,
                 reg949,
                 reg948,
                 reg947,
                 reg946,
                 forvar945,
                 reg944,
                 reg943,
                 forvar942,
                 reg941,
                 reg940,
                 reg939,
                 reg938,
                 reg937,
                 forvar936,
                 reg935,
                 reg934,
                 reg933,
                 reg932,
                 forvar931,
                 reg930,
                 reg929,
                 reg928,
                 forvar927,
                 reg926,
                 reg925,
                 reg924,
                 reg923,
                 forvar922,
                 reg921,
                 reg920,
                 reg919,
                 reg918,
                 reg917,
                 forvar916,
                 reg915,
                 forvar914,
                 reg913,
                 reg912,
                 reg911,
                 reg910,
                 reg909,
                 reg908,
                 forvar907,
                 forvar906,
                 reg905,
                 reg904,
                 reg903,
                 reg902,
                 reg901,
                 reg900,
                 forvar899,
                 reg898,
                 reg897,
                 forvar896,
                 reg895,
                 reg894,
                 reg893,
                 reg892,
                 reg891,
                 reg890,
                 wire889,
                 reg888,
                 reg887,
                 reg886,
                 reg885,
                 reg884,
                 reg883,
                 reg882,
                 reg881,
                 reg880,
                 reg879,
                 forvar878,
                 reg877,
                 reg876,
                 reg875,
                 reg874,
                 forvar873,
                 reg872,
                 forvar871,
                 forvar870,
                 reg869,
                 reg868,
                 reg867,
                 reg866,
                 reg865,
                 reg864,
                 reg863,
                 reg862,
                 reg861,
                 reg860,
                 forvar859,
                 reg858,
                 reg857,
                 reg856,
                 reg855,
                 reg854,
                 reg853,
                 reg852,
                 reg851,
                 reg850,
                 reg849,
                 forvar848,
                 reg847,
                 reg846,
                 reg845,
                 reg844,
                 forvar843,
                 forvar842,
                 reg841,
                 reg840,
                 wire839,
                 reg838,
                 reg837,
                 reg836,
                 reg835,
                 reg834,
                 reg833,
                 reg832,
                 reg831,
                 reg830,
                 forvar829,
                 forvar828,
                 reg827,
                 reg826,
                 forvar825,
                 reg824,
                 reg823,
                 reg822,
                 forvar821,
                 reg820,
                 forvar807,
                 reg819,
                 reg818,
                 forvar810,
                 reg809,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 reg812,
                 reg811,
                 reg810,
                 forvar809,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg802,
                 reg801,
                 reg800,
                 reg799,
                 reg798,
                 reg797,
                 reg796,
                 reg795,
                 reg794,
                 wire793,
                 wire792,
                 wire791,
                 wire790,
                 reg789,
                 reg788,
                 reg787,
                 reg786,
                 wire785,
                 wire784,
                 (1'h0)};
  assign wire784 = wire781;
  assign wire785 = wire781[(3'h5):(2'h3)];
  always
    @(posedge clk) begin
      reg786 = wire781;
      reg787 <= wire780;
      reg788 <= (reg786[(1'h1):(1'h1)] << $unsigned(("R5isGEK9" >= $unsigned(wire784[(3'h7):(2'h3)]))));
      reg789 = wire783[(1'h1):(1'h0)];
    end
  assign wire790 = wire785[(4'h8):(2'h3)];
  assign wire791 = wire783;
  assign wire792 = $signed($unsigned(wire781));
  assign wire793 = $signed((-$signed("s1E")));
  always
    @(posedge clk) begin
      reg794 = wire780[(5'h19):(2'h3)];
      reg795 <= ("YleeF7I2m6BQ49mkvu" ?
          (((!{wire781, wire791}) ?
                  ("P7qbktVe" <= (wire784 >> wire781)) : $signed(wire790)) ?
              wire783 : $signed($signed((wire782 ?
                  reg788 : wire791)))) : wire780);
    end
  always
    @(posedge clk) begin
      reg796 <= ((~"QL2lvQtqY1rq81Gl5qDrOGf") ?
          $unsigned(($unsigned((wire784 << reg794)) ?
              (~"7qSZOoDys0DaKF") : "M3KU")) : (^(!(!"4inPGO"))));
      reg797 <= $signed(((&("rA0zyE3" ?
          $unsigned(wire780) : (wire783 ^ wire790))) >= ($signed(reg788[(2'h3):(2'h3)]) ^~ ((8'hb9) ^~ reg787[(3'h4):(1'h1)]))));
      reg798 = $unsigned((&""));
    end
  always
    @(posedge clk) begin
      reg799 <= ({((+$unsigned((8'ha2))) * reg797),
          reg798} <= reg797[(1'h0):(1'h0)]);
      reg800 = ($signed(reg786) + ((^wire793) > "q4qtFrbzRYKTOcNZOV4H57"));
      reg801 <= "T";
      reg802 <= (~$unsigned((reg801[(4'he):(4'h9)] ?
          "b3" : $signed({(7'h41), reg786}))));
    end
  always
    @(posedge clk) begin
      reg803 = ($unsigned(($signed((reg800 ?
              wire790 : wire783)) != wire781[(3'h5):(3'h5)])) ?
          "rTqraqr2Ct" : "16lBx5i3NYPy");
      if ($signed("swlIWO9lg0RR6f6zenIVpYowZ"))
        begin
          reg804 = $signed($signed(reg803));
          reg805 = $unsigned(wire784);
          reg806 <= $signed("HPlITf1XwmuvlrkFU");
          if ("URr")
            begin
              reg807 <= (&($signed("FX2OuJ2E8wJdhq") ~^ ({(7'h46)} ?
                  (wire785 || (|wire780)) : $unsigned($signed(reg803)))));
              reg808 <= (~^"ZZYYZc4Ia8LX1sooubGS3Il");
              for (forvar809 = (1'h0); (forvar809 < (3'h5)); forvar809 = (forvar809 + (1'h1)))
                begin
                  reg810 = (reg786[(3'h4):(1'h0)] ?
                      "46" : $unsigned((-reg787[(5'h14):(4'hf)])));
                  reg811 <= (reg788 >= (~|"L7M4C2LGBX"));
                  reg812 <= (reg800 ?
                      (7'h41) : (wire790 >= reg797[(1'h1):(1'h0)]));
                  reg813 <= $unsigned({reg800[(2'h3):(1'h0)], reg787});
                  reg814 <= "GWc8a1N8nLXSRYSN";
                  reg815 <= reg801[(3'h4):(1'h1)];
                end
              reg816 = $signed((&({reg805[(3'h6):(2'h3)],
                  "WWZY1Hm1"} && ((^~reg801) < $unsigned(wire782)))));
              reg817 <= (7'h4d);
            end
          else
            begin
              reg807 <= $signed(wire793[(1'h0):(1'h0)]);
              reg808 <= (reg794 ?
                  $unsigned({{(-reg788), $signed(reg799)},
                      (-$signed((8'ha5)))}) : $signed($signed("C5m6rJ4")));
              reg809 <= wire791;
              for (forvar810 = (1'h0); (forvar810 < (1'h1)); forvar810 = (forvar810 + (1'h1)))
                begin
                  reg811 = $signed((~&($signed($unsigned(wire790)) ?
                      (8'hb3) : $unsigned("S28eVVUp4a"))));
                  reg812 = ((-(((+forvar810) ?
                              wire783 : "xKklPCuvAMbcNgk3VvzAch") ?
                          $unsigned(reg816) : reg787)) ?
                      (8'haa) : reg811[(5'h11):(4'hf)]);
                  reg813 <= (((-{(reg807 ? reg814 : (8'ha1))}) + ("3t19U9vK" ?
                          $signed((7'h4e)) : "CBNQfQq0YfOC0n")) ?
                      reg813 : {reg798});
                  reg814 <= reg810;
                end
              reg815 <= $signed($signed({reg788}));
            end
          reg818 <= $signed(reg801);
          reg819 <= $unsigned((~^"NIJzEIIugbXXoRxNl"));
        end
      else
        begin
          reg804 <= $unsigned({($unsigned({reg819, (8'hb3)}) ?
                  wire785[(4'h8):(1'h0)] : ($signed(reg812) ?
                      wire791 : wire783[(3'h5):(3'h4)])),
              (reg808 + {((8'h9d) ~^ (8'hbc))})});
          reg805 <= "WG43tKCG";
          reg806 = {$signed(wire785)};
          for (forvar807 = (1'h0); (forvar807 < (2'h3)); forvar807 = (forvar807 + (1'h1)))
            begin
              reg808 <= $unsigned((~^(~&(+reg809))));
              for (forvar809 = (1'h0); (forvar809 < (2'h3)); forvar809 = (forvar809 + (1'h1)))
                begin
                  reg810 = $unsigned((&$signed(reg803)));
                  reg811 <= reg787[(5'h14):(4'hb)];
                  reg812 <= (~"XVM");
                end
              reg813 <= "pT4";
              reg814 <= (+((wire780 >>> "VfqtN7gPw4qTrPbvm3") ?
                  (~&wire793) : $unsigned("neNWvSgCaz")));
            end
          reg815 = "lk9qAt1WeZlqZLqtV18TAs";
          reg816 <= (!{$unsigned(reg800[(5'h10):(4'hd)])});
        end
      reg820 <= reg796[(5'h11):(4'h8)];
      for (forvar821 = (1'h0); (forvar821 < (1'h0)); forvar821 = (forvar821 + (1'h1)))
        begin
          reg822 <= $unsigned(((($signed(reg786) >= (~^reg819)) ?
                  reg802 : $signed({wire790})) ?
              (^~$signed({(7'h42), (7'h49)})) : reg817[(5'h11):(2'h2)]));
        end
    end
  always
    @(posedge clk) begin
      reg823 = reg811[(3'h6):(3'h5)];
      reg824 <= (~"L3gd3");
    end
  always
    @(posedge clk) begin
      for (forvar825 = (1'h0); (forvar825 < (2'h2)); forvar825 = (forvar825 + (1'h1)))
        begin
          reg826 <= $unsigned(wire790[(4'hb):(4'h8)]);
          reg827 <= ($unsigned((~($unsigned(wire781) ?
              $signed((8'ha9)) : {reg796, reg788}))) ^~ {$unsigned(reg826),
              ({reg823[(5'h16):(5'h14)]} ?
                  reg799 : {{reg822}, reg797[(1'h0):(1'h0)]})});
          for (forvar828 = (1'h0); (forvar828 < (2'h3)); forvar828 = (forvar828 + (1'h1)))
            begin
              for (forvar829 = (1'h0); (forvar829 < (3'h4)); forvar829 = (forvar829 + (1'h1)))
                begin
                  reg830 = $unsigned($unsigned((&(reg816 ?
                      (!reg817) : "mQ8mW74gf"))));
                  reg831 = reg808[(4'h8):(3'h6)];
                  reg832 <= {$signed($signed(reg789))};
                end
              reg833 <= (^{("zuuf0ztkShQZRY1axE" ?
                      reg822 : (^~(reg813 - reg811)))});
            end
          reg834 = $unsigned(reg801[(2'h3):(1'h0)]);
          reg835 <= ((7'h4b) ^ $unsigned((^~forvar810)));
        end
      reg836 = $signed(wire780[(2'h2):(2'h2)]);
      reg837 <= $signed(wire782[(4'h8):(3'h4)]);
      reg838 <= (~^{(reg808[(3'h5):(1'h1)] << ($unsigned((8'hb8)) * "Pyeb06Z59so7BN"))});
    end
  assign wire839 = (reg795[(1'h0):(1'h0)] << wire782[(3'h7):(3'h5)]);
  always
    @(posedge clk) begin
      reg840 <= reg819;
      reg841 = (^(reg801 ? $signed("nY0R1UJv4T6RpL5") : (|wire783)));
      for (forvar842 = (1'h0); (forvar842 < (2'h3)); forvar842 = (forvar842 + (1'h1)))
        begin
          for (forvar843 = (1'h0); (forvar843 < (3'h4)); forvar843 = (forvar843 + (1'h1)))
            begin
              reg844 <= ((reg815 ?
                      "Edf9UUZbr78" : $signed(($signed((7'h42)) | (8'hbb)))) ?
                  (^(((reg831 ~^ forvar821) >= (&forvar809)) && reg787[(3'h5):(1'h0)])) : wire792);
              reg845 <= $unsigned($signed({{(reg827 <<< reg803),
                      {reg834, reg816}}}));
              reg846 <= $signed(wire790);
              reg847 <= reg814[(2'h3):(2'h3)];
              for (forvar848 = (1'h0); (forvar848 < (3'h5)); forvar848 = (forvar848 + (1'h1)))
                begin
                  reg849 = $unsigned(((forvar843[(1'h1):(1'h0)] ?
                      (|$signed(reg814)) : wire780) > wire783[(1'h0):(1'h0)]));
                  reg850 = "JlwNRITg4M6PovcU4B";
                  reg851 <= $unsigned((wire784[(2'h2):(1'h0)] ?
                      reg796 : ((-reg799) || ((reg795 ?
                          reg807 : reg796) <= (~|reg844)))));
                  reg852 <= $signed({"NqZMWL"});
                end
            end
          reg853 <= (((($unsigned(reg832) ?
              $unsigned(wire785) : $unsigned(reg824)) >> (8'hac)) ^~ ("AGb48qCKRoP3H1Jakr2p" && reg806)) + (((8'hae) ?
                  $signed(forvar828[(2'h2):(2'h2)]) : ("dXWHJU6LryvPo6MzW" <= forvar843)) ?
              {(reg794[(3'h4):(2'h2)] >>> reg841[(3'h7):(2'h2)]),
                  ($unsigned(reg800) >>> reg808[(3'h5):(1'h0)])} : reg797[(2'h2):(1'h0)]));
        end
      reg854 <= forvar810;
      reg855 <= reg811;
      reg856 <= $signed($unsigned(({$signed(reg847)} ?
          (7'h45) : "rSiazqGMO7a20NSp")));
    end
  always
    @(posedge clk) begin
      reg857 <= $unsigned((wire784[(2'h3):(2'h3)] ^~ (~$unsigned($unsigned(reg809)))));
      reg858 <= $unsigned((~(!forvar828)));
      for (forvar859 = (1'h0); (forvar859 < (2'h3)); forvar859 = (forvar859 + (1'h1)))
        begin
          reg860 <= $signed($unsigned($signed($signed(reg851[(1'h0):(1'h0)]))));
          if (wire792[(3'h7):(2'h2)])
            begin
              reg861 <= $unsigned($signed($unsigned($unsigned((reg855 ?
                  wire783 : (8'ha9))))));
              if (forvar809[(1'h0):(1'h0)])
                begin
                  reg862 <= $unsigned((reg845 ?
                      (forvar828 ?
                          {wire793[(4'h9):(3'h7)],
                              (reg830 << reg835)} : (reg789 ?
                              reg795[(2'h2):(1'h0)] : (-(8'ha0)))) : ((!(reg804 ?
                              reg858 : reg832)) ?
                          $signed((reg835 ?
                              reg854 : forvar810)) : $unsigned({forvar821,
                              (7'h4c)}))));
                end
              else
                begin
                  reg862 = "XlHLoR41u3rFqn";
                  reg863 = "DncVylp8Ak6A";
                  reg864 <= (~^(forvar810[(3'h7):(2'h2)] ?
                      ((&(reg815 ?
                          (8'ha5) : reg814)) << reg816[(1'h0):(1'h0)]) : {"A0HV40",
                          (reg826[(1'h1):(1'h1)] ?
                              (~^forvar821) : $signed(reg786))}));
                  reg865 <= (^~wire784);
                  reg866 = (8'h9e);
                  reg867 = reg820[(5'h14):(5'h14)];
                end
            end
          else
            begin
              reg861 <= (|$unsigned((($unsigned(forvar829) ?
                  $signed(reg866) : reg810[(1'h1):(1'h1)]) <= (reg846 ?
                  "Ai" : $signed(reg836)))));
              reg862 <= (!(-$signed(($unsigned(reg810) & "Ze"))));
              reg863 <= (~|"xS2B1gIU");
              reg864 <= ($signed("7ldblh") ? "bFOKQzWgglqXiDisOd95sOGaD" : "b");
            end
          reg868 <= {(|(8'h9f)),
              $unsigned(($signed(reg808[(4'ha):(4'h8)]) >> $signed((reg798 ?
                  reg820 : reg808))))};
        end
      reg869 <= reg816[(2'h2):(1'h0)];
    end
  always
    @(posedge clk) begin
      for (forvar870 = (1'h0); (forvar870 < (1'h1)); forvar870 = (forvar870 + (1'h1)))
        begin
          for (forvar871 = (1'h0); (forvar871 < (2'h2)); forvar871 = (forvar871 + (1'h1)))
            begin
              reg872 <= $unsigned("542ght5HyiUCq");
              for (forvar873 = (1'h0); (forvar873 < (1'h1)); forvar873 = (forvar873 + (1'h1)))
                begin
                  reg874 <= (+"SpL");
                  reg875 = "PCL5ag23klwaR";
                  reg876 <= $signed(forvar807);
                  reg877 = "roNAvdC";
                end
              for (forvar878 = (1'h0); (forvar878 < (3'h4)); forvar878 = (forvar878 + (1'h1)))
                begin
                  reg879 <= $unsigned($unsigned($signed(((reg854 ?
                      reg864 : forvar828) ~^ (reg838 <<< (8'hac))))));
                  reg880 <= (-$unsigned("BDveDPt9TdoFLnQfCLc8ow2"));
                  reg881 <= $signed($signed(((!(wire783 ? reg816 : reg834)) ?
                      ((wire781 ? reg868 : reg789) - (reg812 ?
                          reg858 : reg835)) : "McX68kCC27zIEzh")));
                  reg882 <= {(wire791[(1'h0):(1'h0)] ?
                          "" : ((^reg854[(3'h5):(1'h0)]) && "BLPDWgvVoYrN1T98HEbIKK"))};
                end
            end
          reg883 = $unsigned("WlEsd3tbP");
          reg884 <= $unsigned($signed((("uPMuiMNs6c89gqOsZacz6S5" ?
              $signed((8'hb5)) : (reg786 > forvar843)) - "st6kZVfb9TUDSSmsZCu6t")));
        end
      reg885 = $unsigned("Dd1k2mzNZGFVCG");
      reg886 <= {$unsigned((7'h48)), $signed((~"2fvNL1TOxHPnSNf"))};
      reg887 <= {$unsigned(reg836[(5'h10):(1'h1)]),
          ("GR" ? reg856[(1'h0):(1'h0)] : reg813[(3'h4):(1'h1)])};
      reg888 <= forvar848;
    end
  assign wire889 = (reg856[(1'h0):(1'h0)] << (~&reg801[(2'h2):(2'h2)]));
  always
    @(posedge clk) begin
      reg890 <= $unsigned($signed($unsigned($unsigned(reg852[(2'h2):(2'h2)]))));
      reg891 <= ((!(~^(|reg832[(1'h1):(1'h0)]))) ?
          ($signed($unsigned(((8'ha8) <<< forvar870))) || (+$unsigned(wire782))) : (~$signed({reg823[(5'h17):(4'h8)]})));
      reg892 <= $unsigned({reg798, (~&"V0KBPKVO6LD34")});
      reg893 <= (($unsigned(((reg860 ? reg838 : forvar842) | (reg888 ?
                  wire889 : (8'ha7)))) ?
              $signed($signed(reg837)) : $signed({$unsigned(reg816),
                  (reg890 <= reg822)})) ?
          $unsigned(((reg881 >> $signed((8'ha7))) ^ (~(reg813 ?
              (8'ha8) : reg882)))) : (!reg806[(3'h7):(3'h6)]));
      reg894 = ("dtQEkuTbTzWzM0HiG4wnEmT3" ?
          $signed(reg857[(4'hb):(3'h4)]) : $unsigned(((reg819 ?
                  (reg837 >= wire780) : "0YZ") ?
              ({forvar828,
                  reg846} <= "FWSFuvkJxy3C") : $unsigned("iVWnLKu6kyB6"))));
    end
  always
    @(posedge clk) begin
      reg895 <= reg865[(4'hb):(3'h7)];
      for (forvar896 = (1'h0); (forvar896 < (2'h3)); forvar896 = (forvar896 + (1'h1)))
        begin
          reg897 <= $signed({($unsigned((forvar842 ?
                  forvar821 : wire780)) <= reg869),
              (wire791 <<< $signed($signed((8'ha7))))});
        end
      reg898 <= $signed($signed(reg832[(4'h8):(1'h0)]));
      for (forvar899 = (1'h0); (forvar899 < (3'h5)); forvar899 = (forvar899 + (1'h1)))
        begin
          reg900 <= ($unsigned($unsigned(reg809[(4'h8):(2'h3)])) ?
              reg810[(3'h7):(3'h5)] : "rAABh8S3nq6wBxaswgI");
          reg901 <= $signed($signed(wire781[(3'h7):(1'h1)]));
          reg902 = reg812[(3'h5):(2'h3)];
          reg903 <= (reg797 ^ reg832[(3'h7):(3'h4)]);
          reg904 <= {reg890,
              (&(($signed(wire839) >>> $signed((8'haa))) | (reg897 >= "hEysHLUyVQodDLA")))};
        end
    end
  always
    @(posedge clk) begin
      reg905 = "mhsn";
      for (forvar906 = (1'h0); (forvar906 < (3'h5)); forvar906 = (forvar906 + (1'h1)))
        begin
          for (forvar907 = (1'h0); (forvar907 < (1'h0)); forvar907 = (forvar907 + (1'h1)))
            begin
              reg908 <= (|$unsigned(((7'h4e) != ("kkZtI" | $unsigned(reg834)))));
              reg909 <= (reg809[(2'h2):(1'h1)] ?
                  (forvar810[(4'hb):(4'hb)] ?
                      reg812[(3'h4):(3'h4)] : $signed(reg867[(2'h2):(2'h2)])) : {((reg867 ?
                              (reg789 ~^ (8'hb0)) : "tN") ?
                          reg884[(3'h5):(1'h0)] : reg797),
                      (|$signed((reg822 != reg849)))});
              reg910 = $unsigned((&reg865[(3'h4):(2'h2)]));
              reg911 <= $unsigned({reg879,
                  (forvar829 && ((reg886 ? reg879 : reg823) >= (~forvar899)))});
              reg912 <= $unsigned("y9TGVp");
            end
          reg913 <= $signed(reg852);
          for (forvar914 = (1'h0); (forvar914 < (3'h4)); forvar914 = (forvar914 + (1'h1)))
            begin
              reg915 <= (+$signed("w4haPx5n1tAEqYOid2"));
              for (forvar916 = (1'h0); (forvar916 < (1'h1)); forvar916 = (forvar916 + (1'h1)))
                begin
                  reg917 <= $unsigned(((reg808 <= forvar899[(3'h6):(3'h4)]) ?
                      reg834[(2'h2):(1'h1)] : $signed(((~reg872) && (reg851 ^ reg876)))));
                  reg918 <= {(7'h47),
                      ({$unsigned({reg857, reg798}),
                          reg800} >>> reg819[(4'ha):(4'h8)])};
                  reg919 <= $signed($signed(($signed((-reg815)) != ("lNTq3TDt" - reg895))));
                  reg920 <= $signed($signed(reg796[(5'h11):(4'h8)]));
                end
            end
          reg921 <= reg897;
          for (forvar922 = (1'h0); (forvar922 < (1'h1)); forvar922 = (forvar922 + (1'h1)))
            begin
              reg923 <= (reg801[(2'h3):(2'h3)] < ({($unsigned(reg820) < "")} ?
                  (&{reg854[(2'h3):(2'h2)],
                      (reg920 ? reg920 : (7'h44))}) : {{(reg788 - (7'h4e)),
                          (!reg864)}}));
              reg924 <= {(reg921[(2'h3):(2'h3)] ?
                      "tCOAZf3ddr4o4r" : $unsigned((~|$unsigned(reg798))))};
              reg925 <= wire785[(3'h5):(2'h3)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg926 = "2zU1EUSayZ1sIJk72gqQP1";
      for (forvar927 = (1'h0); (forvar927 < (3'h5)); forvar927 = (forvar927 + (1'h1)))
        begin
          reg928 <= ((^~$unsigned("ILqcGTsIZL")) < {($unsigned($unsigned(reg812)) < (8'hbf)),
              reg909});
          reg929 <= reg879[(1'h0):(1'h0)];
          reg930 <= ((reg909[(3'h7):(1'h1)] ? "oWdalYHqkMPJlRfVY7u" : reg866) ?
              (~("qFC4gg3m" ?
                  $signed($signed(reg846)) : reg826)) : reg810[(3'h7):(3'h6)]);
          for (forvar931 = (1'h0); (forvar931 < (1'h0)); forvar931 = (forvar931 + (1'h1)))
            begin
              reg932 <= (~(($signed((forvar829 ? wire780 : reg804)) ?
                  forvar896[(5'h12):(2'h3)] : $unsigned(reg894)) - "KyeLoIvJ"));
              reg933 = ($signed((wire793 && $unsigned((+reg840)))) <<< reg905);
              reg934 <= ("Pol4DCOqM6JJfnWqphyhX" + $unsigned({"", "yI58PQte"}));
            end
          reg935 <= reg851;
          for (forvar936 = (1'h0); (forvar936 < (1'h0)); forvar936 = (forvar936 + (1'h1)))
            begin
              reg937 <= forvar842;
              reg938 <= $unsigned($unsigned($signed($signed((-reg844)))));
              reg939 <= ((((reg892 >>> (reg865 == reg788)) + "fX7LL2Q6X0QNZ7GqfRCpW") * (reg913[(3'h4):(2'h2)] ?
                      ($unsigned(reg932) ?
                          $unsigned(reg832) : reg802[(4'hd):(4'h9)]) : $signed($signed(reg888)))) ?
                  forvar922[(3'h6):(1'h1)] : reg924);
              reg940 = ((^~(reg929[(4'hf):(3'h4)] ?
                  $signed(reg884[(3'h5):(1'h1)]) : ((reg853 | reg887) ?
                      {reg884, reg830} : reg805))) && {("0tNdtOuzmvyuuTdiQxh3" ?
                      $signed($signed(reg937)) : ($signed(reg851) ?
                          reg808[(2'h3):(1'h1)] : (forvar878 ?
                              reg860 : reg809))),
                  (7'h42)});
              reg941 = ((|forvar916[(5'h13):(1'h1)]) ?
                  $unsigned(forvar843) : (8'hbb));
              for (forvar942 = (1'h0); (forvar942 < (1'h0)); forvar942 = (forvar942 + (1'h1)))
                begin
                  reg943 = $signed("6vYkg");
                end
            end
        end
      reg944 = reg883[(3'h7):(3'h4)];
      for (forvar945 = (1'h0); (forvar945 < (2'h2)); forvar945 = (forvar945 + (1'h1)))
        begin
          reg946 <= "Zckce";
          reg947 = (~^reg807[(3'h4):(2'h3)]);
          reg948 <= "";
        end
      reg949 <= {{"YwOLPzmYLL77oH"}, "F0A"};
      reg950 <= "tWKIR";
    end
  always
    @(posedge clk) begin
      reg951 <= ((+$signed(reg831)) ?
          {$unsigned($signed(forvar907[(4'h9):(3'h5)])),
              "fLY4z7o1e3goew8dHPlAmsv"} : {{("MzyitPRxUP1aESV7YmMB" ?
                      (~^reg937) : $unsigned(reg824)),
                  ((reg840 == forvar843) ? reg881 : $signed(wire839))},
              (({reg933} <<< "baElZUEaqYow4CWviCM6Fm") > reg814)});
      reg952 <= reg934;
      reg953 = $signed($signed((~|$unsigned(reg800[(4'ha):(2'h2)]))));
      reg954 <= ((&"nk3x4O39Ux83") >= $unsigned($signed("lm9Iq4")));
      for (forvar955 = (1'h0); (forvar955 < (2'h3)); forvar955 = (forvar955 + (1'h1)))
        begin
          reg956 <= "x2QGy9u1Pik7A";
          reg957 <= reg854;
          reg958 <= $unsigned(reg801[(4'he):(3'h5)]);
          reg959 <= reg796;
          reg960 = $unsigned(reg855[(3'h4):(2'h2)]);
        end
      reg961 <= $signed(reg949);
    end
  always
    @(posedge clk) begin
      reg962 <= reg841;
      reg963 <= wire793[(4'hc):(3'h6)];
      for (forvar964 = (1'h0); (forvar964 < (3'h5)); forvar964 = (forvar964 + (1'h1)))
        begin
          for (forvar965 = (1'h0); (forvar965 < (2'h2)); forvar965 = (forvar965 + (1'h1)))
            begin
              reg966 <= ($unsigned(reg857) ?
                  ((reg904[(2'h3):(1'h1)] > "548QnymDDzOwZ4s5") ?
                      $unsigned((reg822 || "1X49kTDobdfaf6")) : reg903[(2'h3):(1'h1)]) : "R3Jg55y");
            end
          reg967 <= ($signed(forvar922[(3'h4):(2'h3)]) && (($signed(reg962[(1'h0):(1'h0)]) ?
              "Rdh9CcLACMxy" : ((+reg882) ?
                  (+(8'hb0)) : $unsigned(forvar936))) > $signed((forvar842 ?
              $unsigned(reg811) : (+reg818)))));
          reg968 <= $signed("Oc9tp99bIVkdPDLB6gqw6LO");
          for (forvar969 = (1'h0); (forvar969 < (1'h1)); forvar969 = (forvar969 + (1'h1)))
            begin
              reg970 = (reg798 >> (^~$unsigned(reg910)));
            end
          for (forvar971 = (1'h0); (forvar971 < (3'h4)); forvar971 = (forvar971 + (1'h1)))
            begin
              reg972 <= forvar931[(3'h6):(3'h4)];
              for (forvar973 = (1'h0); (forvar973 < (3'h5)); forvar973 = (forvar973 + (1'h1)))
                begin
                  reg974 <= reg837;
                end
              reg975 = ((reg853 ? "f9" : "AwiVOgvCcR5I") ?
                  $unsigned(reg912[(4'hc):(3'h5)]) : reg788[(1'h0):(1'h0)]);
              reg976 <= $signed((|forvar859[(1'h1):(1'h1)]));
            end
          reg977 <= reg948[(3'h5):(3'h5)];
        end
      reg978 <= "I8S7SbbrGX";
    end
  always
    @(posedge clk) begin
      reg979 = reg786;
      reg980 <= reg849[(5'h11):(4'h9)];
      reg981 <= $signed((("i0k7PPE" * {(+(8'hb4)), wire790}) >>> "iIrxNCiZ"));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module560  (y, clk, wire565, wire564, wire563, wire562, wire561);
  output wire [(32'ha33):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire565;
  input wire signed [(5'h19):(1'h0)] wire564;
  input wire signed [(5'h16):(1'h0)] wire563;
  input wire [(3'h5):(1'h0)] wire562;
  input wire [(5'h18):(1'h0)] wire561;
  reg [(4'h9):(1'h0)] reg749 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg748 = (1'h0);
  reg [(4'hd):(1'h0)] reg747 = (1'h0);
  reg [(4'h9):(1'h0)] reg746 = (1'h0);
  reg [(3'h6):(1'h0)] reg745 = (1'h0);
  reg [(5'h12):(1'h0)] reg744 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar743 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg742 = (1'h0);
  reg [(4'hc):(1'h0)] reg741 = (1'h0);
  reg [(4'ha):(1'h0)] reg740 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar739 = (1'h0);
  reg [(4'hd):(1'h0)] reg738 = (1'h0);
  reg [(2'h2):(1'h0)] reg737 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg736 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg735 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg734 = (1'h0);
  reg [(2'h3):(1'h0)] reg733 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar732 = (1'h0);
  reg [(4'hf):(1'h0)] forvar731 = (1'h0);
  reg [(5'h17):(1'h0)] reg730 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg729 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg728 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg727 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar726 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg725 = (1'h0);
  reg [(4'hb):(1'h0)] reg724 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar723 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg722 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg721 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg720 = (1'h0);
  reg [(3'h6):(1'h0)] reg719 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg718 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg717 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg716 = (1'h0);
  reg [(5'h15):(1'h0)] reg715 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg714 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar713 = (1'h0);
  reg [(5'h13):(1'h0)] reg712 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar711 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg710 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg709 = (1'h0);
  reg [(5'h14):(1'h0)] reg708 = (1'h0);
  reg [(5'h15):(1'h0)] forvar707 = (1'h0);
  wire [(3'h7):(1'h0)] wire706;
  wire signed [(4'hb):(1'h0)] wire705;
  reg signed [(5'h13):(1'h0)] reg704 = (1'h0);
  reg [(5'h16):(1'h0)] reg703 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg702 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg701 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg700 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg699 = (1'h0);
  reg [(5'h10):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg697 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg696 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire695;
  reg [(5'h16):(1'h0)] reg694 = (1'h0);
  reg [(5'h12):(1'h0)] reg693 = (1'h0);
  reg [(5'h11):(1'h0)] reg692 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar691 = (1'h0);
  reg [(5'h13):(1'h0)] forvar690 = (1'h0);
  reg signed [(4'he):(1'h0)] reg689 = (1'h0);
  reg [(5'h19):(1'h0)] reg688 = (1'h0);
  reg [(5'h17):(1'h0)] reg687 = (1'h0);
  reg [(4'hc):(1'h0)] forvar683 = (1'h0);
  reg [(5'h16):(1'h0)] reg686 = (1'h0);
  reg [(4'hc):(1'h0)] reg685 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg684 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg681 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg683 = (1'h0);
  reg [(5'h17):(1'h0)] reg682 = (1'h0);
  reg [(4'h9):(1'h0)] forvar681 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg680 = (1'h0);
  reg [(4'hc):(1'h0)] reg679 = (1'h0);
  reg [(5'h16):(1'h0)] reg678 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire677;
  reg signed [(4'hd):(1'h0)] reg676 = (1'h0);
  wire signed [(5'h18):(1'h0)] wire675;
  reg signed [(4'hb):(1'h0)] reg674 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg673 = (1'h0);
  reg [(5'h1a):(1'h0)] reg672 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg671 = (1'h0);
  reg [(4'hd):(1'h0)] reg670 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg669 = (1'h0);
  reg [(4'ha):(1'h0)] reg668 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg667 = (1'h0);
  reg [(5'h12):(1'h0)] reg666 = (1'h0);
  reg [(5'h10):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg664 = (1'h0);
  reg [(5'h1a):(1'h0)] reg663 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar662 = (1'h0);
  reg [(4'hc):(1'h0)] reg661 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar660 = (1'h0);
  reg [(5'h1a):(1'h0)] reg659 = (1'h0);
  reg [(5'h10):(1'h0)] forvar658 = (1'h0);
  reg [(2'h3):(1'h0)] reg657 = (1'h0);
  reg [(4'he):(1'h0)] reg656 = (1'h0);
  reg [(4'he):(1'h0)] reg655 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar654 = (1'h0);
  wire [(3'h5):(1'h0)] wire653;
  wire signed [(4'h9):(1'h0)] wire652;
  reg signed [(4'h8):(1'h0)] reg651 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg650 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg649 = (1'h0);
  reg [(5'h11):(1'h0)] reg648 = (1'h0);
  reg [(5'h15):(1'h0)] reg647 = (1'h0);
  reg [(2'h2):(1'h0)] reg646 = (1'h0);
  reg [(5'h1a):(1'h0)] reg645 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg644 = (1'h0);
  reg [(2'h3):(1'h0)] forvar643 = (1'h0);
  reg [(5'h19):(1'h0)] forvar642 = (1'h0);
  reg [(4'h8):(1'h0)] reg641 = (1'h0);
  reg [(3'h6):(1'h0)] reg640 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg639 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg638 = (1'h0);
  reg [(4'h8):(1'h0)] reg637 = (1'h0);
  reg [(4'hb):(1'h0)] forvar636 = (1'h0);
  reg [(4'h8):(1'h0)] reg635 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg634 = (1'h0);
  reg [(4'hd):(1'h0)] reg633 = (1'h0);
  reg [(5'h11):(1'h0)] reg632 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg631 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg630 = (1'h0);
  reg [(4'hf):(1'h0)] reg629 = (1'h0);
  reg [(3'h4):(1'h0)] reg628 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg627 = (1'h0);
  reg [(4'ha):(1'h0)] reg626 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg623 = (1'h0);
  reg [(4'hd):(1'h0)] reg622 = (1'h0);
  reg [(3'h6):(1'h0)] forvar621 = (1'h0);
  reg [(4'hd):(1'h0)] reg620 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg619 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg618 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg617 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg616 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar615 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg614 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg613 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg612 = (1'h0);
  reg [(4'hf):(1'h0)] reg611 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg610 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg609 = (1'h0);
  reg [(4'hb):(1'h0)] forvar608 = (1'h0);
  reg [(3'h7):(1'h0)] reg607 = (1'h0);
  reg [(2'h2):(1'h0)] reg606 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg605 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg604 = (1'h0);
  wire [(3'h6):(1'h0)] wire603;
  reg signed [(5'h1a):(1'h0)] reg602 = (1'h0);
  reg [(4'h9):(1'h0)] reg601 = (1'h0);
  reg [(5'h18):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg599 = (1'h0);
  reg [(5'h16):(1'h0)] reg598 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg597 = (1'h0);
  reg [(5'h19):(1'h0)] reg596 = (1'h0);
  reg [(4'hf):(1'h0)] reg595 = (1'h0);
  reg [(5'h18):(1'h0)] forvar594 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg593 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar592 = (1'h0);
  reg [(4'hb):(1'h0)] reg591 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg590 = (1'h0);
  reg [(5'h11):(1'h0)] reg589 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar588 = (1'h0);
  reg [(4'hc):(1'h0)] reg587 = (1'h0);
  reg [(4'hc):(1'h0)] reg586 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg585 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg584 = (1'h0);
  reg [(5'h1a):(1'h0)] reg583 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg581 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg580 = (1'h0);
  reg [(5'h13):(1'h0)] reg579 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg578 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg577 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg576 = (1'h0);
  reg [(5'h16):(1'h0)] forvar575 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg574 = (1'h0);
  reg [(3'h4):(1'h0)] reg573 = (1'h0);
  reg [(3'h5):(1'h0)] forvar572 = (1'h0);
  reg [(5'h12):(1'h0)] reg571 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg570 = (1'h0);
  reg [(5'h11):(1'h0)] reg569 = (1'h0);
  reg [(5'h16):(1'h0)] forvar568 = (1'h0);
  reg [(4'hb):(1'h0)] forvar567 = (1'h0);
  reg [(4'h9):(1'h0)] reg566 = (1'h0);
  assign y = {reg749,
                 reg748,
                 reg747,
                 reg746,
                 reg745,
                 reg744,
                 forvar743,
                 reg742,
                 reg741,
                 reg740,
                 forvar739,
                 reg738,
                 reg737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 forvar732,
                 forvar731,
                 reg730,
                 reg729,
                 reg728,
                 reg727,
                 forvar726,
                 reg725,
                 reg724,
                 forvar723,
                 reg722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 forvar713,
                 reg712,
                 forvar711,
                 reg710,
                 reg709,
                 reg708,
                 forvar707,
                 wire706,
                 wire705,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 reg699,
                 reg698,
                 reg697,
                 reg696,
                 wire695,
                 reg694,
                 reg693,
                 reg692,
                 forvar691,
                 forvar690,
                 reg689,
                 reg688,
                 reg687,
                 forvar683,
                 reg686,
                 reg685,
                 reg684,
                 reg681,
                 reg683,
                 reg682,
                 forvar681,
                 reg680,
                 reg679,
                 reg678,
                 wire677,
                 reg676,
                 wire675,
                 reg674,
                 reg673,
                 reg672,
                 reg671,
                 reg670,
                 reg669,
                 reg668,
                 reg667,
                 reg666,
                 reg665,
                 reg664,
                 reg663,
                 forvar662,
                 reg661,
                 forvar660,
                 reg659,
                 forvar658,
                 reg657,
                 reg656,
                 reg655,
                 forvar654,
                 wire653,
                 wire652,
                 reg651,
                 reg650,
                 reg649,
                 reg648,
                 reg647,
                 reg646,
                 reg645,
                 reg644,
                 forvar643,
                 forvar642,
                 reg641,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 forvar636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 forvar621,
                 reg620,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 forvar615,
                 reg614,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 reg609,
                 forvar608,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 wire603,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 forvar594,
                 reg593,
                 forvar592,
                 reg591,
                 reg590,
                 reg589,
                 forvar588,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 reg579,
                 reg578,
                 reg577,
                 reg576,
                 forvar575,
                 reg574,
                 reg573,
                 forvar572,
                 reg571,
                 reg570,
                 reg569,
                 forvar568,
                 forvar567,
                 reg566,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg566 <= (wire562[(1'h0):(1'h0)] ?
          wire565 : $unsigned((wire564[(5'h11):(5'h10)] > {$signed(wire564),
              "P7XSXDE4Oriu7EZKA7NBRy"})));
      for (forvar567 = (1'h0); (forvar567 < (3'h5)); forvar567 = (forvar567 + (1'h1)))
        begin
          for (forvar568 = (1'h0); (forvar568 < (1'h1)); forvar568 = (forvar568 + (1'h1)))
            begin
              reg569 <= $unsigned($unsigned((7'h4b)));
              reg570 <= ($signed($signed(wire561[(4'he):(4'hb)])) | "6mJlpwahAn6mT");
            end
        end
      reg571 <= (wire561[(4'h8):(3'h7)] & "wvoMCErgIaT9M7KSID");
      for (forvar572 = (1'h0); (forvar572 < (2'h2)); forvar572 = (forvar572 + (1'h1)))
        begin
          reg573 <= {$signed($signed("vO1qIeg3y"))};
          reg574 <= (((~($signed((8'hb6)) + {reg569})) ?
              (-"0Aca8Afezfq5mWgg") : wire565[(3'h6):(3'h4)]) | (8'haa));
          for (forvar575 = (1'h0); (forvar575 < (2'h3)); forvar575 = (forvar575 + (1'h1)))
            begin
              if ({$signed("JaqXbPg8g"),
                  $signed(("QNmlUzy" ~^ ((forvar572 ?
                      wire565 : wire564) <<< $unsigned(reg574))))})
                begin
                  reg576 <= $signed((|$unsigned(((reg574 + reg571) ?
                      wire565[(3'h4):(1'h1)] : (reg571 ~^ wire565)))));
                  reg577 <= $signed(forvar572);
                  reg578 = $signed(forvar567);
                  reg579 <= ({(((+wire564) ~^ $signed(reg569)) | "k12p")} ?
                      (+forvar575[(4'hd):(3'h4)]) : reg571[(3'h6):(1'h0)]);
                  reg580 <= (!"WU7R8yHOMa4VSqiYHo0D7bhcs");
                  reg581 <= $signed("FpVtw");
                end
              else
                begin
                  reg576 <= (reg566 ? reg577 : "TGfEc8RB3");
                end
              reg582 <= ((|(8'had)) >> "rLmLK0apg83DxA50HdHDa");
              reg583 = (8'haf);
              reg584 = ("stoybM8CyI8tLS8i3o" > {forvar575});
            end
        end
    end
  always
    @(posedge clk) begin
      reg585 = "woxe3vBJ35muuEhbKJ";
      reg586 <= $signed((~&{reg571, "hBfXFteGx4GQixqWBJU"}));
      reg587 <= "2a1CvPNIZOMMcCDc1";
      for (forvar588 = (1'h0); (forvar588 < (2'h3)); forvar588 = (forvar588 + (1'h1)))
        begin
          reg589 <= wire564[(4'hb):(2'h3)];
          reg590 <= forvar572[(2'h2):(2'h2)];
        end
    end
  always
    @(posedge clk) begin
      reg591 <= "fZZb";
      for (forvar592 = (1'h0); (forvar592 < (2'h2)); forvar592 = (forvar592 + (1'h1)))
        begin
          reg593 = reg582[(2'h2):(1'h1)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar594 = (1'h0); (forvar594 < (3'h5)); forvar594 = (forvar594 + (1'h1)))
        begin
          reg595 = {($signed($unsigned((reg579 < reg593))) ?
                  $signed((|$signed(reg587))) : ($unsigned((^wire563)) | $signed(reg583[(4'h9):(4'h9)]))),
              (8'hb3)};
          reg596 <= $signed((reg569[(4'h8):(3'h4)] ?
              "18mi1QztYegeRoD" : $signed(((8'ha6) ? (^wire565) : reg573))));
          reg597 <= wire562[(3'h5):(3'h5)];
          reg598 <= reg591;
          reg599 <= (reg578 || "hTV2y6u6imAGgCI");
        end
      reg600 <= $unsigned((+{"ZM"}));
      reg601 <= (~^(!((~^forvar594) | $signed(forvar572[(2'h3):(2'h3)]))));
      reg602 <= ($unsigned(reg571[(2'h2):(2'h2)]) < reg587);
    end
  assign wire603 = reg576[(4'hb):(3'h6)];
  always
    @(posedge clk) begin
      reg604 <= reg570[(4'hd):(4'hb)];
      reg605 = reg574;
      reg606 <= {(8'hb9), (~reg604)};
      reg607 <= $signed($signed(reg597));
      for (forvar608 = (1'h0); (forvar608 < (2'h3)); forvar608 = (forvar608 + (1'h1)))
        begin
          reg609 <= reg597;
          reg610 <= ($unsigned(reg571[(4'hc):(3'h7)]) ?
              (~|((^wire564) ?
                  (reg570 ?
                      (&forvar575) : "N8vv9P1uJZFbn") : $unsigned(reg600[(5'h11):(4'hc)]))) : (-(^$signed((forvar588 ?
                  reg591 : reg609)))));
          reg611 <= (+(&reg585[(1'h1):(1'h1)]));
          reg612 <= reg598;
          if ($unsigned({(~(^$signed(reg586))), "4T"}))
            begin
              reg613 <= ($unsigned(reg574) ^ $unsigned({"8bb4TvT", "gBKSL"}));
            end
          else
            begin
              reg613 = wire562;
              reg614 <= $signed($unsigned("mE"));
              for (forvar615 = (1'h0); (forvar615 < (1'h0)); forvar615 = (forvar615 + (1'h1)))
                begin
                  reg616 <= "hp1ADiqRTEfGK";
                  reg617 = (wire564 || ("UeeawwGvhb7DcN1EBvJR" ?
                      reg586[(3'h4):(1'h1)] : (^~"gp4v")));
                  reg618 = reg577;
                  reg619 = $unsigned($unsigned({(reg595[(4'h8):(3'h6)] - {forvar568}),
                      (^"9Xgk10syLqVvIwE0FJbJ")}));
                end
            end
        end
    end
  always
    @(posedge clk) begin
      reg620 = wire561;
      for (forvar621 = (1'h0); (forvar621 < (3'h5)); forvar621 = (forvar621 + (1'h1)))
        begin
          reg622 <= reg574[(2'h3):(2'h2)];
          reg623 <= (+("gM4hJgAyE1XAmmSPV" + (~^$unsigned((forvar588 ?
              reg569 : wire603)))));
          reg624 <= "L0OcCKUpB7UpmTHsR7RDT3wA0";
          reg625 <= reg584;
        end
      reg626 <= $signed(((^~reg576) > reg606[(1'h1):(1'h0)]));
      reg627 <= $unsigned(forvar567[(3'h4):(3'h4)]);
    end
  always
    @(posedge clk) begin
      reg628 <= {({(8'hb9)} ?
              (!((wire603 | forvar572) >>> "dUrbAnPbcb")) : reg614[(5'h18):(3'h5)])};
      reg629 = reg574[(5'h10):(4'ha)];
    end
  always
    @(posedge clk) begin
      reg630 = reg578;
      reg631 <= reg576;
      reg632 <= (reg579[(5'h13):(4'hb)] - wire561[(5'h17):(5'h14)]);
      reg633 <= (forvar572[(1'h0):(1'h0)] >>> "wXHZ7M4");
    end
  always
    @(posedge clk) begin
      reg634 = reg631;
      reg635 <= $unsigned((^~"d"));
      for (forvar636 = (1'h0); (forvar636 < (3'h5)); forvar636 = (forvar636 + (1'h1)))
        begin
          reg637 = (((&"t") ?
              $unsigned(reg600[(3'h7):(3'h7)]) : "Qb") + reg578[(2'h2):(2'h2)]);
          reg638 <= "gG3bxbesmd";
          reg639 <= wire603[(3'h6):(3'h5)];
          reg640 <= $signed("nrJ1kb");
          reg641 <= ("Mz4aIZ7MlOYv" << $signed($signed(reg619[(4'h8):(4'h8)])));
          for (forvar642 = (1'h0); (forvar642 < (2'h2)); forvar642 = (forvar642 + (1'h1)))
            begin
              for (forvar643 = (1'h0); (forvar643 < (3'h5)); forvar643 = (forvar643 + (1'h1)))
                begin
                  reg644 <= wire603;
                  reg645 <= reg577[(2'h2):(1'h1)];
                  reg646 <= ({$signed($unsigned(reg610[(1'h0):(1'h0)]))} ?
                      (("IR3m3GrLLJuwiA" + (reg576 || forvar594[(3'h5):(2'h3)])) ?
                          reg599 : ($signed($unsigned(reg611)) ?
                              reg639 : $signed(((8'hb3) ^ wire563)))) : "2PQZVt");
                  reg647 <= (7'h43);
                  reg648 <= reg630;
                end
              reg649 <= $signed("SkNOGOTlpzzen");
              reg650 <= reg626[(3'h5):(1'h0)];
              reg651 <= forvar615[(2'h3):(2'h3)];
            end
        end
    end
  assign wire652 = reg576;
  assign wire653 = reg591[(4'ha):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar654 = (1'h0); (forvar654 < (2'h3)); forvar654 = (forvar654 + (1'h1)))
        begin
          reg655 <= (reg620[(4'hc):(3'h4)] ? "I7" : "tw83icHf");
          reg656 <= $unsigned(reg646[(1'h0):(1'h0)]);
        end
      reg657 <= $unsigned(reg598);
      for (forvar658 = (1'h0); (forvar658 < (2'h2)); forvar658 = (forvar658 + (1'h1)))
        begin
          reg659 <= wire653;
          for (forvar660 = (1'h0); (forvar660 < (1'h1)); forvar660 = (forvar660 + (1'h1)))
            begin
              reg661 = ((-wire563[(5'h15):(4'h8)]) ? reg570 : "Eex");
              for (forvar662 = (1'h0); (forvar662 < (1'h0)); forvar662 = (forvar662 + (1'h1)))
                begin
                  reg663 <= {"lnCQTXe2h7NWFuTMYmcBb"};
                  reg664 <= "uc";
                  reg665 <= $unsigned({{((reg604 && forvar594) & $signed(forvar575))},
                      $signed((~reg633))});
                end
            end
          reg666 <= reg661[(1'h1):(1'h1)];
          reg667 <= ("qfuQ" | "Jgia8ELVxvIbFGb0");
          reg668 <= "75e8Y";
        end
    end
  always
    @(posedge clk) begin
      reg669 <= $signed((wire603[(2'h3):(1'h0)] || "RQu7ZeWK4KHx9xuq1wTQ0dhqD"));
      reg670 <= reg600[(5'h13):(5'h13)];
      reg671 <= reg639[(2'h3):(2'h3)];
      reg672 <= reg626;
      reg673 = $unsigned($signed($unsigned($unsigned(reg604))));
      reg674 = ((($signed((reg667 && (8'hbc))) ?
          ("tDi" ?
              ((8'hba) ?
                  forvar568 : reg629) : "4IwrD94FKBX4") : (~&(!reg634))) >> (reg625[(4'h9):(3'h7)] && $unsigned((+reg656)))) >>> ($signed(reg579[(4'hb):(3'h7)]) < $signed($signed({reg633}))));
    end
  assign wire675 = $signed("io66Lr3cWr");
  always
    @(posedge clk) begin
      reg676 <= $signed(reg586);
    end
  assign wire677 = reg606[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      reg678 <= $signed($signed((~^reg578)));
      reg679 <= (($signed((~forvar592[(2'h3):(1'h0)])) ^~ reg576[(4'h9):(3'h7)]) <<< (-(^~reg580[(1'h0):(1'h0)])));
      reg680 <= $unsigned({$unsigned((wire564[(2'h2):(1'h1)] ?
              $signed((7'h4e)) : (7'h42))),
          reg590[(2'h2):(1'h1)]});
      if ($signed((~$unsigned(reg638[(1'h1):(1'h1)]))))
        begin
          if ("hs")
            begin
              for (forvar681 = (1'h0); (forvar681 < (3'h5)); forvar681 = (forvar681 + (1'h1)))
                begin
                  reg682 <= (|(8'had));
                end
              reg683 <= $signed($unsigned((forvar568 == $signed($signed(reg678)))));
            end
          else
            begin
              reg681 <= ({reg574,
                  (forvar592[(4'hc):(3'h7)] ?
                      ((~forvar575) * reg613) : (^reg601[(2'h2):(2'h2)]))} <= $unsigned($signed(wire562[(3'h4):(3'h4)])));
              reg682 = $signed($signed($unsigned("WKUyuuwOn")));
            end
          reg684 <= {$unsigned((($signed(forvar568) ?
                  (reg640 && reg609) : reg680) ^~ reg624)),
              $unsigned("roeXFozglL5NABGdX9A")};
          reg685 <= wire561;
          reg686 <= $signed($unsigned(((+(reg645 ~^ wire565)) ?
              $unsigned((8'hbd)) : (~(~|reg641)))));
        end
      else
        begin
          reg681 <= "ycsYpWNhYvZdlNSNsfFPSqEy5";
          reg682 = reg584[(3'h4):(1'h1)];
          for (forvar683 = (1'h0); (forvar683 < (3'h5)); forvar683 = (forvar683 + (1'h1)))
            begin
              reg684 <= $unsigned($signed((~|$signed(reg664))));
            end
          reg685 <= (forvar572[(2'h3):(1'h0)] ?
              ((~&"") >> ($signed($signed(reg570)) ?
                  (8'h9c) : "2d5rrSb")) : (^~"7HMwNN"));
          reg686 <= "B2Gn";
        end
      reg687 <= "Ao0Uy8GaIgVGhiO2DL";
      reg688 = $signed(reg596);
    end
  always
    @(posedge clk) begin
      reg689 <= ((!(-reg688)) ?
          "fzGaZ3Dnt9QlMpWPV" : ((forvar575 >= ((forvar621 ?
                      (8'haf) : (8'ha1)) ?
                  "0RUSGde9" : $unsigned(reg648))) ?
              ((|reg676[(2'h2):(2'h2)]) >>> $signed(forvar592)) : (7'h49)));
      for (forvar690 = (1'h0); (forvar690 < (1'h1)); forvar690 = (forvar690 + (1'h1)))
        begin
          for (forvar691 = (1'h0); (forvar691 < (2'h3)); forvar691 = (forvar691 + (1'h1)))
            begin
              reg692 = reg581;
            end
          reg693 <= ((-$unsigned((^(~|reg645)))) ?
              {$signed((reg623 == (reg681 ? reg634 : (8'h9d)))),
                  {"oBS"}} : (&((forvar621[(2'h2):(2'h2)] ?
                  (wire565 < wire675) : reg571) + {$unsigned(reg610),
                  $signed((8'hb9))})));
        end
      reg694 <= ($signed($unsigned(forvar654[(2'h2):(2'h2)])) <<< $signed(forvar658[(5'h10):(4'h8)]));
    end
  assign wire695 = reg573;
  always
    @(posedge clk) begin
      reg696 <= {(8'ha4), (^~reg581[(3'h7):(1'h1)])};
      reg697 <= (~&{forvar662, $unsigned($unsigned(reg639))});
      reg698 <= reg576;
      reg699 <= $unsigned({(~&("" <= (^~(8'hb0)))), reg616});
      reg700 <= (^~$unsigned((reg684[(3'h7):(3'h5)] ?
          {reg644[(3'h5):(3'h4)], (8'haa)} : "Z0")));
    end
  always
    @(posedge clk) begin
      reg701 = {reg605};
      reg702 <= (reg610[(1'h0):(1'h0)] < ($unsigned($unsigned($signed((8'hb3)))) ?
          (7'h4b) : reg606[(1'h0):(1'h0)]));
      reg703 <= (~&(reg671[(4'he):(1'h0)] == (($signed(reg626) < ((7'h49) ?
          forvar643 : reg602)) + ($signed(reg589) && "csHVrbZTaDcIWuBT7bhY0i"))));
      reg704 <= (("K9mlcFAPD2n" ^ reg676) + reg692[(4'he):(4'hd)]);
    end
  assign wire705 = ((~^$signed(($signed(forvar690) & (reg570 ?
                       reg647 : forvar608)))) ^~ (^~$unsigned(($signed(forvar572) ?
                       (!reg688) : $unsigned((7'h44))))));
  assign wire706 = forvar575;
  always
    @(posedge clk) begin
      for (forvar707 = (1'h0); (forvar707 < (1'h1)); forvar707 = (forvar707 + (1'h1)))
        begin
          reg708 <= "LXgYis930GIt2DqN3LR";
          reg709 <= reg667[(4'h9):(1'h0)];
          reg710 <= ((reg669 * ($unsigned((reg692 <<< reg671)) & (~(~|reg632)))) | reg578[(3'h5):(1'h1)]);
          for (forvar711 = (1'h0); (forvar711 < (3'h5)); forvar711 = (forvar711 + (1'h1)))
            begin
              reg712 <= forvar691[(3'h4):(2'h2)];
              for (forvar713 = (1'h0); (forvar713 < (3'h4)); forvar713 = (forvar713 + (1'h1)))
                begin
                  reg714 = "IU1LIG3nHUi40V1z";
                  reg715 = reg571;
                end
              reg716 = (+$unsigned((reg613 ?
                  $signed($signed(reg630)) : $unsigned($signed(reg628)))));
              reg717 <= reg611;
              reg718 <= reg570[(3'h7):(3'h5)];
            end
          reg719 <= $unsigned((8'hb2));
          reg720 <= reg634[(2'h3):(2'h2)];
        end
    end
  always
    @(posedge clk) begin
      reg721 <= reg700;
      reg722 = reg644[(2'h3):(2'h3)];
    end
  always
    @(posedge clk) begin
      for (forvar723 = (1'h0); (forvar723 < (3'h5)); forvar723 = (forvar723 + (1'h1)))
        begin
          reg724 = (!"OnU41");
        end
      reg725 <= ((reg720[(4'hb):(2'h3)] >> wire695) ?
          (&$signed($unsigned(reg693))) : reg612[(1'h0):(1'h0)]);
      for (forvar726 = (1'h0); (forvar726 < (3'h4)); forvar726 = (forvar726 + (1'h1)))
        begin
          reg727 = reg601;
          reg728 <= reg715[(4'h9):(4'h9)];
          reg729 <= ((("p5h" ?
                  (reg670[(1'h1):(1'h1)] ?
                      "mUH" : (reg697 ? reg693 : reg626)) : (7'h44)) ?
              "" : $signed($unsigned((^reg582)))) + "XbLdBt5KTUDXUd");
          reg730 <= ($signed("xu41YxC3nbqQqxUko5") >= wire652[(2'h2):(2'h2)]);
          for (forvar731 = (1'h0); (forvar731 < (1'h0)); forvar731 = (forvar731 + (1'h1)))
            begin
              for (forvar732 = (1'h0); (forvar732 < (3'h4)); forvar732 = (forvar732 + (1'h1)))
                begin
                  reg733 <= (reg703[(4'hb):(1'h1)] && (("uO3GlOVXs" - ((&reg573) && $signed(forvar713))) ?
                      (((&reg622) ?
                          forvar723 : (~&reg620)) < reg630) : reg579[(2'h2):(1'h0)]));
                  reg734 <= $unsigned(((((wire564 > reg637) ~^ $unsigned(reg678)) == "NrzXWidIDobk") ?
                      (reg598[(2'h2):(2'h2)] ?
                          "E6KyxgKYIiAKfKAh" : "d7BIFJXBngCu") : ((wire705[(3'h6):(1'h0)] <<< "levgomARGwNNh") ^~ "xhD")));
                  reg735 <= "mDuYCmEfQS1omvsVEQpSq";
                  reg736 = {reg634};
                end
              reg737 <= reg671;
              reg738 <= forvar690;
            end
          for (forvar739 = (1'h0); (forvar739 < (3'h4)); forvar739 = (forvar739 + (1'h1)))
            begin
              reg740 <= $signed($unsigned($signed({reg702})));
              reg741 = ({(~|"Sy7kdTm4NCwzR5pbpw8q")} ?
                  reg570[(2'h2):(2'h2)] : "Ih7bIPBh4Uu3gx8L4yzHdv");
              reg742 <= reg655;
              for (forvar743 = (1'h0); (forvar743 < (2'h2)); forvar743 = (forvar743 + (1'h1)))
                begin
                  reg744 = reg622;
                end
              reg745 <= reg595;
              reg746 <= (~|$signed(reg638[(1'h1):(1'h0)]));
            end
        end
      reg747 = "DBwOlJVDadPhW";
    end
  always
    @(posedge clk) begin
      reg748 = reg629[(1'h0):(1'h0)];
      reg749 <= reg742[(3'h5):(1'h0)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module459
#( parameter param557 = ({(~|(((7'h42) & (8'hba)) > (~|(8'hb4))))} ? (((((8'hae) ? (8'haf) : (7'h4c)) && {(8'ha0)}) >>> {(~|(8'ha3))}) == (|({(7'h47)} ? {(7'h4d), (8'hb5)} : ((7'h4d) ? (8'h9c) : (8'hba))))) : {{(-((8'ha2) + (8'hb6))), (((8'hbf) ? (8'haa) : (8'ha7)) ? (~(7'h4a)) : {(8'hbe), (8'hae)})}}) )
(y, clk, wire464, wire463, wire462, wire461, wire460);
  output wire [(32'h504):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire464;
  input wire [(3'h4):(1'h0)] wire463;
  input wire signed [(5'h15):(1'h0)] wire462;
  input wire [(5'h16):(1'h0)] wire461;
  input wire signed [(5'h11):(1'h0)] wire460;
  wire signed [(4'he):(1'h0)] wire556;
  reg signed [(4'h8):(1'h0)] reg555 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg554 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg553 = (1'h0);
  reg [(5'h1a):(1'h0)] reg552 = (1'h0);
  reg [(3'h7):(1'h0)] forvar551 = (1'h0);
  reg [(3'h6):(1'h0)] reg550 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg549 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg548 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg547 = (1'h0);
  reg [(3'h7):(1'h0)] forvar546 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar545 = (1'h0);
  reg [(3'h7):(1'h0)] reg544 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg543 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg542 = (1'h0);
  reg [(5'h1a):(1'h0)] reg541 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg540 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar539 = (1'h0);
  reg [(2'h3):(1'h0)] reg538 = (1'h0);
  reg [(4'hc):(1'h0)] reg537 = (1'h0);
  reg [(4'hc):(1'h0)] reg536 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg535 = (1'h0);
  reg [(2'h3):(1'h0)] reg534 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg533 = (1'h0);
  reg [(2'h2):(1'h0)] reg532 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg531 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg530 = (1'h0);
  reg [(5'h17):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg528 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire527;
  reg [(5'h13):(1'h0)] reg526 = (1'h0);
  wire [(3'h5):(1'h0)] wire525;
  wire [(5'h1a):(1'h0)] wire524;
  reg signed [(4'hb):(1'h0)] reg523 = (1'h0);
  reg [(2'h2):(1'h0)] reg522 = (1'h0);
  reg [(4'hc):(1'h0)] reg521 = (1'h0);
  reg [(5'h19):(1'h0)] reg520 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg519 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg518 = (1'h0);
  reg [(5'h1a):(1'h0)] reg517 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg516 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg515 = (1'h0);
  reg [(4'hd):(1'h0)] reg514 = (1'h0);
  reg [(4'hf):(1'h0)] reg513 = (1'h0);
  reg [(4'he):(1'h0)] reg512 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg511 = (1'h0);
  reg [(5'h19):(1'h0)] reg510 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar508 = (1'h0);
  reg [(4'he):(1'h0)] reg507 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar506 = (1'h0);
  reg [(5'h10):(1'h0)] forvar505 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg504 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg503 = (1'h0);
  reg [(5'h13):(1'h0)] reg502 = (1'h0);
  reg [(4'he):(1'h0)] forvar501 = (1'h0);
  reg [(5'h17):(1'h0)] reg500 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg498 = (1'h0);
  reg [(5'h11):(1'h0)] reg497 = (1'h0);
  reg [(5'h1a):(1'h0)] reg496 = (1'h0);
  reg [(4'hc):(1'h0)] forvar495 = (1'h0);
  reg [(5'h17):(1'h0)] reg494 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar493 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg492 = (1'h0);
  reg [(4'hd):(1'h0)] reg491 = (1'h0);
  reg [(4'hb):(1'h0)] reg490 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg489 = (1'h0);
  reg [(2'h3):(1'h0)] reg488 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg487 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar486 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar485 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar484 = (1'h0);
  reg [(5'h12):(1'h0)] reg483 = (1'h0);
  reg [(2'h2):(1'h0)] reg482 = (1'h0);
  reg [(5'h14):(1'h0)] forvar481 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg480 = (1'h0);
  reg [(5'h17):(1'h0)] reg479 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg478 = (1'h0);
  reg [(4'he):(1'h0)] reg477 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar476 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg475 = (1'h0);
  reg [(5'h19):(1'h0)] reg474 = (1'h0);
  reg [(5'h18):(1'h0)] reg473 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg472 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg471 = (1'h0);
  reg [(3'h4):(1'h0)] forvar470 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg469 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg468 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar467 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg466 = (1'h0);
  wire [(5'h10):(1'h0)] wire465;
  assign y = {wire556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 forvar551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 forvar546,
                 forvar545,
                 reg544,
                 reg543,
                 reg542,
                 reg541,
                 reg540,
                 forvar539,
                 reg538,
                 reg537,
                 reg536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 wire527,
                 reg526,
                 wire525,
                 wire524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 reg517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 forvar508,
                 reg507,
                 forvar506,
                 forvar505,
                 reg504,
                 reg503,
                 reg502,
                 forvar501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 forvar495,
                 reg494,
                 forvar493,
                 reg492,
                 reg491,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 forvar486,
                 forvar485,
                 forvar484,
                 reg483,
                 reg482,
                 forvar481,
                 reg480,
                 reg479,
                 reg478,
                 reg477,
                 forvar476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 forvar470,
                 reg469,
                 reg468,
                 forvar467,
                 reg466,
                 wire465,
                 (1'h0)};
  assign wire465 = $signed(wire460);
  always
    @(posedge clk) begin
      reg466 <= "Bpb";
    end
  always
    @(posedge clk) begin
      for (forvar467 = (1'h0); (forvar467 < (2'h3)); forvar467 = (forvar467 + (1'h1)))
        begin
          reg468 <= $signed(wire465);
          reg469 <= "Oh5LYGzcmEK";
          for (forvar470 = (1'h0); (forvar470 < (3'h4)); forvar470 = (forvar470 + (1'h1)))
            begin
              reg471 <= $signed(($unsigned($signed("oCfdo")) - wire462[(4'hd):(1'h1)]));
              reg472 <= "UmIBNlsazWJ";
              reg473 <= (-$unsigned((^wire461[(4'hc):(4'hc)])));
              reg474 = wire464;
              reg475 <= $signed((&(~&$signed($signed(reg468)))));
              for (forvar476 = (1'h0); (forvar476 < (1'h0)); forvar476 = (forvar476 + (1'h1)))
                begin
                  reg477 <= (wire460 ?
                      (8'ha4) : ((|(wire464 ?
                          $signed((8'hbc)) : "v")) <<< wire460));
                  reg478 <= reg474[(5'h12):(4'h8)];
                  reg479 <= (|((7'h4a) << wire464[(4'h8):(2'h3)]));
                  reg480 <= ({wire462,
                      (reg468 && ((wire463 & reg474) <<< (+(8'hb8))))} ^ (8'hb0));
                end
            end
          for (forvar481 = (1'h0); (forvar481 < (3'h4)); forvar481 = (forvar481 + (1'h1)))
            begin
              reg482 <= reg469;
              reg483 <= (!(~|($signed((!(8'hb0))) || (~^$unsigned(reg478)))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar484 = (1'h0); (forvar484 < (2'h2)); forvar484 = (forvar484 + (1'h1)))
        begin
          for (forvar485 = (1'h0); (forvar485 < (2'h2)); forvar485 = (forvar485 + (1'h1)))
            begin
              for (forvar486 = (1'h0); (forvar486 < (1'h0)); forvar486 = (forvar486 + (1'h1)))
                begin
                  reg487 <= $signed((-("DPp88HZG43wl" ?
                      (reg483[(1'h0):(1'h0)] ?
                          {reg468, wire463} : (+reg475)) : reg466)));
                  reg488 <= (({((reg487 ^~ reg477) ?
                                  "sNFLRTOr0fxOw6JyeeCQC" : forvar476[(4'h8):(3'h4)]),
                              $unsigned($unsigned(wire463))} ?
                          (~&"ZdKViLRzlfQEkIxDL") : "") ?
                      "CtlvLYD6ol92d" : (|"VlsihvyVIVZ"));
                  reg489 = "sRe1pw5IyAYF1iTC";
                  reg490 <= reg466;
                  reg491 <= reg483[(2'h3):(1'h1)];
                end
              reg492 = wire465;
              for (forvar493 = (1'h0); (forvar493 < (1'h1)); forvar493 = (forvar493 + (1'h1)))
                begin
                  reg494 = (wire463 ? reg483[(3'h7):(3'h5)] : "rM");
                end
              for (forvar495 = (1'h0); (forvar495 < (1'h1)); forvar495 = (forvar495 + (1'h1)))
                begin
                  reg496 <= $unsigned(($unsigned(reg490) ^~ "ExeIeqr84qLVg"));
                  reg497 <= reg479[(3'h4):(2'h3)];
                  reg498 <= (~|reg468);
                  reg499 = (~^$unsigned(((reg494[(1'h1):(1'h0)] ?
                      (reg474 ?
                          (8'ha7) : reg487) : {forvar486}) * $signed(reg496[(2'h2):(1'h0)]))));
                end
              reg500 <= (^~(+reg496[(4'hd):(4'hd)]));
            end
          for (forvar501 = (1'h0); (forvar501 < (3'h4)); forvar501 = (forvar501 + (1'h1)))
            begin
              reg502 <= "3FpoTG4FrGN";
              reg503 = reg478;
              reg504 <= ((^(^~$signed($unsigned(forvar467)))) && (!((&{reg491}) ?
                  (~^"CUqbBnPAzf3evxGh579X") : (+wire460[(3'h4):(1'h1)]))));
            end
        end
      for (forvar505 = (1'h0); (forvar505 < (1'h1)); forvar505 = (forvar505 + (1'h1)))
        begin
          for (forvar506 = (1'h0); (forvar506 < (1'h1)); forvar506 = (forvar506 + (1'h1)))
            begin
              reg507 <= "";
              for (forvar508 = (1'h0); (forvar508 < (2'h3)); forvar508 = (forvar508 + (1'h1)))
                begin
                  reg509 <= (&reg483[(4'hc):(2'h2)]);
                  reg510 <= "VcfkN4ZMubQEwB8eY1";
                  reg511 <= "fh5ON9J";
                  reg512 <= reg498[(1'h0):(1'h0)];
                  reg513 <= $unsigned((reg497 <= reg502));
                  reg514 <= "cyqMC";
                end
              reg515 <= reg471;
              reg516 <= reg479[(5'h10):(1'h1)];
            end
          reg517 <= ("diDAk" && $unsigned($signed({$unsigned(reg489),
              forvar481})));
        end
    end
  always
    @(posedge clk) begin
      reg518 <= "cIGRYmVZF7";
    end
  always
    @(posedge clk) begin
      reg519 <= "7IE4LgRkJstn37ch";
      reg520 = $signed(reg469);
      reg521 <= (8'hbc);
      reg522 <= (reg512 & forvar485);
      reg523 <= ((forvar501[(4'h9):(2'h2)] ?
              (reg509[(1'h0):(1'h0)] == $signed(wire463)) : reg468[(3'h4):(2'h3)]) ?
          (reg518[(2'h3):(1'h0)] ?
              reg494 : forvar481[(5'h13):(3'h7)]) : {((~|(reg496 ?
                  reg469 : (8'hbf))) > "7Qh4TbvTk"),
              (({reg483, reg483} ? "b" : reg510) ?
                  forvar476 : (&wire461[(5'h16):(4'h8)]))});
    end
  assign wire524 = ($unsigned($signed($signed(((7'h4e) ? reg512 : reg510)))) ?
                       (&reg521) : "Erren0tMTNg7NXqpxt");
  assign wire525 = forvar506[(3'h5):(2'h2)];
  always
    @(posedge clk) begin
      reg526 <= $unsigned((&(-reg490)));
    end
  assign wire527 = reg496;
  always
    @(posedge clk) begin
      reg528 <= reg502[(2'h3):(2'h3)];
      reg529 <= (+$signed(({reg522} ?
          "Ua" : ($signed((8'hb9)) ? (+reg528) : forvar470[(1'h1):(1'h1)]))));
      reg530 <= reg511;
      reg531 <= ((^"fVk") ?
          "n0b2QBaoS7dIllMzda" : (-$signed(($signed(wire462) ?
              $unsigned(reg519) : "fZO6B4rcMqsGzNB5MHe9y7Usc"))));
      reg532 <= (+(7'h49));
    end
  always
    @(posedge clk) begin
      reg533 <= forvar476[(2'h2):(2'h2)];
      reg534 <= forvar505;
    end
  always
    @(posedge clk) begin
      reg535 <= "uMx7";
      reg536 <= $signed(reg490[(1'h1):(1'h1)]);
      reg537 <= (("JM4vTNm" + $signed(reg528)) ^~ $signed((reg473 * wire460[(4'hf):(3'h7)])));
      reg538 <= (((reg536[(4'hc):(1'h1)] ? "AohTJmWscxsSehA0VGo" : reg504) ?
              wire465[(4'he):(4'hd)] : wire525[(2'h3):(1'h0)]) ?
          $signed((({reg500, (8'hb2)} > (~^forvar470)) ?
              (reg521 ? (reg468 || reg500) : (!reg474)) : forvar506)) : reg526);
    end
  always
    @(posedge clk) begin
      for (forvar539 = (1'h0); (forvar539 < (3'h5)); forvar539 = (forvar539 + (1'h1)))
        begin
          reg540 <= $signed(reg526[(3'h5):(2'h2)]);
          reg541 <= "P";
          reg542 = "iVeqKcHUdrC0HdeoKb";
        end
      reg543 <= "Jyy5WSPNv60";
      reg544 <= $unsigned((reg538[(2'h2):(1'h0)] == (-forvar539)));
    end
  always
    @(posedge clk) begin
      for (forvar545 = (1'h0); (forvar545 < (1'h0)); forvar545 = (forvar545 + (1'h1)))
        begin
          for (forvar546 = (1'h0); (forvar546 < (3'h5)); forvar546 = (forvar546 + (1'h1)))
            begin
              reg547 = reg480;
              reg548 = reg515[(4'hb):(2'h3)];
              reg549 <= "SIOL5x9vr";
            end
          reg550 <= "2tr189RtWpTx2eh5Dusr";
        end
      for (forvar551 = (1'h0); (forvar551 < (1'h0)); forvar551 = (forvar551 + (1'h1)))
        begin
          reg552 <= "gN1x";
          reg553 <= ((+$unsigned({""})) ?
              "b" : ($unsigned("BScbrbNPGIP4vvGLvJgK") == ("0FSCSZ1n2yvpilkEalcsUu" ?
                  ((reg522 >= reg487) * $unsigned(reg509)) : $unsigned(reg538[(2'h3):(2'h2)]))));
        end
      reg554 <= (8'ha6);
      reg555 <= ($unsigned($signed(reg515)) ?
          {(-"T6QAmbWKAAn"),
              "22xm1Mbc6wumGU1kZF"} : ({"RzT3AOXZt1KqQn"} | ($unsigned(((8'ha4) & reg516)) ?
              reg487[(5'h10):(1'h0)] : "nMyYcnJ2rJs2yWeiy")));
    end
  assign wire556 = reg554[(4'hc):(3'h5)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module219
#( parameter param444 = ((7'h4b) ? ({({(8'hbd), (8'haa)} - (~^(8'hbb)))} * (^{((7'h43) ? (7'h40) : (8'h9c))})) : {(((&(8'haf)) >> (&(8'ha9))) >= ((~|(8'ha7)) ? {(8'hb9)} : (~&(8'ha7))))})
, parameter param445 = (param444 ~^ param444) )
(y, clk, wire223, wire222, wire221, wire220);
  output wire [(32'hc96):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire223;
  input wire [(5'h12):(1'h0)] wire222;
  input wire signed [(4'h8):(1'h0)] wire221;
  input wire [(4'ha):(1'h0)] wire220;
  wire [(5'h17):(1'h0)] wire443;
  wire signed [(5'h18):(1'h0)] wire442;
  wire [(5'h19):(1'h0)] wire441;
  wire signed [(5'h13):(1'h0)] wire440;
  reg signed [(5'h18):(1'h0)] reg439 = (1'h0);
  reg [(3'h5):(1'h0)] reg438 = (1'h0);
  reg [(3'h6):(1'h0)] reg437 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg436 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg435 = (1'h0);
  reg [(4'h8):(1'h0)] reg434 = (1'h0);
  reg [(3'h7):(1'h0)] reg433 = (1'h0);
  reg [(5'h17):(1'h0)] reg432 = (1'h0);
  reg [(5'h11):(1'h0)] forvar431 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg430 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg415 = (1'h0);
  reg [(3'h6):(1'h0)] reg429 = (1'h0);
  reg [(5'h13):(1'h0)] reg428 = (1'h0);
  reg [(5'h17):(1'h0)] reg427 = (1'h0);
  reg [(4'h9):(1'h0)] reg426 = (1'h0);
  reg [(3'h7):(1'h0)] reg425 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg424 = (1'h0);
  reg [(4'hc):(1'h0)] reg423 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg422 = (1'h0);
  reg [(3'h7):(1'h0)] forvar421 = (1'h0);
  reg [(3'h4):(1'h0)] reg420 = (1'h0);
  reg [(5'h1a):(1'h0)] reg419 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg418 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg417 = (1'h0);
  reg [(5'h18):(1'h0)] reg416 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar415 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg414 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg413 = (1'h0);
  reg [(3'h5):(1'h0)] forvar412 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire411;
  reg [(5'h10):(1'h0)] reg410 = (1'h0);
  reg [(3'h6):(1'h0)] reg409 = (1'h0);
  reg [(4'hf):(1'h0)] reg408 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg407 = (1'h0);
  reg [(5'h18):(1'h0)] reg406 = (1'h0);
  reg [(4'h9):(1'h0)] reg405 = (1'h0);
  reg [(2'h3):(1'h0)] forvar404 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg403 = (1'h0);
  reg [(2'h2):(1'h0)] reg402 = (1'h0);
  reg [(4'hc):(1'h0)] reg401 = (1'h0);
  reg [(5'h13):(1'h0)] reg400 = (1'h0);
  reg [(2'h2):(1'h0)] reg399 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg398 = (1'h0);
  reg [(2'h3):(1'h0)] forvar397 = (1'h0);
  reg [(5'h18):(1'h0)] forvar396 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg394 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg393 = (1'h0);
  reg [(5'h12):(1'h0)] reg392 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg391 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg390 = (1'h0);
  reg [(3'h7):(1'h0)] reg389 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg388 = (1'h0);
  reg [(5'h19):(1'h0)] reg387 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg386 = (1'h0);
  reg [(4'h8):(1'h0)] reg385 = (1'h0);
  reg [(4'h9):(1'h0)] forvar384 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg383 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg382 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg381 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar380 = (1'h0);
  reg [(5'h1a):(1'h0)] reg379 = (1'h0);
  reg [(5'h15):(1'h0)] reg378 = (1'h0);
  reg [(5'h19):(1'h0)] reg377 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar376 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg375 = (1'h0);
  reg [(5'h16):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg373 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar372 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar371 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg370 = (1'h0);
  reg [(5'h16):(1'h0)] reg369 = (1'h0);
  reg [(4'h9):(1'h0)] reg368 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg367 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg366 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg365 = (1'h0);
  reg [(3'h6):(1'h0)] reg364 = (1'h0);
  reg [(4'h9):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg362 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar361 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar360 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar359 = (1'h0);
  reg [(5'h14):(1'h0)] reg358 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg357 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg356 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar355 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg354 = (1'h0);
  reg [(4'h8):(1'h0)] reg353 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar352 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg351 = (1'h0);
  reg [(5'h13):(1'h0)] reg350 = (1'h0);
  reg [(5'h15):(1'h0)] reg349 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg348 = (1'h0);
  reg [(2'h2):(1'h0)] reg347 = (1'h0);
  reg [(5'h12):(1'h0)] reg346 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar345 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar344 = (1'h0);
  reg [(5'h1a):(1'h0)] reg343 = (1'h0);
  reg [(5'h10):(1'h0)] reg342 = (1'h0);
  reg [(5'h12):(1'h0)] reg341 = (1'h0);
  reg [(4'hb):(1'h0)] reg340 = (1'h0);
  reg [(5'h19):(1'h0)] reg339 = (1'h0);
  reg [(2'h2):(1'h0)] reg338 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg337 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg336 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg335 = (1'h0);
  reg [(3'h6):(1'h0)] reg334 = (1'h0);
  reg [(5'h11):(1'h0)] reg333 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar332 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg331 = (1'h0);
  reg [(3'h4):(1'h0)] forvar330 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar329 = (1'h0);
  reg [(3'h6):(1'h0)] reg328 = (1'h0);
  reg [(5'h1a):(1'h0)] reg327 = (1'h0);
  reg [(5'h16):(1'h0)] reg326 = (1'h0);
  reg signed [(4'he):(1'h0)] reg325 = (1'h0);
  reg [(4'hd):(1'h0)] reg324 = (1'h0);
  reg [(5'h13):(1'h0)] reg323 = (1'h0);
  reg [(5'h14):(1'h0)] forvar322 = (1'h0);
  reg [(4'hb):(1'h0)] reg321 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar320 = (1'h0);
  reg [(3'h4):(1'h0)] reg319 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar316 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg315 = (1'h0);
  reg [(4'h9):(1'h0)] reg314 = (1'h0);
  reg [(2'h3):(1'h0)] reg313 = (1'h0);
  reg [(4'h8):(1'h0)] forvar312 = (1'h0);
  reg [(4'hc):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar310 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg308 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg307 = (1'h0);
  reg [(4'hb):(1'h0)] reg306 = (1'h0);
  reg [(2'h3):(1'h0)] reg305 = (1'h0);
  reg [(2'h3):(1'h0)] reg304 = (1'h0);
  reg [(2'h2):(1'h0)] forvar299 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar298 = (1'h0);
  reg signed [(4'he):(1'h0)] reg297 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg303 = (1'h0);
  reg [(5'h14):(1'h0)] reg302 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg301 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg300 = (1'h0);
  reg [(5'h10):(1'h0)] reg299 = (1'h0);
  reg [(2'h2):(1'h0)] reg298 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar297 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg296 = (1'h0);
  reg [(4'hf):(1'h0)] reg295 = (1'h0);
  reg [(5'h19):(1'h0)] reg294 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg293 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar292 = (1'h0);
  reg [(4'he):(1'h0)] forvar291 = (1'h0);
  reg [(5'h12):(1'h0)] reg290 = (1'h0);
  reg [(5'h13):(1'h0)] reg289 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire288;
  reg signed [(4'hd):(1'h0)] reg287 = (1'h0);
  reg [(3'h4):(1'h0)] reg286 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg285 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg284 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg283 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar282 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg281 = (1'h0);
  reg [(5'h1a):(1'h0)] reg280 = (1'h0);
  reg [(5'h10):(1'h0)] reg279 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg278 = (1'h0);
  reg [(5'h11):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg276 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg275 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg274 = (1'h0);
  reg [(4'hb):(1'h0)] forvar273 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg272 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg271 = (1'h0);
  reg [(5'h12):(1'h0)] forvar270 = (1'h0);
  reg [(4'h8):(1'h0)] reg269 = (1'h0);
  reg [(5'h1a):(1'h0)] reg268 = (1'h0);
  reg [(5'h17):(1'h0)] reg267 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar266 = (1'h0);
  reg [(4'he):(1'h0)] reg265 = (1'h0);
  reg [(5'h17):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg263 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg262 = (1'h0);
  reg [(3'h4):(1'h0)] reg261 = (1'h0);
  reg [(5'h1a):(1'h0)] reg260 = (1'h0);
  reg [(4'h8):(1'h0)] reg259 = (1'h0);
  reg [(4'hc):(1'h0)] forvar258 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar257 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg256 = (1'h0);
  reg [(5'h18):(1'h0)] reg255 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg254 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg253 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg252 = (1'h0);
  reg [(5'h19):(1'h0)] reg251 = (1'h0);
  reg [(5'h15):(1'h0)] reg250 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar249 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg248 = (1'h0);
  reg [(4'h9):(1'h0)] reg247 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg246 = (1'h0);
  reg [(5'h10):(1'h0)] reg245 = (1'h0);
  reg [(5'h15):(1'h0)] reg244 = (1'h0);
  reg [(5'h15):(1'h0)] reg243 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg241 = (1'h0);
  reg [(5'h17):(1'h0)] forvar239 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar238 = (1'h0);
  reg [(5'h13):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg240 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg239 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg238 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg237 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg236 = (1'h0);
  reg [(5'h1a):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar234 = (1'h0);
  wire [(3'h7):(1'h0)] wire233;
  wire signed [(4'hc):(1'h0)] wire232;
  reg [(3'h7):(1'h0)] reg231 = (1'h0);
  reg [(5'h19):(1'h0)] reg230 = (1'h0);
  reg [(4'hd):(1'h0)] reg229 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg228 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg227 = (1'h0);
  reg [(4'ha):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg225 = (1'h0);
  reg [(5'h15):(1'h0)] reg224 = (1'h0);
  assign y = {wire443,
                 wire442,
                 wire441,
                 wire440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 forvar431,
                 reg430,
                 reg415,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 forvar421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 forvar415,
                 reg414,
                 reg413,
                 forvar412,
                 wire411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 forvar404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 forvar397,
                 forvar396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 forvar384,
                 reg383,
                 reg382,
                 reg381,
                 forvar380,
                 reg379,
                 reg378,
                 reg377,
                 forvar376,
                 reg375,
                 reg374,
                 reg373,
                 forvar372,
                 forvar371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 reg362,
                 forvar361,
                 forvar360,
                 forvar359,
                 reg358,
                 reg357,
                 reg356,
                 forvar355,
                 reg354,
                 reg353,
                 forvar352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 forvar345,
                 forvar344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 forvar332,
                 reg331,
                 forvar330,
                 forvar329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 reg323,
                 forvar322,
                 reg321,
                 forvar320,
                 reg319,
                 reg318,
                 reg317,
                 forvar316,
                 reg315,
                 reg314,
                 reg313,
                 forvar312,
                 reg311,
                 forvar310,
                 reg309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 forvar299,
                 forvar298,
                 reg297,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 forvar297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 forvar292,
                 forvar291,
                 reg290,
                 reg289,
                 wire288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 forvar282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 forvar273,
                 reg272,
                 reg271,
                 forvar270,
                 reg269,
                 reg268,
                 reg267,
                 forvar266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 forvar258,
                 forvar257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 forvar249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 forvar239,
                 forvar238,
                 reg234,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 forvar234,
                 wire233,
                 wire232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg224 <= ("B" < $signed(wire220[(2'h3):(1'h0)]));
      reg225 <= wire222;
      reg226 <= (^wire221);
      reg227 = ((+wire221) ?
          (wire223[(1'h1):(1'h0)] <<< $signed({$signed((8'hac)),
              $unsigned((8'hbe))})) : (!{reg226[(1'h0):(1'h0)],
              "L2kEnMeX8tGPvvXQCPQHuM4"}));
      reg228 = "B2zkM95ZCO7WT6tezw";
      reg229 = wire221;
    end
  always
    @(posedge clk) begin
      reg230 <= ((((((8'hb0) ?
              reg226 : reg224) == $unsigned(wire221)) ^ "pGK47") ?
          reg224[(1'h1):(1'h0)] : (~^$signed($signed(reg225)))) <<< reg228);
      reg231 <= (8'haf);
    end
  assign wire232 = reg227;
  assign wire233 = ({{$signed("ielkFaOM1q"), (!reg228[(1'h1):(1'h0)])},
                           "EXrTfTCOzMkmLfyc"} ?
                       $unsigned(("d2RgfKWf3E3kB152Tel8yyH" ^ reg229[(1'h0):(1'h0)])) : "VczWnYyCvzQWbxUTgXGQfh");
  always
    @(posedge clk) begin
      if ({$unsigned(((^(reg231 ?
              wire233 : (8'ha8))) <<< $unsigned("SdrZBs1Ymz1HxUd")))})
        begin
          for (forvar234 = (1'h0); (forvar234 < (2'h2)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 <= forvar234[(1'h1):(1'h1)];
              reg236 <= $unsigned("dzPldclfKCtoHR");
            end
          reg237 = ((+(^$unsigned((reg230 ^ wire232)))) ?
              reg227 : wire223[(1'h1):(1'h1)]);
          reg238 <= {"Y43", $unsigned("edVM")};
          reg239 <= reg235[(2'h2):(1'h0)];
          reg240 = (~^wire221);
        end
      else
        begin
          reg234 <= (~|$unsigned($unsigned($signed((wire223 << wire220)))));
          reg235 = (reg240 ? reg227[(5'h11):(4'hd)] : wire223[(2'h3):(1'h0)]);
          reg236 <= "hhVLPg9uEr";
          reg237 <= {reg235[(3'h7):(2'h2)]};
          for (forvar238 = (1'h0); (forvar238 < (1'h1)); forvar238 = (forvar238 + (1'h1)))
            begin
              for (forvar239 = (1'h0); (forvar239 < (2'h3)); forvar239 = (forvar239 + (1'h1)))
                begin
                  reg240 <= ({(~&({forvar239} ?
                              $signed(reg226) : $signed((7'h48)))),
                          $signed(reg238)} ?
                      (wire233 > (("x8ok7U6NHp" ? (reg236 ^ reg239) : reg235) ?
                          (reg237[(2'h3):(1'h0)] != (forvar234 ?
                              wire220 : reg235)) : {"vvLsp7qpcGY"})) : (~((7'h40) ^ {{reg234,
                              reg238},
                          (reg235 < reg238)})));
                end
              reg241 <= $unsigned($unsigned(wire232));
              reg242 <= "EY2kUbz8f";
              reg243 <= ("QAC4eLzlmwSiAaxoP" > $signed($signed(("SzNErE" < (-reg229)))));
            end
          reg244 = (forvar234 * (|$signed(($signed(reg228) >> (reg234 >> reg229)))));
        end
      reg245 <= (reg225[(5'h14):(5'h11)] ? "ZU13apxrcyF1SCqy42Vr" : (+"X"));
      reg246 <= (8'ha7);
      reg247 = (~&((&({reg243, wire220} & "z64eIV")) & reg237));
      reg248 <= $signed($unsigned(("XG" ^ (^~wire221[(3'h5):(3'h4)]))));
    end
  always
    @(posedge clk) begin
      for (forvar249 = (1'h0); (forvar249 < (2'h3)); forvar249 = (forvar249 + (1'h1)))
        begin
          reg250 <= (($unsigned({(-reg245),
                  "MpBm689z"}) <= (^~{$unsigned(reg225)})) ?
              wire222 : wire232[(3'h5):(3'h4)]);
          reg251 <= {$unsigned((("2CwPhtOwDxtqHPQWaCNUcDrp" ?
                  "MqVqvWVxWc7FfqnX8" : wire221[(3'h5):(1'h1)]) >= ((reg243 ?
                  wire233 : wire232) != (reg241 ? reg237 : reg239)))),
              ((|"6fBIK") ? "hWRMJREh" : wire222[(3'h7):(3'h5)])};
        end
      reg252 <= reg246[(3'h5):(1'h0)];
      reg253 <= reg244[(4'ha):(3'h6)];
    end
  always
    @(posedge clk) begin
      reg254 <= $signed(("06xA1ubCacm1GP4bP" ?
          "E9h8x3uMJoPqVYFEcaLUXx" : reg239[(4'he):(3'h6)]));
      reg255 <= "tDc7C4x70RmZFC0vRFhlxG";
      reg256 <= $unsigned(reg255[(5'h10):(4'h8)]);
      for (forvar257 = (1'h0); (forvar257 < (2'h3)); forvar257 = (forvar257 + (1'h1)))
        begin
          for (forvar258 = (1'h0); (forvar258 < (3'h5)); forvar258 = (forvar258 + (1'h1)))
            begin
              reg259 <= wire233[(1'h1):(1'h1)];
              reg260 <= (~reg252[(1'h1):(1'h1)]);
              reg261 <= {$signed(($signed($unsigned(wire223)) >= "PeDDQM8snoGK1AZMDsi0")),
                  reg247[(3'h6):(3'h6)]};
              reg262 <= $signed(wire233);
              reg263 <= $signed(((forvar234 < (~^(reg256 - (8'ha1)))) ?
                  $unsigned((reg253[(5'h13):(1'h1)] & (wire221 ?
                      reg228 : reg227))) : (^~reg251)));
            end
          reg264 <= forvar234[(4'h9):(3'h6)];
          reg265 = {reg248};
          for (forvar266 = (1'h0); (forvar266 < (3'h4)); forvar266 = (forvar266 + (1'h1)))
            begin
              reg267 <= {reg264[(4'ha):(2'h3)]};
              reg268 <= ($unsigned((($signed(reg259) ?
                  $signed(reg228) : $signed(reg224)) == ($signed((8'hb3)) ?
                  $signed(reg235) : (-reg224)))) - $unsigned((((^forvar239) ?
                      "wr8AcAahS" : $signed(reg254)) ?
                  ((reg244 ?
                      reg230 : (8'h9e)) >= forvar249[(4'h9):(3'h4)]) : "Epn")));
            end
          reg269 <= wire222[(4'h9):(4'h8)];
        end
      for (forvar270 = (1'h0); (forvar270 < (1'h1)); forvar270 = (forvar270 + (1'h1)))
        begin
          reg271 <= reg237[(3'h6):(1'h0)];
          reg272 <= $unsigned($signed("C6X7CEhvpPQh1WlIhE3VrGsRK"));
          for (forvar273 = (1'h0); (forvar273 < (2'h2)); forvar273 = (forvar273 + (1'h1)))
            begin
              if ((^~$signed({(-(reg255 != (7'h4c)))})))
                begin
                  reg274 = "lY9vVAkNEwuAh8Y";
                  reg275 <= $unsigned($unsigned({"HZqA"}));
                  reg276 <= "";
                end
              else
                begin
                  reg274 <= reg236[(4'ha):(2'h3)];
                  reg275 <= (~($signed({$signed(reg238)}) ?
                      forvar258[(1'h0):(1'h0)] : (!$unsigned({reg261}))));
                end
              reg277 <= {(reg228[(2'h3):(1'h1)] ?
                      reg274 : ({$unsigned(forvar238),
                          (reg239 >= (7'h44))} << "v3tHM5u7yvfdu")),
                  $unsigned($unsigned((&$signed(reg228))))};
              if ($signed(("r" ?
                  (forvar239[(1'h0):(1'h0)] >> reg241[(4'ha):(2'h3)]) : (&reg256))))
                begin
                  reg278 <= (~&(~^{$unsigned(reg268),
                      ("bw2fGRRcgzBrk5WkDa6LlnVAT" ?
                          forvar273 : (^forvar249))}));
                  reg279 <= reg268[(5'h11):(3'h6)];
                end
              else
                begin
                  reg278 <= (reg244[(1'h1):(1'h1)] ?
                      (reg265[(4'hc):(4'ha)] ?
                          "HiYzyNOCrl" : ($signed({reg254,
                              reg238}) & reg252[(4'hc):(4'h8)])) : "tY4Pt1HFuPEUSEJxivyO2UsS");
                end
            end
          reg280 = "cgkVoVecGWlX";
          reg281 <= $unsigned($unsigned($unsigned(((reg227 < reg250) ?
              reg274 : (~reg271)))));
        end
      for (forvar282 = (1'h0); (forvar282 < (2'h3)); forvar282 = (forvar282 + (1'h1)))
        begin
          reg283 <= reg241[(4'h8):(3'h6)];
          reg284 <= (^(reg262 ?
              ($unsigned($unsigned(reg225)) >> reg255[(1'h1):(1'h0)]) : (-$unsigned((~&reg275)))));
        end
    end
  always
    @(posedge clk) begin
      reg285 <= {(&$signed($signed("YKNHhNnB"))), (^reg262)};
      reg286 = reg243;
      reg287 <= ((~^reg253[(4'ha):(4'h8)]) ?
          reg234[(4'hd):(4'h8)] : ("kT" || "IHwfS78AiHkJLoq"));
    end
  assign wire288 = $signed(forvar238);
  always
    @(posedge clk) begin
      reg289 <= reg231;
      reg290 = $unsigned(forvar258[(2'h3):(1'h0)]);
      for (forvar291 = (1'h0); (forvar291 < (3'h5)); forvar291 = (forvar291 + (1'h1)))
        begin
          for (forvar292 = (1'h0); (forvar292 < (3'h4)); forvar292 = (forvar292 + (1'h1)))
            begin
              reg293 <= (((wire288[(4'hf):(2'h3)] ?
                  ((reg261 ? reg274 : reg285) ?
                      (8'hb6) : $signed(forvar239)) : ($signed(reg231) ?
                      (reg275 ?
                          forvar266 : wire233) : (reg280 - (7'h47)))) > (("QAdK0" ?
                      "a4" : "AsSeB77zcAYADhuBiz") ?
                  $unsigned(reg239[(4'he):(3'h5)]) : ("t2kD3gwKuCTRy815I0r71JKJY" > "Lv8yfSyMmzUO"))) ^~ "Fmy0JWWndo");
            end
        end
      reg294 <= wire288[(3'h4):(1'h0)];
      if ((-$unsigned((wire223 << (8'ha0)))))
        begin
          reg295 = $signed($unsigned({$unsigned((8'hb0)),
              ("53xHKYS9qBLYZf8v5zvpeCV0" * $unsigned(reg230))}));
          reg296 <= (forvar266[(1'h0):(1'h0)] ?
              $unsigned($unsigned("qqKCiVqiIci")) : (8'ha7));
          for (forvar297 = (1'h0); (forvar297 < (2'h3)); forvar297 = (forvar297 + (1'h1)))
            begin
              if ($unsigned(((~|((~reg241) << (+reg242))) ?
                  {$unsigned("a"), $unsigned({reg245})} : reg245)))
                begin
                  reg298 <= "1ZaAsFWd714z5Rm2w3BJ";
                  reg299 <= $unsigned($signed("lA22d"));
                  reg300 <= {"DueIAurolwKH7aq7F", "4FDNs6aNLGJ27hlBKA4q1Y"};
                end
              else
                begin
                  reg298 <= (|reg279[(1'h0):(1'h0)]);
                end
              reg301 <= $signed(wire222[(2'h2):(2'h2)]);
              reg302 = {"XpF8u"};
            end
          reg303 <= {(($unsigned((reg267 ?
                  reg276 : forvar257)) <= $signed(reg302)) <<< reg275[(2'h2):(1'h0)])};
        end
      else
        begin
          reg295 <= ((~reg299[(4'hc):(1'h1)]) | ($unsigned(reg231[(1'h0):(1'h0)]) * ({"s6aQT",
                  (forvar258 >>> reg295)} ?
              "r1Ab" : "QUPo1ozGVWK8oSUmKow")));
          reg296 <= (^~{($unsigned($signed(reg252)) >= ("xVVOtHDUnqO" ?
                  $unsigned(reg286) : reg253[(1'h1):(1'h1)]))});
          reg297 <= $unsigned($signed(((reg241[(4'hf):(3'h6)] > reg295[(4'hb):(2'h2)]) ?
              reg235 : forvar249)));
          for (forvar298 = (1'h0); (forvar298 < (3'h4)); forvar298 = (forvar298 + (1'h1)))
            begin
              for (forvar299 = (1'h0); (forvar299 < (1'h0)); forvar299 = (forvar299 + (1'h1)))
                begin
                  reg300 <= (7'h40);
                  reg301 <= (reg240[(4'hb):(4'hb)] ?
                      (&reg286[(1'h1):(1'h0)]) : ($signed(reg293) ?
                          $unsigned(reg247) : (~reg225)));
                  reg302 <= $signed(({$unsigned($unsigned(reg279))} ?
                      ((-(7'h45)) ?
                          (8'ha8) : ("eEarMrl4dzrkSKkFVM" ?
                              reg234 : $unsigned(reg224))) : (^~$unsigned(reg239))));
                  reg303 <= reg284;
                end
              reg304 <= $unsigned(reg298);
              reg305 = ("qTCO8" << (8'haa));
              reg306 <= {(((reg287[(2'h2):(1'h1)] ?
                              (~^wire223) : (wire223 * reg261)) ?
                          $signed(reg297[(4'hc):(3'h6)]) : reg303[(2'h2):(1'h1)]) ?
                      $signed($unsigned((&reg301))) : reg253),
                  (+(-"n0S2I6ItVdD4"))};
              reg307 <= (8'ha8);
              reg308 = $unsigned((+$signed(reg279[(4'hf):(3'h6)])));
            end
          reg309 = ((~^((!reg299) ?
              "EVTH" : "gfLr2LPUd3YGWrtD")) + $signed((($unsigned(wire288) >= (~&reg275)) == reg242[(4'hc):(3'h7)])));
          for (forvar310 = (1'h0); (forvar310 < (3'h4)); forvar310 = (forvar310 + (1'h1)))
            begin
              reg311 <= $unsigned({{$signed((reg278 ~^ reg287))},
                  $unsigned((~((8'hbb) && reg267)))});
              for (forvar312 = (1'h0); (forvar312 < (1'h1)); forvar312 = (forvar312 + (1'h1)))
                begin
                  reg313 = "1ZmKYO";
                end
              reg314 <= reg234[(5'h13):(1'h1)];
            end
        end
      reg315 <= ({($signed(((7'h41) ? forvar292 : reg242)) ?
                  (|{reg275, reg287}) : $signed(reg237)),
              reg280[(5'h12):(4'hf)]} ?
          ({(~^(8'hbc)), $signed("VXsUaowqLdzANP4")} ?
              (&$signed((reg307 >> (7'h42)))) : ((-$unsigned(reg259)) == ($unsigned(reg300) ?
                  (^(8'hac)) : (forvar299 + (8'hb1))))) : reg267[(3'h7):(2'h3)]);
    end
  always
    @(posedge clk) begin
      for (forvar316 = (1'h0); (forvar316 < (2'h3)); forvar316 = (forvar316 + (1'h1)))
        begin
          reg317 <= forvar234[(4'hc):(3'h4)];
          reg318 <= $unsigned("f5iQKkDLEZks2mmQ7nn3");
          reg319 <= {(~|{reg309[(4'ha):(4'h9)]}),
              {{$unsigned("zv8tb2UCbrniJHE"), reg267}}};
          for (forvar320 = (1'h0); (forvar320 < (2'h3)); forvar320 = (forvar320 + (1'h1)))
            begin
              reg321 = reg298;
              for (forvar322 = (1'h0); (forvar322 < (2'h2)); forvar322 = (forvar322 + (1'h1)))
                begin
                  reg323 <= ($unsigned(reg307) && ("TMpgQN7d" + "0XF1Q83Cw1"));
                  reg324 <= (^~forvar292);
                  reg325 <= "4fw";
                end
            end
          reg326 = forvar291[(2'h2):(1'h1)];
          reg327 <= (~reg301[(2'h2):(1'h0)]);
        end
      reg328 <= (reg323 <<< (((^{reg289}) && $signed({(8'ha1), reg302})) ?
          $signed({forvar239[(5'h13):(3'h5)],
              forvar298[(4'hc):(4'hc)]}) : (-{reg269[(3'h7):(3'h7)],
              (reg285 >>> reg268)})));
      for (forvar329 = (1'h0); (forvar329 < (2'h3)); forvar329 = (forvar329 + (1'h1)))
        begin
          for (forvar330 = (1'h0); (forvar330 < (2'h3)); forvar330 = (forvar330 + (1'h1)))
            begin
              reg331 <= ("q1ETDMDN" <= reg301);
              for (forvar332 = (1'h0); (forvar332 < (2'h2)); forvar332 = (forvar332 + (1'h1)))
                begin
                  reg333 <= (reg239[(4'hd):(2'h3)] ? reg272 : (8'hb8));
                  reg334 <= $unsigned($unsigned($unsigned(($signed(reg293) >> forvar310[(5'h12):(4'h9)]))));
                  reg335 <= $unsigned(reg250);
                  reg336 <= "NVh9wakFCpsp0F";
                  reg337 <= "MqiW9Oeewzq9m8q";
                  reg338 <= (^~(-($unsigned($unsigned(reg295)) >>> reg315)));
                end
              reg339 = (~|reg263[(5'h10):(4'hf)]);
              reg340 <= $unsigned(reg243[(3'h4):(3'h4)]);
              reg341 = (wire288 ?
                  ("2tDf7W72E" || ($unsigned($unsigned(reg290)) | "biGX4Rt8yUsgTEcY9")) : "Tzn3Q7E2smJY1NDV");
              reg342 <= ({(forvar297[(5'h16):(4'hc)] ?
                      {(^reg302), reg271[(1'h0):(1'h0)]} : ((~|wire288) ?
                          (~|reg281) : (^~reg295)))} <<< reg255[(4'hf):(3'h7)]);
            end
          reg343 <= $unsigned(("6hDAQLRwQ6hzrtuNws" << ((7'h40) ?
              "SXs86qrkm" : reg256)));
          for (forvar344 = (1'h0); (forvar344 < (3'h4)); forvar344 = (forvar344 + (1'h1)))
            begin
              for (forvar345 = (1'h0); (forvar345 < (2'h3)); forvar345 = (forvar345 + (1'h1)))
                begin
                  reg346 <= $unsigned((&{((reg269 ^~ reg340) ?
                          $signed(reg308) : reg262[(3'h6):(3'h5)]),
                      (-(reg254 ? (8'ha7) : wire232))}));
                  reg347 <= forvar273[(3'h5):(3'h4)];
                  reg348 <= reg341[(5'h11):(3'h4)];
                  reg349 <= "u1XB2XPew3";
                  reg350 <= reg338[(1'h0):(1'h0)];
                end
              reg351 <= {$signed($unsigned({(reg304 * reg286)})),
                  "2BU36YpCZ7gt"};
              for (forvar352 = (1'h0); (forvar352 < (1'h1)); forvar352 = (forvar352 + (1'h1)))
                begin
                  reg353 = reg245[(4'hc):(4'h8)];
                end
              reg354 <= forvar316[(4'hf):(4'hc)];
            end
          for (forvar355 = (1'h0); (forvar355 < (1'h1)); forvar355 = (forvar355 + (1'h1)))
            begin
              reg356 <= (+(reg340[(2'h3):(2'h3)] ^ "izM1UbOAzJZ5eXN8i1b2eQ"));
              reg357 <= {$unsigned(((~|$unsigned(forvar332)) ?
                      (forvar355[(3'h4):(2'h3)] ?
                          "00GldaXsctsZFD2pd" : reg324[(4'hd):(1'h0)]) : $unsigned("llprxGElP")))};
            end
        end
      reg358 <= (($unsigned($signed("xX6Zpt0rbz7pyhiCi")) ?
              $signed(forvar320) : $unsigned($signed((reg247 ?
                  (8'ha5) : reg279)))) ?
          (~|(~($signed(reg317) ?
              (forvar258 | wire222) : reg263[(4'he):(1'h0)]))) : forvar270);
    end
  always
    @(posedge clk) begin
      for (forvar359 = (1'h0); (forvar359 < (3'h5)); forvar359 = (forvar359 + (1'h1)))
        begin
          for (forvar360 = (1'h0); (forvar360 < (2'h2)); forvar360 = (forvar360 + (1'h1)))
            begin
              for (forvar361 = (1'h0); (forvar361 < (2'h2)); forvar361 = (forvar361 + (1'h1)))
                begin
                  reg362 = $signed(($signed($unsigned("JX")) ?
                      $signed($unsigned((~|forvar234))) : $unsigned((~(reg313 * forvar266)))));
                  reg363 <= "vxY0iMmJFqhPWy3";
                  reg364 = (forvar355[(2'h2):(1'h0)] ~^ "nyUQJduDnWuYl");
                  reg365 = ("lo" ?
                      ((reg318[(3'h4):(2'h3)] * "3X5xfZHceXF") ?
                          reg313[(2'h2):(2'h2)] : $signed($signed(forvar322[(4'ha):(4'ha)]))) : (!($unsigned((!reg271)) ^ reg354[(1'h0):(1'h0)])));
                end
              reg366 <= reg333;
              reg367 <= $unsigned(($signed($unsigned($signed((8'hbf)))) ?
                  {reg261[(2'h2):(2'h2)],
                      (&(reg331 << (8'h9d)))} : ($unsigned((-reg350)) != $unsigned("1aAVx8v6Kb7x"))));
            end
          reg368 <= $signed(reg239);
          reg369 = reg309[(3'h5):(2'h2)];
        end
      reg370 <= ($unsigned($unsigned(reg227[(2'h3):(1'h1)])) ?
          (reg341[(4'h9):(3'h4)] | (~(!"ToN7zORkZrmO81v8"))) : {"zW",
              forvar360[(1'h1):(1'h0)]});
      for (forvar371 = (1'h0); (forvar371 < (1'h1)); forvar371 = (forvar371 + (1'h1)))
        begin
          for (forvar372 = (1'h0); (forvar372 < (3'h5)); forvar372 = (forvar372 + (1'h1)))
            begin
              reg373 <= $unsigned(forvar361[(5'h11):(3'h7)]);
              reg374 <= reg278[(1'h0):(1'h0)];
              reg375 <= $signed("SN3vQTgMuM5XBcewTyKne");
              for (forvar376 = (1'h0); (forvar376 < (2'h2)); forvar376 = (forvar376 + (1'h1)))
                begin
                  reg377 = ((+$signed(reg357[(5'h15):(4'hb)])) < reg348);
                  reg378 = (|wire232);
                  reg379 = (~^((-(~^$unsigned(reg255))) ?
                      $unsigned($unsigned($unsigned((8'hba)))) : reg262));
                end
            end
          for (forvar380 = (1'h0); (forvar380 < (3'h5)); forvar380 = (forvar380 + (1'h1)))
            begin
              reg381 <= ((reg259 + $signed((forvar270 ?
                  (+forvar360) : reg243[(4'ha):(3'h7)]))) < (($signed((forvar257 ?
                          (8'ha3) : reg279)) ?
                      $unsigned(forvar355[(2'h2):(1'h1)]) : reg315) ?
                  (^~reg369) : ($signed((reg341 ?
                      reg334 : forvar330)) != (reg296 != $unsigned(reg319)))));
              reg382 = (reg362 ?
                  (forvar355[(3'h5):(3'h5)] ?
                      (wire221 ?
                          reg289 : $signed((reg300 <= reg287))) : (-$signed(forvar332[(1'h0):(1'h0)]))) : reg281);
              reg383 <= $unsigned({(reg230[(5'h13):(1'h0)] ?
                      (|reg365) : $signed({reg301, reg271}))});
              for (forvar384 = (1'h0); (forvar384 < (1'h1)); forvar384 = (forvar384 + (1'h1)))
                begin
                  reg385 <= $signed("Ol26H3UGbiTdvuYczX");
                  reg386 <= ("GuzSASOBUdscC7UYN0XPPTzO" ?
                      ($signed(reg366) ?
                          (((+reg237) ?
                                  (reg336 ? reg297 : reg346) : (forvar322 ?
                                      reg367 : reg304)) ?
                              {"GQDZ0SS9k7A"} : (^~(forvar322 ?
                                  forvar345 : reg271))) : forvar310[(5'h13):(4'hc)]) : {((reg340[(1'h1):(1'h1)] != "I5IiXaIFpB") ?
                              reg335 : reg331[(4'h9):(1'h1)])});
                  reg387 <= forvar316[(4'hc):(4'ha)];
                  reg388 <= reg374;
                  reg389 <= {"", $unsigned(reg239[(4'he):(3'h6)])};
                end
              if ({"1T387E8i2pq9ozs9"})
                begin
                  reg390 <= ({reg242[(4'hf):(4'h8)],
                          (~|(^~((8'hb7) ? reg260 : forvar352)))} ?
                      reg328[(3'h6):(2'h3)] : reg309);
                  reg391 = reg382;
                  reg392 <= ($unsigned("9ZDcJY") ?
                      $signed((($signed(reg250) << (reg391 && forvar257)) ?
                          reg343[(5'h17):(5'h12)] : $unsigned({reg287}))) : "0oI2DTdIY");
                  reg393 <= $unsigned((~|reg324));
                  reg394 <= {((|"x2qXX43eU1vNa3ypT9OQhBYK") ?
                          reg237[(3'h4):(2'h3)] : (-reg351)),
                      reg301[(3'h6):(1'h1)]};
                  reg395 <= ((~^forvar371) ?
                      $unsigned($unsigned($unsigned((forvar270 ?
                          wire232 : (7'h44))))) : $unsigned((8'ha4)));
                end
              else
                begin
                  reg390 = $unsigned((reg336[(3'h4):(3'h4)] ?
                      (^~reg227[(2'h3):(2'h2)]) : $signed(("aF3YcgzrPYJ6c9dZ61yy3e" <= $signed(reg295)))));
                  reg391 <= (~|$unsigned(reg274[(4'hf):(4'hf)]));
                  reg392 <= $unsigned($unsigned(forvar292));
                  reg393 = ((+(-{$signed((7'h40))})) ?
                      reg247 : {"OFzPkSXrsa6XcCwJLQuxo"});
                  reg394 <= ($unsigned("TR7fW8") ?
                      "u0nBXD2S0V" : ($unsigned((reg323 ?
                              (&(8'ha3)) : wire232[(2'h3):(2'h3)])) ?
                          ($signed("nRSY") & "pblMxobNUkkP") : (~^$signed($signed((8'ha0))))));
                end
            end
          for (forvar396 = (1'h0); (forvar396 < (1'h0)); forvar396 = (forvar396 + (1'h1)))
            begin
              for (forvar397 = (1'h0); (forvar397 < (2'h2)); forvar397 = (forvar397 + (1'h1)))
                begin
                  reg398 <= "6Yaw0d9AgTrHEMv";
                  reg399 <= "5tLiiBwqQ9OWsaXdc";
                  reg400 <= $unsigned((~$signed("hO0q")));
                  reg401 <= forvar332[(1'h0):(1'h0)];
                  reg402 <= reg333;
                end
              reg403 <= (7'h49);
              for (forvar404 = (1'h0); (forvar404 < (2'h2)); forvar404 = (forvar404 + (1'h1)))
                begin
                  reg405 = reg381[(3'h6):(3'h4)];
                  reg406 <= (-"");
                  reg407 <= ("X0X8qvP301ProoJ" ?
                      (|($unsigned($unsigned((8'haf))) ?
                          (forvar282[(2'h3):(1'h0)] + $unsigned(reg255)) : ((wire221 & reg298) <= "SsBMf0Mn7SCb6wD"))) : (wire221 && ($unsigned($signed(forvar316)) ?
                          "8HrcBa" : forvar298)));
                end
            end
          reg408 <= $signed((!(^~$signed((^~reg269)))));
        end
      reg409 <= ($unsigned(("hZyUrWih799128cQLED" >= ($signed((8'h9f)) ~^ $signed(reg327)))) ?
          "xYvAFLMRzEVK2IUD" : $unsigned((|"7XvPRypK3tEP6zLaJu6eo")));
    end
  always
    @(posedge clk) begin
      reg410 = ("1" ? "pWWimsw2o" : "");
    end
  assign wire411 = $signed("aRROy9pS25GfoXWN");
  always
    @(posedge clk) begin
      for (forvar412 = (1'h0); (forvar412 < (2'h3)); forvar412 = (forvar412 + (1'h1)))
        begin
          reg413 <= ($unsigned((reg353 != ("LR1uRGXy6chfKgEsSKBG" ?
              forvar310[(4'he):(1'h0)] : (~reg315)))) - {reg342,
              reg264[(4'hd):(2'h3)]});
          if ($signed(((forvar361[(4'h9):(4'h8)] ?
                  reg363[(4'h9):(2'h3)] : ((reg358 ^~ forvar397) ?
                      "MPXspKR0hehmAbhrtK" : (reg227 ? reg252 : reg362))) ?
              wire232[(3'h4):(2'h3)] : (8'hb8))))
            begin
              reg414 <= reg256[(3'h4):(1'h0)];
              for (forvar415 = (1'h0); (forvar415 < (3'h5)); forvar415 = (forvar415 + (1'h1)))
                begin
                  reg416 <= "MSpQqaLybbweROhlhKo";
                  reg417 <= $signed((reg239[(4'ha):(3'h4)] ?
                      (forvar397 ?
                          "Sg0DKtdQC" : (7'h4d)) : $signed(forvar292)));
                  reg418 <= reg324;
                  reg419 <= (~(-(^$signed($signed(reg374)))));
                  reg420 = "OPOW";
                end
              for (forvar421 = (1'h0); (forvar421 < (2'h3)); forvar421 = (forvar421 + (1'h1)))
                begin
                  reg422 <= $unsigned("Z8c");
                  reg423 <= reg251;
                  reg424 <= "hJAwmNq4F5V0IkstfM9f";
                  reg425 <= $signed("7Q2MyuXRPP7wOtHoPsB");
                  reg426 <= ("wPEeAdB9gBmy" * (-{(reg419[(5'h16):(3'h6)] ?
                          $signed(wire233) : (reg407 && reg422))}));
                end
              reg427 = reg325[(4'hc):(3'h5)];
              reg428 <= $signed(reg413[(3'h7):(3'h5)]);
              reg429 <= reg418[(3'h5):(2'h2)];
            end
          else
            begin
              reg414 <= ("" ? "vuEZJJ42atch" : reg328);
              reg415 = (8'h9c);
            end
          reg430 = reg234[(2'h2):(2'h2)];
          for (forvar431 = (1'h0); (forvar431 < (3'h5)); forvar431 = (forvar431 + (1'h1)))
            begin
              reg432 <= (!($signed(reg398[(3'h7):(3'h5)]) ^~ forvar258[(4'hb):(3'h4)]));
              reg433 = reg309[(4'he):(4'hb)];
              reg434 <= reg370[(1'h1):(1'h1)];
              reg435 <= reg419;
              reg436 <= (&$unsigned(($unsigned((8'hbf)) ?
                  (reg290[(4'ha):(3'h5)] ~^ ((8'h9f) & reg294)) : $signed((reg305 ?
                      reg358 : reg429)))));
            end
        end
      reg437 <= ($signed($signed({(^~reg381)})) << $unsigned((^{"hSJT6Zi9Uc8tRkYc"})));
      reg438 = ($unsigned(((|$signed(reg410)) ^ forvar234)) ?
          $signed(reg377) : (&$signed(reg302[(2'h3):(1'h0)])));
      reg439 = (~$signed((-reg262[(2'h2):(2'h2)])));
    end
  assign wire440 = (reg430 << reg277);
  assign wire441 = ((^~$signed($unsigned(((7'h46) < (8'hbd))))) ?
                       $unsigned(forvar344[(1'h1):(1'h1)]) : ((("npLUbqTy09w8vxIwH4" && "XRlz5BCk") ?
                           ({reg378} ?
                               "yEHbc22oyRQWae36" : (reg238 ?
                                   reg374 : reg416)) : $unsigned((~|(8'hbf)))) >> reg307[(4'h9):(3'h6)]));
  assign wire442 = $signed($signed("DdJ5azJQ74eU"));
  assign wire443 = (~(reg313[(1'h0):(1'h0)] ^~ (8'hb9)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module93
#( parameter param173 = ({(^~(~&(+(8'h9d))))} ? (^~(&(((7'h4d) ? (7'h46) : (7'h41)) ? ((7'h45) ? (7'h48) : (8'hb2)) : (7'h40)))) : ((((~|(7'h45)) + ((8'hb9) << (8'h9e))) > {{(8'ha8), (8'hb2)}}) ? ((!((8'haf) ? (8'haf) : (8'h9c))) >> (((7'h4a) ? (8'h9f) : (7'h4c)) || ((7'h44) - (7'h4e)))) : {(~|(~^(8'ha3)))}))
, parameter param174 = param173 )
(y, clk, wire97, wire96, wire95, wire94);
  output wire [(32'h432):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire97;
  input wire [(4'ha):(1'h0)] wire96;
  input wire signed [(5'h12):(1'h0)] wire95;
  input wire [(4'hd):(1'h0)] wire94;
  wire signed [(5'h12):(1'h0)] wire172;
  reg [(3'h5):(1'h0)] reg171 = (1'h0);
  reg [(4'h9):(1'h0)] reg170 = (1'h0);
  reg [(5'h17):(1'h0)] reg169 = (1'h0);
  reg [(5'h19):(1'h0)] reg168 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg167 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg166 = (1'h0);
  reg [(4'he):(1'h0)] reg165 = (1'h0);
  reg [(5'h17):(1'h0)] reg164 = (1'h0);
  reg [(4'he):(1'h0)] reg163 = (1'h0);
  reg [(5'h14):(1'h0)] forvar162 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar161 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg160 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg159 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire158;
  reg signed [(3'h6):(1'h0)] reg157 = (1'h0);
  wire [(5'h10):(1'h0)] wire156;
  wire signed [(5'h12):(1'h0)] wire155;
  reg signed [(3'h4):(1'h0)] reg154 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg152 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg150 = (1'h0);
  reg [(5'h15):(1'h0)] reg149 = (1'h0);
  reg [(2'h2):(1'h0)] reg148 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar147 = (1'h0);
  reg signed [(4'he):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar145 = (1'h0);
  reg [(3'h7):(1'h0)] reg144 = (1'h0);
  reg [(3'h5):(1'h0)] reg143 = (1'h0);
  reg [(4'he):(1'h0)] reg142 = (1'h0);
  reg [(5'h16):(1'h0)] reg141 = (1'h0);
  reg [(5'h1a):(1'h0)] reg140 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg139 = (1'h0);
  reg [(4'hb):(1'h0)] reg138 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg137 = (1'h0);
  reg [(4'hc):(1'h0)] reg136 = (1'h0);
  reg [(3'h5):(1'h0)] forvar135 = (1'h0);
  reg [(5'h16):(1'h0)] forvar134 = (1'h0);
  reg [(5'h14):(1'h0)] forvar133 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg132 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg131 = (1'h0);
  reg [(5'h15):(1'h0)] reg130 = (1'h0);
  reg [(4'hb):(1'h0)] forvar129 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg127 = (1'h0);
  reg [(5'h13):(1'h0)] reg126 = (1'h0);
  reg [(3'h4):(1'h0)] reg125 = (1'h0);
  reg [(5'h16):(1'h0)] reg124 = (1'h0);
  reg [(4'he):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar122 = (1'h0);
  reg [(5'h17):(1'h0)] reg121 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg120 = (1'h0);
  reg signed [(4'he):(1'h0)] reg119 = (1'h0);
  reg [(5'h14):(1'h0)] reg118 = (1'h0);
  reg [(4'he):(1'h0)] reg117 = (1'h0);
  reg [(4'he):(1'h0)] forvar116 = (1'h0);
  reg [(5'h15):(1'h0)] reg115 = (1'h0);
  reg [(5'h14):(1'h0)] reg114 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg113 = (1'h0);
  reg [(5'h15):(1'h0)] forvar112 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg111 = (1'h0);
  reg [(4'ha):(1'h0)] reg110 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar109 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar108 = (1'h0);
  reg [(4'he):(1'h0)] reg107 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg106 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg105 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg104 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire103;
  wire [(4'hd):(1'h0)] wire102;
  reg signed [(5'h13):(1'h0)] reg101 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar100 = (1'h0);
  wire [(3'h7):(1'h0)] wire99;
  wire [(4'h8):(1'h0)] wire98;
  assign y = {wire172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 forvar162,
                 forvar161,
                 reg160,
                 reg159,
                 wire158,
                 reg157,
                 wire156,
                 wire155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 forvar147,
                 reg146,
                 forvar145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 forvar135,
                 forvar134,
                 forvar133,
                 reg132,
                 reg131,
                 reg130,
                 forvar129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 forvar122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 forvar116,
                 reg115,
                 reg114,
                 reg113,
                 forvar112,
                 reg111,
                 reg110,
                 forvar109,
                 forvar108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 wire103,
                 wire102,
                 reg101,
                 forvar100,
                 wire99,
                 wire98,
                 (1'h0)};
  assign wire98 = $signed(wire96[(3'h5):(2'h2)]);
  assign wire99 = $unsigned(wire95[(5'h12):(5'h10)]);
  always
    @(posedge clk) begin
      for (forvar100 = (1'h0); (forvar100 < (2'h3)); forvar100 = (forvar100 + (1'h1)))
        begin
          reg101 <= wire94[(3'h6):(1'h1)];
        end
    end
  assign wire102 = wire99;
  assign wire103 = ((^~wire94[(2'h3):(1'h0)]) ~^ (wire98[(1'h0):(1'h0)] ?
                       wire99[(2'h2):(1'h1)] : ({wire95} ?
                           (7'h4a) : ((wire99 ? (7'h4d) : forvar100) ?
                               $signed(wire97) : $signed(wire94)))));
  always
    @(posedge clk) begin
      reg104 <= {($signed((wire94[(3'h7):(3'h7)] * forvar100[(3'h4):(2'h2)])) <<< ((wire98 ?
              $signed(wire99) : (forvar100 >>> wire94)) ^~ forvar100))};
      reg105 <= wire98[(2'h3):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg106 <= $unsigned((~^(^(&(wire96 >>> wire103)))));
      reg107 <= ($signed((8'hb5)) != ("iPSONwFf9Y1fUQL" ?
          ($unsigned($signed(wire95)) > ((reg101 ?
              reg101 : forvar100) <= $signed(wire95))) : reg105[(2'h2):(1'h0)]));
      for (forvar108 = (1'h0); (forvar108 < (3'h5)); forvar108 = (forvar108 + (1'h1)))
        begin
          for (forvar109 = (1'h0); (forvar109 < (1'h0)); forvar109 = (forvar109 + (1'h1)))
            begin
              reg110 <= $unsigned((~|(&(+(7'h48)))));
              reg111 <= (!$unsigned({wire102[(4'hc):(3'h5)],
                  "s6iu484TnRTCrypoaAfqbpE"}));
            end
          for (forvar112 = (1'h0); (forvar112 < (3'h4)); forvar112 = (forvar112 + (1'h1)))
            begin
              reg113 <= $signed(wire94);
              reg114 = ((wire96 ?
                  $unsigned(({wire103, wire96} ?
                      reg105[(1'h1):(1'h1)] : $unsigned(reg106))) : wire103[(3'h7):(2'h2)]) ~^ (-$unsigned($unsigned("zNk3JcrM8JAiYnBsCpT"))));
              reg115 <= (((&("xlN4" ~^ wire95)) ?
                  $unsigned("") : ((-$unsigned(wire102)) + (~^forvar109[(2'h3):(2'h2)]))) || wire95);
              for (forvar116 = (1'h0); (forvar116 < (3'h5)); forvar116 = (forvar116 + (1'h1)))
                begin
                  reg117 <= reg101;
                  reg118 = ((|"3C") ?
                      ($unsigned((reg104[(2'h2):(1'h0)] << (+reg104))) << $unsigned(wire103)) : ((reg117[(4'hc):(4'h9)] || "NDUwV1JDY5votuukfIsiq1U") ?
                          "vB0J70ElggmzK41khQBNpQ" : (~{(~|wire103),
                              (reg106 >> reg115)})));
                  reg119 = (($signed($signed((reg110 < (8'ha7)))) != "Q0co") < forvar100[(1'h1):(1'h1)]);
                  reg120 <= forvar116[(4'h8):(1'h0)];
                  reg121 = $unsigned((reg120[(2'h3):(2'h3)] ?
                      forvar116 : $signed((((8'hab) ?
                          wire103 : reg106) * (reg105 ? forvar100 : reg101)))));
                end
              for (forvar122 = (1'h0); (forvar122 < (3'h5)); forvar122 = (forvar122 + (1'h1)))
                begin
                  reg123 <= ((-($unsigned((~^(8'haf))) ?
                          wire99[(2'h2):(1'h1)] : forvar109[(1'h0):(1'h0)])) ?
                      ($signed($signed((8'hbe))) ~^ (("puWBmNOOz33vTRQfGXY1" ?
                              (+wire102) : "vFVBx8WkI8iK9vrCHvCb") ?
                          $unsigned((forvar109 <= forvar100)) : $unsigned(reg115))) : (-(~((reg105 || wire96) ?
                          (wire103 ? reg115 : (7'h4b)) : (&forvar108)))));
                  reg124 <= forvar112[(4'hc):(3'h7)];
                  reg125 <= (reg120 <= (+(reg105[(1'h1):(1'h0)] <<< ((!forvar100) ?
                      (~^reg104) : (~|reg119)))));
                end
              reg126 <= wire96[(3'h6):(2'h2)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg127 = (8'ha4);
      reg128 <= {reg115, reg121[(4'hf):(2'h3)]};
      for (forvar129 = (1'h0); (forvar129 < (1'h1)); forvar129 = (forvar129 + (1'h1)))
        begin
          reg130 <= (!{($unsigned(reg121[(4'hf):(4'hc)]) << wire102),
              ({(reg124 ? (8'hb4) : (7'h4a))} >> ({reg118} & {reg111}))});
          reg131 <= ($signed($signed({$unsigned(wire94)})) && $signed(({((8'h9d) ~^ wire95)} ?
              (8'hae) : "6f8nueuXEmX")));
        end
      reg132 <= $unsigned(reg118[(3'h6):(2'h3)]);
      for (forvar133 = (1'h0); (forvar133 < (1'h0)); forvar133 = (forvar133 + (1'h1)))
        begin
          for (forvar134 = (1'h0); (forvar134 < (3'h4)); forvar134 = (forvar134 + (1'h1)))
            begin
              for (forvar135 = (1'h0); (forvar135 < (2'h2)); forvar135 = (forvar135 + (1'h1)))
                begin
                  reg136 <= $unsigned($unsigned(reg107));
                  reg137 = reg124[(5'h15):(2'h3)];
                  reg138 <= "QiJ";
                end
              reg139 <= (~|wire103[(1'h1):(1'h0)]);
              reg140 <= reg121[(5'h16):(5'h15)];
            end
          reg141 = {{((-(wire99 != wire98)) ?
                      $unsigned(forvar134[(1'h0):(1'h0)]) : reg104[(2'h2):(1'h0)])},
              $unsigned($signed($signed("AoATDFnpcwMAgyB")))};
          reg142 <= ((|(!({wire94,
              reg127} >= "Ny9aEW1WesqxoJ"))) + $unsigned((!((reg111 ?
              wire102 : wire99) != $unsigned(forvar129)))));
          reg143 <= $unsigned((-(+(reg120 ?
              reg110[(3'h7):(3'h4)] : (forvar108 ~^ (8'hac))))));
          reg144 <= (reg125 ?
              (~^(($signed(reg140) ?
                  $signed((7'h40)) : (reg104 + reg113)) <= (~$signed(reg114)))) : (~&((reg106 ?
                      reg117[(2'h3):(1'h0)] : wire99) ?
                  reg123[(3'h5):(2'h3)] : $signed(wire95))));
          for (forvar145 = (1'h0); (forvar145 < (3'h4)); forvar145 = (forvar145 + (1'h1)))
            begin
              reg146 <= (&"g4tXeGoJ");
              for (forvar147 = (1'h0); (forvar147 < (2'h3)); forvar147 = (forvar147 + (1'h1)))
                begin
                  reg148 <= "7c391upk";
                  reg149 <= "c";
                  reg150 = {(wire97 ? $signed((!{reg149})) : forvar108)};
                end
              reg151 <= (reg144[(3'h4):(2'h3)] | $signed((("Ls5IdTgmxMoR0e2K9f" <<< forvar112[(5'h12):(5'h11)]) ?
                  ((reg125 + reg119) || (!(8'hb0))) : $unsigned($unsigned(reg148)))));
              reg152 <= $unsigned("vSNZ");
              reg153 <= ("zhIotZZ6TvYEuQQ" ?
                  $signed(($signed((reg140 ? reg120 : reg130)) ?
                      (~&reg125) : $unsigned($unsigned(reg101)))) : ("0dmMtnToPl0Lh" ?
                      ((forvar133 ?
                          "03Rs" : reg127[(5'h11):(3'h4)]) != (forvar147 << $unsigned((8'ha3)))) : (!$signed(reg130))));
            end
        end
      reg154 <= "mgdoY73sPwotrEdSa9rn6FWiS";
    end
  assign wire155 = ((&((reg141[(3'h5):(3'h5)] == "82XD9QxPHrNI5WvLZlPOoiik") ?
                           reg121[(4'hf):(1'h1)] : ((!reg127) != $signed(reg113)))) ?
                       (~|((|(wire98 ? reg132 : reg153)) ?
                           $signed(reg123[(4'ha):(1'h1)]) : "")) : reg121);
  assign wire156 = reg105;
  always
    @(posedge clk) begin
      reg157 = forvar109[(2'h2):(2'h2)];
    end
  assign wire158 = (&(~^reg105));
  always
    @(posedge clk) begin
      reg159 = $unsigned($unsigned(((!"8CVfLC") ?
          $signed((~^reg146)) : $signed(reg152[(1'h0):(1'h0)]))));
      reg160 = ($unsigned((((reg110 << reg104) * (~(8'hab))) & $unsigned({(7'h43)}))) ?
          "B52uPrDopnIIMk" : forvar135);
      for (forvar161 = (1'h0); (forvar161 < (2'h2)); forvar161 = (forvar161 + (1'h1)))
        begin
          for (forvar162 = (1'h0); (forvar162 < (1'h0)); forvar162 = (forvar162 + (1'h1)))
            begin
              reg163 <= $unsigned(((~^(~&$unsigned((8'ha9)))) ?
                  ((~&(&forvar108)) >>> reg104) : $signed((-(wire96 ?
                      (8'hb0) : reg153)))));
              if ((^($unsigned((reg114[(4'hd):(1'h0)] ?
                  ((7'h40) & (8'ha7)) : $signed(wire103))) + ("X36vkOiY0hkAA0yVQHS" << "8XsJByqPMWqec9blzP"))))
                begin
                  reg164 = wire155[(5'h11):(4'hc)];
                  reg165 <= $signed($signed(forvar122));
                  reg166 = (~|(reg151 ?
                      "ANPZihBqy2iKCNI1Pko" : (|"N69xaSqZd")));
                end
              else
                begin
                  reg164 <= reg111;
                end
              reg167 <= $signed((("DhxQyQ7HaBS" || forvar135) ?
                  (!(forvar108 & (forvar109 ? (8'hb3) : reg104))) : (8'h9e)));
            end
          reg168 <= reg127;
          reg169 <= $signed((^~"VQMOZGHfnFgprxo"));
        end
      reg170 <= reg169;
      reg171 <= $signed($signed(((&{forvar134, reg106}) ?
          $unsigned(reg165[(3'h5):(1'h0)]) : $signed(wire155[(4'ha):(3'h7)]))));
    end
  assign wire172 = (^(|((reg168[(3'h6):(3'h6)] == $unsigned(wire95)) && (^(|forvar133)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4117  (y, clk, wire4121, wire4120, wire4119, wire4118);
  output wire [(32'h3f9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire4121;
  input wire signed [(5'h18):(1'h0)] wire4120;
  input wire [(5'h13):(1'h0)] wire4119;
  input wire [(5'h19):(1'h0)] wire4118;
  reg signed [(3'h5):(1'h0)] reg4187 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire4186;
  wire [(5'h11):(1'h0)] wire4185;
  wire [(4'hd):(1'h0)] wire4184;
  wire [(5'h19):(1'h0)] wire4183;
  wire [(4'he):(1'h0)] wire4182;
  wire signed [(5'h18):(1'h0)] wire4181;
  wire signed [(4'ha):(1'h0)] wire4180;
  wire signed [(5'h19):(1'h0)] wire4179;
  reg [(5'h11):(1'h0)] reg4178 = (1'h0);
  reg [(5'h11):(1'h0)] reg4177 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4176 = (1'h0);
  reg [(5'h16):(1'h0)] reg4175 = (1'h0);
  reg [(3'h4):(1'h0)] reg4174 = (1'h0);
  reg [(4'hb):(1'h0)] reg4173 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4172 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg4171 = (1'h0);
  reg [(5'h11):(1'h0)] reg4170 = (1'h0);
  reg [(5'h14):(1'h0)] forvar4169 = (1'h0);
  reg [(5'h11):(1'h0)] reg4168 = (1'h0);
  reg [(5'h15):(1'h0)] reg4167 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4166 = (1'h0);
  reg [(4'he):(1'h0)] reg4165 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg4164 = (1'h0);
  reg [(5'h11):(1'h0)] reg4163 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4162 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4161 = (1'h0);
  reg [(3'h5):(1'h0)] reg4160 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire4159;
  reg [(5'h10):(1'h0)] reg4158 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4157 = (1'h0);
  wire [(5'h15):(1'h0)] wire4156;
  reg [(5'h14):(1'h0)] reg4155 = (1'h0);
  reg [(3'h5):(1'h0)] reg4154 = (1'h0);
  wire [(5'h19):(1'h0)] wire4153;
  wire [(4'h8):(1'h0)] wire4152;
  wire [(2'h3):(1'h0)] wire4151;
  reg signed [(5'h13):(1'h0)] reg4150 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg4149 = (1'h0);
  reg [(5'h18):(1'h0)] reg4148 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4147 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg4146 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg4145 = (1'h0);
  reg [(4'hf):(1'h0)] reg4144 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4143 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar4142 = (1'h0);
  reg [(5'h15):(1'h0)] reg4141 = (1'h0);
  reg [(4'h8):(1'h0)] reg4140 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg4139 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire4138;
  wire [(5'h12):(1'h0)] wire4137;
  wire [(5'h13):(1'h0)] wire4136;
  reg signed [(5'h19):(1'h0)] reg4135 = (1'h0);
  reg [(5'h11):(1'h0)] reg4134 = (1'h0);
  reg [(5'h11):(1'h0)] reg4133 = (1'h0);
  reg [(5'h15):(1'h0)] reg4132 = (1'h0);
  wire [(2'h3):(1'h0)] wire4131;
  wire [(5'h10):(1'h0)] wire4130;
  reg [(3'h4):(1'h0)] reg4129 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg4128 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4127 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4126 = (1'h0);
  reg [(5'h17):(1'h0)] forvar4125 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4124 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4123 = (1'h0);
  reg [(4'h8):(1'h0)] reg4122 = (1'h0);
  assign y = {reg4187,
                 wire4186,
                 wire4185,
                 wire4184,
                 wire4183,
                 wire4182,
                 wire4181,
                 wire4180,
                 wire4179,
                 reg4178,
                 reg4177,
                 reg4176,
                 reg4175,
                 reg4174,
                 reg4173,
                 forvar4172,
                 reg4171,
                 reg4170,
                 forvar4169,
                 reg4168,
                 reg4167,
                 reg4166,
                 reg4165,
                 reg4164,
                 reg4163,
                 reg4162,
                 forvar4161,
                 reg4160,
                 wire4159,
                 reg4158,
                 reg4157,
                 wire4156,
                 reg4155,
                 reg4154,
                 wire4153,
                 wire4152,
                 wire4151,
                 reg4150,
                 reg4149,
                 reg4148,
                 reg4147,
                 reg4146,
                 reg4145,
                 reg4144,
                 reg4143,
                 forvar4142,
                 reg4141,
                 reg4140,
                 reg4139,
                 wire4138,
                 wire4137,
                 wire4136,
                 reg4135,
                 reg4134,
                 reg4133,
                 reg4132,
                 wire4131,
                 wire4130,
                 reg4129,
                 reg4128,
                 reg4127,
                 reg4126,
                 forvar4125,
                 reg4124,
                 reg4123,
                 reg4122,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg4122 = {$unsigned("JGA82Qtq4tPk8XJrtBGwLrVVs")};
      reg4123 = wire4119;
      reg4124 = wire4118[(1'h0):(1'h0)];
      for (forvar4125 = (1'h0); (forvar4125 < (1'h1)); forvar4125 = (forvar4125 + (1'h1)))
        begin
          reg4126 = wire4120[(1'h0):(1'h0)];
          reg4127 = reg4124;
          reg4128 = (wire4119 ?
              (wire4119[(4'hb):(3'h4)] ?
                  (^((|forvar4125) ?
                      (8'h9e) : wire4119)) : wire4119) : $unsigned($signed((reg4126[(2'h3):(2'h3)] ?
                  wire4119[(5'h13):(5'h12)] : $unsigned(reg4127)))));
          reg4129 <= $unsigned(wire4118[(4'h8):(2'h2)]);
        end
    end
  assign wire4130 = wire4121;
  assign wire4131 = $signed(({(((8'hb0) == (8'hb9)) >> "d"),
                            $unsigned((&(8'hb6)))} ?
                        ("3v6c" >= (~&reg4129[(2'h2):(1'h0)])) : (&reg4123[(3'h6):(2'h3)])));
  always
    @(posedge clk) begin
      reg4132 <= reg4123[(2'h2):(1'h0)];
      reg4133 <= (($signed(reg4132[(3'h4):(2'h2)]) >= wire4121) | "KaxvFG1u7P7cZ8KuWk8I");
      reg4134 <= reg4132[(3'h4):(3'h4)];
      reg4135 <= $signed({("46l" - $signed({wire4120}))});
    end
  assign wire4136 = reg4122[(3'h7):(2'h3)];
  assign wire4137 = $unsigned(($signed((wire4120 ?
                            ((8'ha1) && reg4134) : (reg4129 >> reg4123))) ?
                        reg4134 : ($unsigned("zncak1Ph3zB") & $unsigned((reg4132 ?
                            reg4122 : wire4118)))));
  assign wire4138 = (reg4123 ?
                        (-(((|(8'ha9)) <<< ((8'hbd) ? (7'h4c) : reg4126)) ?
                            "f6c3BFJ" : ((&reg4133) ?
                                $signed((8'haf)) : (wire4137 ?
                                    forvar4125 : reg4135)))) : $unsigned(wire4136));
  always
    @(posedge clk) begin
      reg4139 <= {reg4129};
      if (("bVcdEnnXklplrFkkDM9Eni1" ~^ forvar4125))
        begin
          reg4140 <= ((("" - reg4133[(4'hb):(1'h1)]) ^~ wire4137[(5'h11):(4'hc)]) ?
              reg4133[(2'h3):(1'h0)] : (!(8'hab)));
          reg4141 <= $signed(wire4118[(4'ha):(3'h5)]);
          for (forvar4142 = (1'h0); (forvar4142 < (2'h3)); forvar4142 = (forvar4142 + (1'h1)))
            begin
              reg4143 <= ((~$unsigned(reg4139[(3'h7):(2'h2)])) ?
                  reg4127[(2'h2):(2'h2)] : (~reg4126[(2'h2):(1'h0)]));
              reg4144 <= reg4123;
            end
          reg4145 <= "7pdfggOoV1UPit0u0meRyS98";
          reg4146 <= reg4132[(5'h11):(4'h8)];
        end
      else
        begin
          reg4140 <= $signed("1FrffayIPiV4B0wP3N2Xs3I");
        end
      reg4147 <= reg4123[(2'h3):(2'h2)];
      reg4148 <= ($signed("PTeWngamHFiJu") > $unsigned({$signed(((8'hb4) * wire4118)),
          ($signed(reg4134) ? $signed(reg4135) : $unsigned(reg4140))}));
      reg4149 <= {(~"pHuZdI0lc51lksD")};
      reg4150 = {reg4140[(3'h4):(2'h2)], reg4149[(4'h9):(3'h5)]};
    end
  assign wire4151 = (^~$unsigned($unsigned(wire4119[(4'hb):(3'h4)])));
  assign wire4152 = "S378yp0gutZSzgiYhPU7G";
  assign wire4153 = reg4122[(3'h7):(1'h0)];
  always
    @(posedge clk) begin
      reg4154 <= reg4148[(1'h0):(1'h0)];
      reg4155 = $signed(wire4130);
    end
  assign wire4156 = (|reg4133);
  always
    @(posedge clk) begin
      reg4157 <= "xnJJTQT5z";
      reg4158 <= {$signed($unsigned((!{(7'h4d)})))};
    end
  assign wire4159 = reg4135[(3'h6):(3'h5)];
  always
    @(posedge clk) begin
      reg4160 <= "Dp";
      for (forvar4161 = (1'h0); (forvar4161 < (1'h1)); forvar4161 = (forvar4161 + (1'h1)))
        begin
          reg4162 = "PRY";
          reg4163 <= ((|reg4127[(4'h9):(4'h8)]) + ($signed(wire4121[(2'h2):(1'h0)]) - (8'haa)));
          reg4164 <= (^~(($signed({reg4140, (8'ha1)}) ?
              "IVB3sVihH2Vz" : $signed("APucDWoBRzEGw")) << "3w7vP2LTiVi4gzncL4L8eKL"));
          reg4165 = (|{reg4143[(5'h11):(4'he)]});
        end
      reg4166 <= {reg4124[(3'h5):(3'h4)]};
      reg4167 = (^"d5b");
      reg4168 = {$unsigned(wire4137)};
    end
  always
    @(posedge clk) begin
      for (forvar4169 = (1'h0); (forvar4169 < (2'h2)); forvar4169 = (forvar4169 + (1'h1)))
        begin
          reg4170 <= (7'h4b);
          reg4171 <= ({{{(~|reg4146), reg4162[(3'h4):(1'h1)]},
                  wire4120}} && "queRHaobB7Iu0tKB3rDaf8f");
          for (forvar4172 = (1'h0); (forvar4172 < (3'h5)); forvar4172 = (forvar4172 + (1'h1)))
            begin
              reg4173 <= reg4140;
              reg4174 <= $signed(reg4154);
              reg4175 <= ((reg4157[(2'h3):(1'h1)] > ({$signed(reg4163),
                      (!wire4120)} - $signed((reg4133 >= reg4157)))) ?
                  $signed(forvar4161[(3'h6):(2'h2)]) : $signed("Lq9qQvugEz5wXGGEs"));
              reg4176 <= wire4119;
            end
          reg4177 = "d2U0MAiUA5BDyNCc";
          reg4178 = reg4162;
        end
    end
  assign wire4179 = "DQQ";
  assign wire4180 = "1kW1O9";
  assign wire4181 = reg4127[(2'h3):(1'h1)];
  assign wire4182 = $signed($signed($unsigned((~&reg4123))));
  assign wire4183 = (8'hba);
  assign wire4184 = $unsigned((({reg4122, reg4170[(4'hf):(4'hd)]} ?
                            "98wO1AmmLTdhBg4fTt13" : {(reg4133 <<< forvar4169)}) ?
                        {("H" ? (&reg4135) : $unsigned(reg4124)),
                            $unsigned({reg4133,
                                forvar4172})} : (("ALRqwyTB06CuYyxhetDh" == $signed(wire4179)) + $signed(((7'h4b) ^ reg4166)))));
  assign wire4185 = ("E0YD3rEZoT4hhsDhoIZCkSFnc" ^~ {{"tMY52FGdOA"}});
  assign wire4186 = (!$unsigned(reg4122));
  always
    @(posedge clk) begin
      reg4187 <= $unsigned(({forvar4142[(5'h14):(4'h9)]} ^ ((~&"Oz8yL") ?
          "" : $unsigned((7'h42)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4024  (y, clk, wire4029, wire4028, wire4027, wire4026, wire4025);
  output wire [(32'h45a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire4029;
  input wire signed [(4'hc):(1'h0)] wire4028;
  input wire [(5'h14):(1'h0)] wire4027;
  input wire signed [(3'h4):(1'h0)] wire4026;
  input wire signed [(4'h8):(1'h0)] wire4025;
  reg [(4'ha):(1'h0)] reg4113 = (1'h0);
  wire [(2'h2):(1'h0)] wire4112;
  reg [(4'he):(1'h0)] reg4111 = (1'h0);
  reg [(4'h8):(1'h0)] reg4110 = (1'h0);
  reg [(2'h3):(1'h0)] reg4109 = (1'h0);
  reg [(5'h13):(1'h0)] reg4108 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4107 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4106 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire4105;
  reg [(3'h7):(1'h0)] reg4104 = (1'h0);
  reg [(3'h7):(1'h0)] reg4103 = (1'h0);
  reg [(4'hf):(1'h0)] reg4102 = (1'h0);
  reg [(3'h7):(1'h0)] reg4101 = (1'h0);
  reg [(5'h17):(1'h0)] reg4100 = (1'h0);
  reg [(2'h2):(1'h0)] reg4099 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4098 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar4097 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar4096 = (1'h0);
  reg [(3'h7):(1'h0)] reg4095 = (1'h0);
  reg [(4'hc):(1'h0)] reg4094 = (1'h0);
  reg [(2'h3):(1'h0)] reg4093 = (1'h0);
  reg [(3'h5):(1'h0)] reg4092 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4091 = (1'h0);
  reg [(4'hb):(1'h0)] reg4090 = (1'h0);
  reg [(5'h12):(1'h0)] forvar4089 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4088 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4087 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire4086;
  reg signed [(4'hf):(1'h0)] reg4085 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4084 = (1'h0);
  reg [(5'h12):(1'h0)] reg4083 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg4082 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar4081 = (1'h0);
  reg [(4'hf):(1'h0)] reg4080 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4079 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4078 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg4077 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg4076 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire4075;
  wire [(4'hd):(1'h0)] wire4074;
  reg [(4'he):(1'h0)] reg4073 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4072 = (1'h0);
  reg [(4'hb):(1'h0)] reg4071 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4070 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4069 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4068 = (1'h0);
  reg [(5'h17):(1'h0)] reg4067 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4066 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4065 = (1'h0);
  reg [(5'h12):(1'h0)] reg4064 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4063 = (1'h0);
  reg [(5'h14):(1'h0)] reg4062 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar4061 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg4060 = (1'h0);
  reg [(4'hc):(1'h0)] reg4059 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg4058 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4057 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4056 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4055 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4054 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire4053;
  wire [(4'hf):(1'h0)] wire4052;
  reg signed [(3'h7):(1'h0)] reg4051 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg4050 = (1'h0);
  reg [(3'h7):(1'h0)] reg4049 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg4048 = (1'h0);
  reg [(4'h9):(1'h0)] reg4047 = (1'h0);
  reg [(5'h1a):(1'h0)] reg4046 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg4045 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4044 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4043 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg4042 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4041 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire4040;
  reg signed [(5'h12):(1'h0)] reg4039 = (1'h0);
  reg [(2'h3):(1'h0)] reg4038 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg4037 = (1'h0);
  reg [(5'h1a):(1'h0)] reg4036 = (1'h0);
  reg [(5'h17):(1'h0)] reg4035 = (1'h0);
  reg [(3'h6):(1'h0)] reg4034 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar4033 = (1'h0);
  reg [(3'h4):(1'h0)] reg4032 = (1'h0);
  reg [(4'h9):(1'h0)] reg4031 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg4030 = (1'h0);
  assign y = {reg4113,
                 wire4112,
                 reg4111,
                 reg4110,
                 reg4109,
                 reg4108,
                 reg4107,
                 reg4106,
                 wire4105,
                 reg4104,
                 reg4103,
                 reg4102,
                 reg4101,
                 reg4100,
                 reg4099,
                 reg4098,
                 forvar4097,
                 forvar4096,
                 reg4095,
                 reg4094,
                 reg4093,
                 reg4092,
                 forvar4091,
                 reg4090,
                 forvar4089,
                 reg4088,
                 reg4087,
                 wire4086,
                 reg4085,
                 reg4084,
                 reg4083,
                 reg4082,
                 forvar4081,
                 reg4080,
                 reg4079,
                 reg4078,
                 reg4077,
                 reg4076,
                 wire4075,
                 wire4074,
                 reg4073,
                 reg4072,
                 reg4071,
                 reg4070,
                 reg4069,
                 forvar4068,
                 reg4067,
                 reg4066,
                 reg4065,
                 reg4064,
                 reg4063,
                 reg4062,
                 forvar4061,
                 reg4060,
                 reg4059,
                 reg4058,
                 forvar4057,
                 reg4056,
                 forvar4055,
                 reg4054,
                 wire4053,
                 wire4052,
                 reg4051,
                 reg4050,
                 reg4049,
                 reg4048,
                 reg4047,
                 reg4046,
                 reg4045,
                 forvar4044,
                 reg4043,
                 reg4042,
                 reg4041,
                 wire4040,
                 reg4039,
                 reg4038,
                 reg4037,
                 reg4036,
                 reg4035,
                 reg4034,
                 forvar4033,
                 reg4032,
                 reg4031,
                 reg4030,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg4030 = "KzUoYhyW";
      reg4031 <= "fdDOJbpEzzmquBxH9Z";
      reg4032 <= (!wire4025);
      for (forvar4033 = (1'h0); (forvar4033 < (2'h2)); forvar4033 = (forvar4033 + (1'h1)))
        begin
          reg4034 = $unsigned($signed($signed("Thf25Y")));
          reg4035 = $unsigned($unsigned((8'ha8)));
          reg4036 <= (((((~(8'h9f)) ?
                  reg4034 : wire4026[(3'h4):(3'h4)]) >>> (~&(+wire4028))) || reg4032) ?
              $unsigned(($unsigned(((8'hb1) ?
                  (8'hbb) : wire4025)) <<< ((~|wire4027) < ((7'h47) ?
                  wire4026 : (8'hbf))))) : wire4026[(2'h3):(1'h0)]);
          reg4037 = (($unsigned((reg4034[(1'h1):(1'h1)] ?
                      "83oLNoEoABn6" : forvar4033)) ?
                  (~&(8'h9d)) : reg4030) ?
              ($signed($unsigned((reg4034 ?
                  reg4030 : wire4027))) ^~ $signed($signed(wire4029[(1'h1):(1'h1)]))) : ((reg4035 ?
                      wire4029 : reg4036[(4'hd):(2'h2)]) ?
                  ((|(!reg4030)) ~^ {(~reg4036),
                      (wire4029 << wire4029)}) : $signed("1hWrufRH0pGYymhQPNXW")));
        end
      reg4038 = wire4028[(3'h5):(1'h1)];
      reg4039 <= reg4035;
    end
  assign wire4040 = $unsigned("tJnueDngnrF95roHVfGrC");
  always
    @(posedge clk) begin
      reg4041 = $unsigned((("vy7" || reg4036) ?
          $unsigned(wire4040) : reg4034[(3'h6):(1'h1)]));
      reg4042 <= $unsigned(reg4035[(4'hd):(4'hb)]);
    end
  always
    @(posedge clk) begin
      reg4043 = $signed("6NpoCTGweCTPqc5gCGDt");
      for (forvar4044 = (1'h0); (forvar4044 < (2'h3)); forvar4044 = (forvar4044 + (1'h1)))
        begin
          reg4045 <= "vO";
          reg4046 <= reg4041;
          reg4047 <= ("6asfP" ? $unsigned("") : $signed(wire4028));
        end
      reg4048 <= (7'h4d);
      reg4049 <= (($unsigned($signed(wire4029)) ? "7" : "temGkosHh8ro8m") ?
          ("onKWx1xqdpUfwvHBNb9ikLkIv" ?
              reg4037 : {(wire4028[(1'h1):(1'h0)] * reg4037),
                  "mZS"}) : reg4043);
      reg4050 = reg4037;
      reg4051 <= "";
    end
  assign wire4052 = $signed(reg4049);
  assign wire4053 = "t4CRsmoEa";
  always
    @(posedge clk) begin
      reg4054 <= (~($unsigned({(reg4039 * wire4052)}) ?
          "9yIVCu" : $unsigned((+$signed(reg4034)))));
      for (forvar4055 = (1'h0); (forvar4055 < (3'h4)); forvar4055 = (forvar4055 + (1'h1)))
        begin
          reg4056 <= reg4038;
          for (forvar4057 = (1'h0); (forvar4057 < (2'h2)); forvar4057 = (forvar4057 + (1'h1)))
            begin
              reg4058 <= ($unsigned(reg4036[(5'h13):(5'h12)]) ?
                  reg4041[(4'he):(2'h3)] : ($unsigned((!(^wire4052))) && {(^~(wire4040 ?
                          wire4029 : reg4041))}));
              reg4059 <= "t36ZkJ7Wei7ey1YhNab8";
              reg4060 <= $signed(reg4042[(4'hc):(4'ha)]);
              for (forvar4061 = (1'h0); (forvar4061 < (3'h4)); forvar4061 = (forvar4061 + (1'h1)))
                begin
                  reg4062 = reg4042;
                  reg4063 = ((((+(+(8'hbc))) & ((reg4039 >= reg4054) ~^ $unsigned(reg4051))) ?
                          $unsigned({(reg4050 > reg4062),
                              (reg4045 | reg4036)}) : $unsigned("")) ?
                      "5e" : (^~($unsigned((~wire4026)) ?
                          "dogQS7z5X4OyixsAtHcKf3" : ($unsigned(wire4053) & (~reg4050)))));
                  reg4064 <= (~reg4056);
                  reg4065 = reg4048[(1'h1):(1'h0)];
                  reg4066 <= (($unsigned(({reg4037} ?
                          forvar4044[(1'h1):(1'h1)] : (reg4037 ?
                              reg4037 : reg4043))) ?
                      $unsigned(($signed(reg4058) ?
                          (-reg4034) : (!reg4049))) : (~^$unsigned("UC"))) && (wire4026 ?
                      {$signed("WDNVxiiEZLI5qMz32")} : wire4053[(5'h13):(5'h13)]));
                  reg4067 <= reg4046;
                end
              for (forvar4068 = (1'h0); (forvar4068 < (1'h0)); forvar4068 = (forvar4068 + (1'h1)))
                begin
                  reg4069 <= (&$signed(reg4051));
                  reg4070 <= $signed((8'hbf));
                end
            end
          reg4071 = (^($signed($unsigned((forvar4044 ? reg4047 : reg4056))) ?
              $signed(forvar4061) : $unsigned(reg4059[(4'h9):(3'h7)])));
          reg4072 <= reg4067;
          reg4073 <= $signed($signed("rt"));
        end
    end
  assign wire4074 = $signed({{"J644kJldq6Kk4lnDbNrVsndQ",
                            $unsigned((~^reg4048))}});
  assign wire4075 = "NR38";
  always
    @(posedge clk) begin
      reg4076 <= $signed((($signed($signed(wire4028)) <<< {(wire4053 ^ reg4039)}) << reg4060));
      reg4077 <= ($signed((reg4067[(4'ha):(1'h1)] & (~^$signed(reg4038)))) ~^ (reg4058 - $unsigned(($unsigned(reg4032) || {reg4045}))));
      reg4078 = ((($unsigned({wire4025}) ? reg4037 : wire4074) ?
          {(~^{(8'hb0)})} : $signed("967J97KBz20vJs")) + $unsigned(reg4077));
      reg4079 <= (reg4054[(2'h3):(1'h0)] ^~ {forvar4055[(4'hb):(4'hb)],
          {("g2VrIz8aKndkZJBvWvh7VRc" && reg4031)}});
      reg4080 = "cpbvuWunoafPGB07NLoG";
      for (forvar4081 = (1'h0); (forvar4081 < (2'h2)); forvar4081 = (forvar4081 + (1'h1)))
        begin
          reg4082 = (|("z4uWy8XM24n" ?
              reg4046 : (~^$unsigned((reg4077 ^ reg4045)))));
          reg4083 = "wKiq3ImZnXdDDhhaELiXJYwT";
          reg4084 <= $signed($signed($unsigned((+$unsigned(forvar4081)))));
        end
    end
  always
    @(posedge clk) begin
      reg4085 <= $signed(($signed(($unsigned(reg4067) ?
              {forvar4044} : $signed(reg4056))) ?
          (!wire4053[(4'hc):(4'hb)]) : "RqLvRGIPr"));
    end
  assign wire4086 = $unsigned($signed(($unsigned("iUQ1U0BJ") ?
                        forvar4081[(5'h10):(3'h5)] : ("MKTsPEoqe5xE93TEbYDNVxEWz" ?
                            (reg4059 || reg4048) : reg4060[(4'hf):(4'he)]))));
  always
    @(posedge clk) begin
      reg4087 = $signed(reg4050);
      reg4088 <= {((~|((reg4060 ? wire4074 : reg4064) ?
              reg4049[(3'h5):(1'h1)] : (reg4070 >= forvar4068))) <<< (^~{(reg4065 <<< reg4031)})),
          $unsigned((("w3CKr" ~^ $signed(reg4073)) == (|"0LRuY0KTe")))};
      for (forvar4089 = (1'h0); (forvar4089 < (3'h4)); forvar4089 = (forvar4089 + (1'h1)))
        begin
          reg4090 = $unsigned($signed((wire4052 - reg4041[(4'hb):(4'ha)])));
          for (forvar4091 = (1'h0); (forvar4091 < (2'h3)); forvar4091 = (forvar4091 + (1'h1)))
            begin
              reg4092 <= "k1HmSdbmFINFUl";
              reg4093 = wire4029;
              reg4094 = "ownpGtDahv9SWK2Bk";
              reg4095 <= reg4087;
            end
          for (forvar4096 = (1'h0); (forvar4096 < (1'h0)); forvar4096 = (forvar4096 + (1'h1)))
            begin
              for (forvar4097 = (1'h0); (forvar4097 < (3'h4)); forvar4097 = (forvar4097 + (1'h1)))
                begin
                  reg4098 <= (((+wire4086) * (^(~^$unsigned(reg4038)))) ^~ (!$unsigned(("X" <= (~&wire4075)))));
                  reg4099 <= $unsigned("hLeKyfv0NoMJ");
                end
              reg4100 <= "lJtcIY8uJuS0J8R1k0lE";
              reg4101 <= "QMshmxgfBJfS3GAoTCkYrq";
              reg4102 <= (~^$unsigned("7hYpeOLrGbb"));
              reg4103 <= wire4052;
            end
          reg4104 <= $signed("");
        end
    end
  assign wire4105 = forvar4033;
  always
    @(posedge clk) begin
      reg4106 <= "5tR59dXxTzbPH7ssgzD";
      reg4107 <= $signed((~&$signed(($unsigned(forvar4091) ?
          $signed(reg4054) : "YARKv"))));
      reg4108 <= "Ot5cgQdDVXcqgd0WxX14CfVG9";
      reg4109 <= {{{(-reg4080[(3'h4):(2'h3)]), (|$signed(reg4069))},
              $unsigned(((reg4032 == forvar4097) << (|reg4070)))}};
      reg4110 <= $signed($signed($signed("FL1ZpxnTEqWwf3rht")));
      reg4111 <= "SGi7";
    end
  assign wire4112 = (!"zVATG6XH0pDK94B8LmOcOJKH");
  always
    @(posedge clk) begin
      reg4113 <= "ytbWWnzeP";
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3981  (y, clk, wire3985, wire3984, wire3983, wire3982);
  output wire [(32'h14f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire3985;
  input wire signed [(4'ha):(1'h0)] wire3984;
  input wire [(5'h12):(1'h0)] wire3983;
  input wire signed [(5'h1a):(1'h0)] wire3982;
  wire [(5'h18):(1'h0)] wire4005;
  reg [(5'h19):(1'h0)] reg4004 = (1'h0);
  reg [(5'h17):(1'h0)] reg4003 = (1'h0);
  reg [(3'h7):(1'h0)] reg4002 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg4001 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar4000 = (1'h0);
  reg [(5'h19):(1'h0)] reg3999 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3998 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3997 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3996 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar3995 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3994 = (1'h0);
  reg [(5'h13):(1'h0)] forvar3993 = (1'h0);
  reg [(5'h14):(1'h0)] reg3992 = (1'h0);
  reg [(5'h13):(1'h0)] forvar3991 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3990 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3989 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3988 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3987 = (1'h0);
  reg [(4'he):(1'h0)] reg3986 = (1'h0);
  assign y = {wire4005,
                 reg4004,
                 reg4003,
                 reg4002,
                 reg4001,
                 forvar4000,
                 reg3999,
                 reg3998,
                 reg3997,
                 reg3996,
                 forvar3995,
                 reg3994,
                 forvar3993,
                 reg3992,
                 forvar3991,
                 reg3990,
                 forvar3989,
                 reg3988,
                 reg3987,
                 reg3986,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg3986 = wire3983[(3'h6):(3'h6)];
      reg3987 = $signed((~^(~$unsigned("y5DwEE"))));
    end
  always
    @(posedge clk) begin
      reg3988 <= $signed(wire3982[(2'h2):(2'h2)]);
    end
  always
    @(posedge clk) begin
      for (forvar3989 = (1'h0); (forvar3989 < (2'h2)); forvar3989 = (forvar3989 + (1'h1)))
        begin
          reg3990 = $signed($unsigned(wire3983[(5'h10):(4'hd)]));
        end
      for (forvar3991 = (1'h0); (forvar3991 < (3'h4)); forvar3991 = (forvar3991 + (1'h1)))
        begin
          reg3992 = $unsigned(wire3985);
          for (forvar3993 = (1'h0); (forvar3993 < (2'h3)); forvar3993 = (forvar3993 + (1'h1)))
            begin
              reg3994 <= forvar3993;
              for (forvar3995 = (1'h0); (forvar3995 < (3'h4)); forvar3995 = (forvar3995 + (1'h1)))
                begin
                  reg3996 <= reg3986[(4'hc):(4'hc)];
                  reg3997 <= "3fIssXANheiZb8Y7Qy1vwf";
                end
              reg3998 = $unsigned(reg3992[(4'h8):(3'h5)]);
            end
          reg3999 <= wire3985[(2'h2):(1'h0)];
        end
      for (forvar4000 = (1'h0); (forvar4000 < (2'h2)); forvar4000 = (forvar4000 + (1'h1)))
        begin
          reg4001 = reg3999[(4'hb):(3'h4)];
          reg4002 <= forvar3991;
          reg4003 = (~(~|$unsigned(forvar3991)));
        end
      reg4004 <= (7'h40);
    end
  assign wire4005 = (^(~(((reg3986 ? reg4002 : forvar3995) ?
                        reg4003 : (reg4004 ?
                            forvar3991 : forvar3989)) & ({reg4001} >>> (reg4001 ?
                        (8'ha4) : reg3986)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3696
#( parameter param3975 = ((|(~|((~|(7'h4d)) | (&(8'ha8))))) << (((((7'h42) ? (7'h40) : (7'h46)) > {(8'hb7), (8'hbf)}) ? ((-(8'hbd)) ? {(8'hba)} : ((8'ha6) >>> (7'h4a))) : ({(8'hb2)} ? {(8'hbf)} : {(8'hb8)})) ? (+(((8'hba) ? (8'hb2) : (7'h49)) ? (8'hb1) : (^~(8'hbf)))) : {(((8'ha4) & (8'hb8)) ? (8'hb8) : ((8'ha4) || (8'hbd))), {(8'ha6), ((8'ha9) ? (8'ha6) : (7'h4b))}}))
, parameter param3976 = ((~(^(~^param3975))) == (-(+(-(~|param3975))))) )
(y, clk, wire3701, wire3700, wire3699, wire3698, wire3697);
  output wire [(32'hf4f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire3701;
  input wire signed [(3'h4):(1'h0)] wire3700;
  input wire signed [(4'he):(1'h0)] wire3699;
  input wire signed [(5'h1a):(1'h0)] wire3698;
  input wire signed [(4'he):(1'h0)] wire3697;
  reg [(5'h14):(1'h0)] reg3974 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3973 = (1'h0);
  reg [(5'h19):(1'h0)] reg3972 = (1'h0);
  reg [(5'h17):(1'h0)] reg3971 = (1'h0);
  reg [(5'h11):(1'h0)] forvar3970 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3969 = (1'h0);
  reg [(4'he):(1'h0)] forvar3968 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3967 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3966 = (1'h0);
  reg [(3'h6):(1'h0)] reg3965 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3964 = (1'h0);
  reg [(4'hf):(1'h0)] reg3963 = (1'h0);
  reg [(5'h15):(1'h0)] forvar3962 = (1'h0);
  reg [(5'h16):(1'h0)] reg3961 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3960 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3959 = (1'h0);
  reg [(3'h5):(1'h0)] reg3958 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3957 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3956 = (1'h0);
  reg [(4'hd):(1'h0)] reg3955 = (1'h0);
  reg [(5'h14):(1'h0)] reg3954 = (1'h0);
  reg [(2'h2):(1'h0)] reg3953 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3952 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3951 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3950 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3949 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3948 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3947 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3946 = (1'h0);
  reg [(4'hc):(1'h0)] reg3945 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3944 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3943 = (1'h0);
  reg [(5'h12):(1'h0)] reg3942 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3941 = (1'h0);
  reg [(3'h6):(1'h0)] reg3940 = (1'h0);
  reg [(4'h8):(1'h0)] reg3939 = (1'h0);
  reg [(5'h12):(1'h0)] reg3938 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3937 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3936 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3935 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3934 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3933 = (1'h0);
  reg [(5'h15):(1'h0)] reg3932 = (1'h0);
  reg [(4'hd):(1'h0)] reg3931 = (1'h0);
  reg [(4'hd):(1'h0)] reg3930 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar3929 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3928 = (1'h0);
  reg [(5'h19):(1'h0)] reg3927 = (1'h0);
  reg [(4'hd):(1'h0)] reg3926 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3925 = (1'h0);
  reg [(5'h17):(1'h0)] reg3924 = (1'h0);
  reg [(5'h16):(1'h0)] forvar3923 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3922 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3921 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3920 = (1'h0);
  reg [(4'hf):(1'h0)] reg3919 = (1'h0);
  reg [(5'h19):(1'h0)] forvar3918 = (1'h0);
  reg [(4'h9):(1'h0)] reg3917 = (1'h0);
  reg [(4'he):(1'h0)] reg3916 = (1'h0);
  reg [(5'h17):(1'h0)] reg3915 = (1'h0);
  reg [(3'h7):(1'h0)] reg3914 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3913 = (1'h0);
  reg [(5'h17):(1'h0)] reg3912 = (1'h0);
  reg [(4'hb):(1'h0)] reg3911 = (1'h0);
  reg [(5'h18):(1'h0)] reg3910 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3909 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3908 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3907 = (1'h0);
  reg [(3'h6):(1'h0)] reg3906 = (1'h0);
  reg [(2'h2):(1'h0)] reg3905 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3904 = (1'h0);
  reg [(4'hb):(1'h0)] reg3903 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3902 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3901 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3900 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3899 = (1'h0);
  reg [(5'h11):(1'h0)] forvar3898 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3897 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3896 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3895 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3894 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3893 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3892 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3891 = (1'h0);
  reg [(4'hb):(1'h0)] reg3890 = (1'h0);
  reg [(4'hb):(1'h0)] reg3889 = (1'h0);
  reg [(5'h16):(1'h0)] forvar3888 = (1'h0);
  reg [(5'h12):(1'h0)] reg3887 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3886 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3885 = (1'h0);
  reg [(4'hd):(1'h0)] reg3884 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3883 = (1'h0);
  reg [(4'h8):(1'h0)] reg3882 = (1'h0);
  reg [(2'h2):(1'h0)] reg3881 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3880 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3879 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3878 = (1'h0);
  reg [(4'ha):(1'h0)] reg3877 = (1'h0);
  reg [(5'h12):(1'h0)] reg3876 = (1'h0);
  reg [(5'h19):(1'h0)] reg3875 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3874 = (1'h0);
  reg [(5'h17):(1'h0)] reg3873 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3872 = (1'h0);
  reg [(2'h3):(1'h0)] reg3871 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3870 = (1'h0);
  reg [(5'h15):(1'h0)] reg3869 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3868 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3867 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar3866 = (1'h0);
  reg [(2'h3):(1'h0)] reg3865 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3864 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3863 = (1'h0);
  reg [(5'h19):(1'h0)] reg3862 = (1'h0);
  reg [(3'h7):(1'h0)] reg3861 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3860 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3859 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3858 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3857 = (1'h0);
  reg [(5'h14):(1'h0)] forvar3856 = (1'h0);
  wire [(5'h1a):(1'h0)] wire3855;
  reg [(4'h8):(1'h0)] reg3854 = (1'h0);
  reg [(5'h19):(1'h0)] reg3853 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3852 = (1'h0);
  wire [(4'he):(1'h0)] wire3851;
  reg signed [(4'h8):(1'h0)] reg3850 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3849 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3848 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3847 = (1'h0);
  reg [(5'h10):(1'h0)] reg3846 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3845 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3844 = (1'h0);
  reg [(4'hb):(1'h0)] reg3843 = (1'h0);
  reg [(4'h9):(1'h0)] reg3842 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3841 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3840 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3839 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3838 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3837 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3836 = (1'h0);
  reg [(2'h2):(1'h0)] reg3835 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3834 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3833 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3832 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3831 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3830 = (1'h0);
  reg [(2'h2):(1'h0)] reg3829 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3828 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire3827;
  reg signed [(2'h2):(1'h0)] reg3826 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3825 = (1'h0);
  reg [(5'h14):(1'h0)] reg3824 = (1'h0);
  reg [(5'h17):(1'h0)] reg3823 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3822 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3821 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3820 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3819 = (1'h0);
  reg [(5'h11):(1'h0)] reg3818 = (1'h0);
  reg [(5'h10):(1'h0)] reg3817 = (1'h0);
  reg [(5'h15):(1'h0)] reg3816 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3815 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3814 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3813 = (1'h0);
  reg [(3'h6):(1'h0)] reg3812 = (1'h0);
  reg [(2'h3):(1'h0)] reg3811 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar3810 = (1'h0);
  reg [(4'hd):(1'h0)] reg3809 = (1'h0);
  reg [(4'ha):(1'h0)] reg3808 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3807 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3806 = (1'h0);
  reg [(5'h13):(1'h0)] reg3805 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3804 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3803 = (1'h0);
  reg [(5'h16):(1'h0)] reg3802 = (1'h0);
  reg [(5'h16):(1'h0)] reg3801 = (1'h0);
  reg [(5'h12):(1'h0)] reg3800 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3799 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3798 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar3797 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar3796 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3795 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar3794 = (1'h0);
  reg [(3'h7):(1'h0)] reg3793 = (1'h0);
  reg [(4'hd):(1'h0)] reg3792 = (1'h0);
  reg [(4'hf):(1'h0)] reg3791 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3790 = (1'h0);
  reg [(5'h11):(1'h0)] forvar3789 = (1'h0);
  reg [(4'ha):(1'h0)] reg3788 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3787 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3786 = (1'h0);
  reg [(2'h3):(1'h0)] reg3785 = (1'h0);
  reg [(4'h8):(1'h0)] reg3784 = (1'h0);
  reg [(5'h11):(1'h0)] forvar3783 = (1'h0);
  reg [(4'hb):(1'h0)] reg3782 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3781 = (1'h0);
  reg [(2'h2):(1'h0)] reg3780 = (1'h0);
  reg [(5'h14):(1'h0)] reg3779 = (1'h0);
  reg [(2'h3):(1'h0)] reg3778 = (1'h0);
  reg [(4'hb):(1'h0)] reg3777 = (1'h0);
  reg [(5'h10):(1'h0)] reg3776 = (1'h0);
  reg [(4'he):(1'h0)] reg3775 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3774 = (1'h0);
  reg [(5'h13):(1'h0)] reg3773 = (1'h0);
  reg [(5'h18):(1'h0)] reg3772 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar3770 = (1'h0);
  reg [(2'h2):(1'h0)] reg3769 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3766 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar3764 = (1'h0);
  reg [(2'h3):(1'h0)] reg3763 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3762 = (1'h0);
  reg [(5'h16):(1'h0)] reg3771 = (1'h0);
  reg [(4'ha):(1'h0)] reg3770 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3769 = (1'h0);
  reg [(5'h15):(1'h0)] reg3768 = (1'h0);
  reg [(5'h12):(1'h0)] reg3767 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3766 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3765 = (1'h0);
  reg [(4'h8):(1'h0)] reg3764 = (1'h0);
  reg [(5'h15):(1'h0)] forvar3763 = (1'h0);
  reg [(4'he):(1'h0)] forvar3762 = (1'h0);
  reg [(5'h17):(1'h0)] reg3761 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3760 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3759 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3758 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3757 = (1'h0);
  reg [(4'hd):(1'h0)] reg3756 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3755 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3754 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar3753 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3752 = (1'h0);
  reg [(5'h15):(1'h0)] reg3751 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3750 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3749 = (1'h0);
  reg [(3'h7):(1'h0)] reg3748 = (1'h0);
  reg [(5'h18):(1'h0)] reg3747 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3746 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3745 = (1'h0);
  reg [(3'h4):(1'h0)] reg3744 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3743 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3742 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3741 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3740 = (1'h0);
  reg [(3'h6):(1'h0)] reg3739 = (1'h0);
  reg [(3'h4):(1'h0)] reg3738 = (1'h0);
  reg [(5'h12):(1'h0)] forvar3737 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar3736 = (1'h0);
  reg [(5'h17):(1'h0)] reg3735 = (1'h0);
  reg [(5'h10):(1'h0)] reg3734 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3733 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3732 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3730 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3728 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3731 = (1'h0);
  reg [(3'h6):(1'h0)] reg3730 = (1'h0);
  reg [(4'h9):(1'h0)] reg3729 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3728 = (1'h0);
  reg [(5'h14):(1'h0)] reg3727 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3726 = (1'h0);
  reg [(5'h18):(1'h0)] reg3725 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3724 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3723 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3722 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3721 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3720 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar3719 = (1'h0);
  reg [(5'h19):(1'h0)] reg3718 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3717 = (1'h0);
  reg [(5'h15):(1'h0)] reg3716 = (1'h0);
  reg [(4'hd):(1'h0)] reg3715 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3714 = (1'h0);
  reg [(4'h8):(1'h0)] reg3713 = (1'h0);
  wire signed [(5'h19):(1'h0)] wire3712;
  reg signed [(4'hc):(1'h0)] reg3711 = (1'h0);
  reg [(3'h5):(1'h0)] reg3710 = (1'h0);
  reg [(5'h15):(1'h0)] reg3709 = (1'h0);
  reg [(5'h10):(1'h0)] reg3708 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3707 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3706 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3705 = (1'h0);
  reg [(3'h5):(1'h0)] reg3704 = (1'h0);
  reg [(5'h14):(1'h0)] reg3703 = (1'h0);
  reg [(4'he):(1'h0)] reg3702 = (1'h0);
  assign y = {reg3974,
                 reg3973,
                 reg3972,
                 reg3971,
                 forvar3970,
                 reg3969,
                 forvar3968,
                 reg3967,
                 reg3966,
                 reg3965,
                 reg3964,
                 reg3963,
                 forvar3962,
                 reg3961,
                 forvar3960,
                 reg3959,
                 reg3958,
                 reg3957,
                 reg3956,
                 reg3955,
                 reg3954,
                 reg3953,
                 reg3952,
                 forvar3951,
                 reg3950,
                 reg3949,
                 reg3948,
                 reg3947,
                 reg3946,
                 reg3945,
                 forvar3944,
                 forvar3943,
                 reg3942,
                 forvar3941,
                 reg3940,
                 reg3939,
                 reg3938,
                 reg3937,
                 reg3936,
                 reg3935,
                 forvar3934,
                 reg3933,
                 reg3932,
                 reg3931,
                 reg3930,
                 forvar3929,
                 forvar3928,
                 reg3927,
                 reg3926,
                 forvar3925,
                 reg3924,
                 forvar3923,
                 reg3922,
                 forvar3921,
                 reg3920,
                 reg3919,
                 forvar3918,
                 reg3917,
                 reg3916,
                 reg3915,
                 reg3914,
                 forvar3913,
                 reg3912,
                 reg3911,
                 reg3910,
                 reg3909,
                 forvar3908,
                 reg3907,
                 reg3906,
                 reg3905,
                 reg3904,
                 reg3903,
                 reg3902,
                 reg3901,
                 forvar3900,
                 reg3899,
                 forvar3898,
                 reg3897,
                 reg3896,
                 reg3895,
                 reg3894,
                 reg3893,
                 forvar3892,
                 forvar3891,
                 reg3890,
                 reg3889,
                 forvar3888,
                 reg3887,
                 reg3886,
                 reg3885,
                 reg3884,
                 reg3883,
                 reg3882,
                 reg3881,
                 forvar3880,
                 reg3879,
                 reg3878,
                 reg3877,
                 reg3876,
                 reg3875,
                 reg3874,
                 reg3873,
                 forvar3872,
                 reg3871,
                 forvar3870,
                 reg3869,
                 reg3868,
                 reg3867,
                 forvar3866,
                 reg3865,
                 reg3864,
                 reg3863,
                 reg3862,
                 reg3861,
                 reg3860,
                 forvar3859,
                 reg3858,
                 reg3857,
                 forvar3856,
                 wire3855,
                 reg3854,
                 reg3853,
                 reg3852,
                 wire3851,
                 reg3850,
                 reg3849,
                 forvar3848,
                 reg3847,
                 reg3846,
                 reg3845,
                 forvar3844,
                 reg3843,
                 reg3842,
                 reg3841,
                 reg3840,
                 reg3839,
                 reg3838,
                 forvar3837,
                 reg3836,
                 reg3835,
                 reg3834,
                 reg3833,
                 reg3832,
                 forvar3831,
                 forvar3830,
                 reg3829,
                 reg3828,
                 wire3827,
                 reg3826,
                 reg3825,
                 reg3824,
                 reg3823,
                 reg3822,
                 forvar3821,
                 reg3820,
                 reg3819,
                 reg3818,
                 reg3817,
                 reg3816,
                 reg3815,
                 reg3814,
                 reg3813,
                 reg3812,
                 reg3811,
                 forvar3810,
                 reg3809,
                 reg3808,
                 reg3807,
                 reg3806,
                 reg3805,
                 forvar3804,
                 forvar3803,
                 reg3802,
                 reg3801,
                 reg3800,
                 reg3799,
                 reg3798,
                 forvar3797,
                 forvar3796,
                 reg3795,
                 forvar3794,
                 reg3793,
                 reg3792,
                 reg3791,
                 forvar3790,
                 forvar3789,
                 reg3788,
                 reg3787,
                 reg3786,
                 reg3785,
                 reg3784,
                 forvar3783,
                 reg3782,
                 forvar3781,
                 reg3780,
                 reg3779,
                 reg3778,
                 reg3777,
                 reg3776,
                 reg3775,
                 reg3774,
                 reg3773,
                 reg3772,
                 forvar3770,
                 reg3769,
                 forvar3766,
                 forvar3764,
                 reg3763,
                 reg3762,
                 reg3771,
                 reg3770,
                 forvar3769,
                 reg3768,
                 reg3767,
                 reg3766,
                 reg3765,
                 reg3764,
                 forvar3763,
                 forvar3762,
                 reg3761,
                 reg3760,
                 reg3759,
                 reg3758,
                 reg3757,
                 reg3756,
                 forvar3755,
                 reg3754,
                 forvar3753,
                 reg3752,
                 reg3751,
                 reg3750,
                 reg3749,
                 reg3748,
                 reg3747,
                 reg3746,
                 reg3745,
                 reg3744,
                 reg3743,
                 reg3742,
                 reg3741,
                 reg3740,
                 reg3739,
                 reg3738,
                 forvar3737,
                 forvar3736,
                 reg3735,
                 reg3734,
                 reg3733,
                 reg3732,
                 forvar3730,
                 reg3728,
                 reg3731,
                 reg3730,
                 reg3729,
                 forvar3728,
                 reg3727,
                 reg3726,
                 reg3725,
                 reg3724,
                 reg3723,
                 reg3722,
                 reg3721,
                 reg3720,
                 forvar3719,
                 reg3718,
                 reg3717,
                 reg3716,
                 reg3715,
                 forvar3714,
                 reg3713,
                 wire3712,
                 reg3711,
                 reg3710,
                 reg3709,
                 reg3708,
                 reg3707,
                 reg3706,
                 forvar3705,
                 reg3704,
                 reg3703,
                 reg3702,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg3702 = wire3699;
      reg3703 <= (^~(reg3702 ^~ $signed({(~&wire3699)})));
      reg3704 <= {wire3701};
    end
  always
    @(posedge clk) begin
      for (forvar3705 = (1'h0); (forvar3705 < (1'h1)); forvar3705 = (forvar3705 + (1'h1)))
        begin
          reg3706 <= reg3702;
          reg3707 <= $signed($unsigned(("NikA0msCVRC1CC3o" ?
              ("UAxcTMJ2MgWT37L2" << {reg3706}) : "WVaLrF0a7gDKA57SdO")));
          reg3708 <= reg3702[(2'h2):(1'h0)];
          reg3709 <= wire3701;
          reg3710 <= "DXTTYCaLDPNuaManWueNzX";
          reg3711 <= $unsigned(reg3707);
        end
    end
  assign wire3712 = $signed(wire3700);
  always
    @(posedge clk) begin
      reg3713 <= forvar3705;
      for (forvar3714 = (1'h0); (forvar3714 < (1'h1)); forvar3714 = (forvar3714 + (1'h1)))
        begin
          reg3715 = (wire3701[(1'h0):(1'h0)] ?
              $signed($signed(($unsigned((8'hae)) ?
                  ((7'h4b) <<< reg3706) : (reg3706 ?
                      reg3707 : wire3698)))) : (("gyBCmXYC1bIseQq" ?
                      ((-wire3697) ~^ (reg3706 ?
                          (8'hbe) : reg3709)) : "kXODuGBCIS") ?
                  (^~(wire3698 ?
                      wire3701 : (~|(7'h41)))) : $unsigned(($signed(reg3710) ?
                      (+wire3700) : "FGWW3z31FP4A4xVbt"))));
          reg3716 <= wire3697;
          reg3717 <= ((+((reg3715 ? $unsigned(wire3701) : $unsigned(reg3713)) ?
              (~^{reg3713}) : reg3709)) - {("d4THw" ?
                  (&$unsigned(forvar3705)) : ({wire3700,
                      reg3708} <= $signed(reg3703)))});
          reg3718 = reg3709;
          for (forvar3719 = (1'h0); (forvar3719 < (3'h4)); forvar3719 = (forvar3719 + (1'h1)))
            begin
              reg3720 <= $unsigned(($signed(({(8'ha4)} ?
                  reg3717 : reg3717[(2'h2):(2'h2)])) ^ $unsigned(forvar3705[(1'h1):(1'h1)])));
              reg3721 <= ("BxIO" > reg3702[(3'h4):(1'h1)]);
              reg3722 <= ($signed((^($signed(wire3701) >> "PS9ybpxPgyw4v22zDMoCnso7"))) ?
                  forvar3714 : ("cnzwmiKCoFDQ4cL9ZpTUBAlTF" + reg3720));
            end
          reg3723 <= ({(forvar3719 ?
                  reg3718 : reg3721[(4'hd):(4'h9)])} <= $signed($signed((~^wire3699))));
        end
      reg3724 = {reg3704};
      reg3725 <= (((8'ha7) ?
          $unsigned((reg3709 >= forvar3714)) : (7'h49)) ~^ $unsigned((~$unsigned($unsigned(reg3711)))));
      reg3726 <= "wnRb0Ixz";
    end
  always
    @(posedge clk) begin
      reg3727 <= $unsigned(reg3725);
      if (wire3698)
        begin
          for (forvar3728 = (1'h0); (forvar3728 < (3'h5)); forvar3728 = (forvar3728 + (1'h1)))
            begin
              reg3729 <= $signed(((!($unsigned(reg3721) ?
                      (~reg3709) : reg3715)) ?
                  $signed($unsigned({forvar3728, reg3720})) : (wire3699 ?
                      "xkGQ267yS6TmXKiAC73WDkdYn" : reg3717[(3'h5):(1'h1)])));
              reg3730 <= {{$unsigned($unsigned(((8'hb1) < (8'hbb)))),
                      ($unsigned((reg3726 ? (7'h4e) : reg3729)) ?
                          (reg3703 ?
                              (forvar3705 > wire3712) : (reg3726 ?
                                  reg3708 : reg3706)) : {wire3701[(1'h1):(1'h1)],
                              (reg3713 ^ wire3698)})}};
            end
          reg3731 = ((8'ha5) ?
              reg3711 : {({$unsigned(reg3706), $signed(wire3701)} ?
                      {reg3711, $unsigned(reg3713)} : "F45JpH4dste")});
        end
      else
        begin
          if (reg3708[(2'h3):(2'h3)])
            begin
              reg3728 <= (^~(~"BOewT0"));
              reg3729 = $signed((^~reg3709[(4'hf):(2'h2)]));
              for (forvar3730 = (1'h0); (forvar3730 < (1'h1)); forvar3730 = (forvar3730 + (1'h1)))
                begin
                  reg3731 <= wire3701[(1'h0):(1'h0)];
                  reg3732 <= ((+reg3716) == reg3730);
                  reg3733 <= (-(~|$signed(wire3698[(4'h8):(2'h2)])));
                end
              reg3734 <= reg3718;
            end
          else
            begin
              reg3728 <= "QhdhzXPTN1qN";
              reg3729 <= reg3728;
              for (forvar3730 = (1'h0); (forvar3730 < (1'h0)); forvar3730 = (forvar3730 + (1'h1)))
                begin
                  reg3731 = $signed($unsigned((^~(-(wire3698 ~^ (8'h9e))))));
                  reg3732 = reg3724;
                  reg3733 <= reg3722[(3'h4):(2'h3)];
                  reg3734 <= (((7'h44) ?
                      reg3709 : (8'h9c)) & $signed(("pqS" | ((8'haa) > forvar3719))));
                end
            end
          reg3735 <= "9kqRoa3HGum";
          for (forvar3736 = (1'h0); (forvar3736 < (3'h4)); forvar3736 = (forvar3736 + (1'h1)))
            begin
              for (forvar3737 = (1'h0); (forvar3737 < (3'h4)); forvar3737 = (forvar3737 + (1'h1)))
                begin
                  reg3738 <= (~reg3721[(4'h9):(2'h2)]);
                  reg3739 = (!($unsigned({$unsigned(reg3722)}) ?
                      ($unsigned($unsigned(wire3699)) + wire3712) : reg3722));
                  reg3740 <= reg3738;
                  reg3741 = "CyDVfbx";
                  reg3742 <= $signed($unsigned((reg3702[(2'h2):(1'h1)] ?
                      ((~reg3730) | $signed(forvar3728)) : $signed($signed(reg3709)))));
                  reg3743 <= {reg3703[(4'h8):(3'h4)]};
                end
              reg3744 = "4Jki0XxpLwWz5S0";
              reg3745 <= reg3742;
              reg3746 = $signed(reg3728[(3'h4):(2'h3)]);
            end
          reg3747 <= $signed(reg3721[(5'h15):(5'h11)]);
          reg3748 = reg3738;
        end
      reg3749 = ($unsigned(wire3701[(2'h3):(1'h0)]) != reg3720[(3'h4):(2'h2)]);
      if ((~$signed("VyuxW5QJLEKOvF4WiYTsR5t")))
        begin
          reg3750 <= ($signed((reg3710 ?
              $unsigned((reg3748 >> forvar3737)) : (!(forvar3705 >> reg3724)))) != (~|(8'ha8)));
        end
      else
        begin
          reg3750 <= reg3745[(4'h8):(3'h7)];
          reg3751 = (({(~&"8FIkegBRwlVmBTK7PpIrXo1")} - reg3721) << "eiiJ");
          reg3752 = reg3724[(4'h9):(4'h9)];
          for (forvar3753 = (1'h0); (forvar3753 < (1'h0)); forvar3753 = (forvar3753 + (1'h1)))
            begin
              reg3754 = $signed({wire3699, $signed((^~((8'hbc) ^ reg3713)))});
              for (forvar3755 = (1'h0); (forvar3755 < (1'h0)); forvar3755 = (forvar3755 + (1'h1)))
                begin
                  reg3756 <= $unsigned((reg3752[(1'h0):(1'h0)] ?
                      (~|reg3724) : {reg3721}));
                  reg3757 = wire3712[(5'h12):(4'ha)];
                  reg3758 <= (+($signed((reg3740 ?
                          reg3725[(4'h9):(3'h7)] : (-reg3734))) ?
                      (~"dSOMe9lVCYd9r1") : $signed($unsigned("9Ahf01sMHXqz0l"))));
                end
            end
          reg3759 = {$signed(((reg3729 < $unsigned(reg3746)) ?
                  $unsigned(reg3711[(4'hb):(4'ha)]) : $signed((forvar3753 ?
                      (8'haa) : reg3745))))};
          reg3760 <= (forvar3730[(3'h7):(2'h3)] < (($signed(reg3739[(1'h1):(1'h0)]) ?
                  (reg3752 ?
                      $signed(forvar3714) : "oeqfndKhQwIg7LU016m") : forvar3719[(1'h0):(1'h0)]) ?
              $unsigned({$unsigned(reg3742), reg3728}) : "wUDUCHF8Fu4wiCZ60"));
        end
      if ($signed((!"TL6QOUXT4")))
        begin
          reg3761 <= (wire3697 ?
              ((^$signed(reg3708)) + "loLQw02LfsN4LIKH5qbwQht") : $unsigned(reg3747));
          for (forvar3762 = (1'h0); (forvar3762 < (2'h3)); forvar3762 = (forvar3762 + (1'h1)))
            begin
              for (forvar3763 = (1'h0); (forvar3763 < (1'h0)); forvar3763 = (forvar3763 + (1'h1)))
                begin
                  reg3764 <= "II";
                  reg3765 = $unsigned((reg3722[(3'h6):(3'h4)] ?
                      ((|reg3723) & {(-forvar3762)}) : reg3703));
                  reg3766 = reg3704;
                end
            end
          reg3767 = (reg3722 ? "5g" : wire3699[(1'h1):(1'h1)]);
          reg3768 <= (+(forvar3728 > "VdgpPB1aSL1lZ"));
          for (forvar3769 = (1'h0); (forvar3769 < (2'h3)); forvar3769 = (forvar3769 + (1'h1)))
            begin
              reg3770 = $signed($unsigned(wire3699[(3'h7):(2'h2)]));
              reg3771 <= {$signed((~^$unsigned(wire3698))), $signed(reg3733)};
            end
        end
      else
        begin
          reg3761 = $unsigned({$unsigned((~^(~&(8'h9f)))),
              (($unsigned(forvar3769) ?
                  $signed(reg3741) : "I4tmBvDoPpHQL") <<< $unsigned("r1kcwJU41"))});
          reg3762 <= ((8'ha3) ?
              (~|reg3727) : ($signed(($unsigned(reg3728) <= {wire3698,
                  reg3713})) >>> reg3768));
          reg3763 <= (reg3746 ? $signed($unsigned(reg3760)) : reg3724);
          for (forvar3764 = (1'h0); (forvar3764 < (3'h4)); forvar3764 = (forvar3764 + (1'h1)))
            begin
              reg3765 = (reg3717[(3'h5):(3'h4)] >>> (^~reg3754[(1'h1):(1'h1)]));
              for (forvar3766 = (1'h0); (forvar3766 < (2'h2)); forvar3766 = (forvar3766 + (1'h1)))
                begin
                  reg3767 <= reg3747[(4'he):(1'h0)];
                  reg3768 <= reg3735[(5'h10):(3'h4)];
                  reg3769 <= (("ebclIAiX2f4IX5Z0sv8bc0K" ?
                          forvar3714[(1'h1):(1'h0)] : {forvar3736[(1'h1):(1'h1)],
                              (!reg3756)}) ?
                      ((&$signed($signed(reg3754))) ?
                          reg3743[(4'h8):(3'h6)] : forvar3737[(4'hd):(4'hd)]) : $unsigned($unsigned(reg3759)));
                end
              for (forvar3770 = (1'h0); (forvar3770 < (2'h3)); forvar3770 = (forvar3770 + (1'h1)))
                begin
                  reg3771 <= reg3762;
                  reg3772 <= $signed($unsigned(($unsigned("qIWwiDGU09hrlzLMda") ?
                      ((^wire3697) ?
                          $unsigned(reg3757) : $signed(reg3704)) : (8'ha0))));
                  reg3773 <= $signed($signed((($signed(reg3772) - reg3762[(3'h4):(1'h0)]) && (reg3731[(4'h9):(3'h6)] ?
                      (reg3750 ? (8'hac) : forvar3719) : (!forvar3737)))));
                  reg3774 = reg3748;
                  reg3775 <= (-("IKMl" - "TH9vCYtiTofS45a"));
                  reg3776 <= (^reg3722[(5'h12):(4'hd)]);
                end
            end
          reg3777 <= (("" ?
              (reg3750[(4'ha):(3'h7)] ?
                  $signed(((7'h42) ?
                      reg3750 : (7'h40))) : "b99JPrkRtehyW1caaHvNBNe") : "ppIbHAy8oyDZi4YTBFAWxF") ~^ reg3724);
          reg3778 <= $signed((&{(wire3700 >>> ((8'hb1) > reg3715))}));
        end
      reg3779 <= reg3769[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg3780 <= $unsigned((^~reg3710));
      for (forvar3781 = (1'h0); (forvar3781 < (1'h0)); forvar3781 = (forvar3781 + (1'h1)))
        begin
          reg3782 <= reg3757[(2'h3):(1'h1)];
          for (forvar3783 = (1'h0); (forvar3783 < (3'h5)); forvar3783 = (forvar3783 + (1'h1)))
            begin
              reg3784 <= (|reg3762);
              reg3785 <= (+$unsigned(reg3758[(1'h0):(1'h0)]));
              reg3786 <= ("Dnpl4KwO2xfmnoub9I1M3FMU3" >= ((reg3739[(1'h0):(1'h0)] ?
                      ((!(8'h9c)) ?
                          $unsigned(reg3740) : reg3728) : "FnoKmKRz63bVeupXkpY") ?
                  wire3697[(1'h0):(1'h0)] : reg3751));
            end
          reg3787 <= (^~$unsigned(((^(~reg3727)) ?
              (^~"XqN9645LuXq74") : reg3724)));
          reg3788 = "605qZkrtbWv9ZAq";
        end
      for (forvar3789 = (1'h0); (forvar3789 < (2'h2)); forvar3789 = (forvar3789 + (1'h1)))
        begin
          for (forvar3790 = (1'h0); (forvar3790 < (3'h4)); forvar3790 = (forvar3790 + (1'h1)))
            begin
              reg3791 <= (^(($signed((reg3739 & reg3784)) ?
                      reg3746[(2'h3):(1'h1)] : (reg3706[(5'h13):(1'h0)] || $signed(reg3735))) ?
                  ((~&wire3700) << forvar3770[(1'h1):(1'h1)]) : $signed((~&{reg3788}))));
              reg3792 = (8'haf);
              reg3793 <= (((^(forvar3789 >> "rvVTEBfBF9uGt7cmb")) ?
                  (+{forvar3755}) : ($signed(reg3738[(3'h4):(3'h4)]) ?
                      (forvar3781[(2'h3):(1'h0)] ?
                          (reg3760 + reg3734) : $signed(reg3788)) : "vX07x16FRQqI9122ZNJYtAPK")) & $unsigned(("8DDwtBHIzePwNBUlQcFQ" ?
                  forvar3764[(1'h0):(1'h0)] : forvar3755)));
              for (forvar3794 = (1'h0); (forvar3794 < (1'h1)); forvar3794 = (forvar3794 + (1'h1)))
                begin
                  reg3795 <= (reg3750[(5'h16):(4'ha)] ?
                      $unsigned((reg3752[(1'h0):(1'h0)] ?
                          (reg3702[(3'h7):(1'h1)] >>> (reg3754 & reg3758)) : $signed($signed((8'hac))))) : reg3757);
                end
            end
          for (forvar3796 = (1'h0); (forvar3796 < (1'h0)); forvar3796 = (forvar3796 + (1'h1)))
            begin
              for (forvar3797 = (1'h0); (forvar3797 < (3'h4)); forvar3797 = (forvar3797 + (1'h1)))
                begin
                  reg3798 <= "FildSERr0A";
                  reg3799 <= ("5ZKJgV8OInNC4BI0ci5QsXzz" >>> (($signed((reg3717 ?
                          (8'hae) : reg3730)) <<< reg3786) ?
                      "6SeN" : {(forvar3766 < $signed((8'hb2))),
                          $signed($signed(reg3716))}));
                end
              reg3800 = {$signed(((^~(~reg3720)) < $signed("TawipfhK2XaEJmwCf79WudmYp"))),
                  (^~$signed(((-reg3792) * (forvar3730 * reg3768))))};
              reg3801 <= reg3706;
              reg3802 <= reg3740;
            end
          for (forvar3803 = (1'h0); (forvar3803 < (1'h0)); forvar3803 = (forvar3803 + (1'h1)))
            begin
              for (forvar3804 = (1'h0); (forvar3804 < (1'h0)); forvar3804 = (forvar3804 + (1'h1)))
                begin
                  reg3805 = (~^"5YsJcqeReY8LCTMKDJht");
                  reg3806 <= (-"UI9Lt4q8AIbRGPZ");
                  reg3807 <= "ZkovMsUWrFpMdPA6";
                  reg3808 = {(reg3723 ? (!"i3bF") : "u8c9SPwlq1")};
                  reg3809 <= (~|(+(&$unsigned($unsigned((8'hb9))))));
                end
            end
          for (forvar3810 = (1'h0); (forvar3810 < (3'h5)); forvar3810 = (forvar3810 + (1'h1)))
            begin
              reg3811 <= ($signed($signed((((7'h4a) > reg3762) ?
                  reg3801[(4'ha):(4'h9)] : "nZkg1R"))) >> ($signed(((reg3757 | reg3785) - (reg3809 & (8'hb6)))) ?
                  $unsigned($unsigned(((8'h9f) ?
                      reg3788 : reg3766))) : "KogmAZPx5SPOIBLsGC6BAP"));
              reg3812 <= $signed($signed($unsigned(forvar3794[(3'h6):(2'h3)])));
              reg3813 <= $unsigned((($signed(reg3746[(2'h2):(1'h1)]) ?
                      reg3749 : (|(reg3743 ? reg3746 : forvar3764))) ?
                  $signed("ORh4ihr") : (&$unsigned(wire3701))));
              reg3814 <= (8'h9c);
              reg3815 = $signed((8'hb4));
            end
          reg3816 <= (reg3802 ? reg3706[(3'h7):(3'h5)] : "p");
          reg3817 <= "3bTbAkKtXflh90MrM4h4";
        end
      reg3818 <= {("ZArIxPKIWlrEGZzV" ?
              $unsigned($unsigned((^~reg3793))) : {$signed("bcNbFPxU2")})};
    end
  always
    @(posedge clk) begin
      reg3819 = reg3813;
      reg3820 = $signed(forvar3796);
      for (forvar3821 = (1'h0); (forvar3821 < (1'h0)); forvar3821 = (forvar3821 + (1'h1)))
        begin
          reg3822 <= ((~&$signed(("03BvxCIy" ?
              forvar3796 : $unsigned(reg3771)))) >>> $unsigned(reg3754[(1'h0):(1'h0)]));
          reg3823 = {reg3812[(1'h1):(1'h1)],
              (^~$unsigned((((8'ha3) && wire3712) ?
                  ((8'hb0) == wire3700) : $signed(reg3711))))};
          reg3824 <= ((!(-(-(&(7'h4a))))) << "WMQH7SSOrwYpZhJQDIyCiW9Sy");
          reg3825 <= $unsigned(forvar3755);
        end
      reg3826 <= $signed((($signed({reg3799}) ? (!"JLGkHyN6BD") : "eg4") ?
          (("ozYacBenOUqvi0XbDnPncrdo" ? (!(8'ha7)) : $signed(reg3763)) ?
              $signed($unsigned(reg3809)) : reg3795[(4'h8):(3'h7)]) : forvar3790[(1'h1):(1'h0)]));
    end
  assign wire3827 = reg3776[(4'h9):(3'h6)];
  always
    @(posedge clk) begin
      reg3828 <= $signed($unsigned(((+reg3763[(2'h3):(1'h0)]) == (reg3715 ?
          (reg3763 ? forvar3728 : (7'h41)) : (forvar3796 != reg3704)))));
      reg3829 <= forvar3719;
      for (forvar3830 = (1'h0); (forvar3830 < (3'h4)); forvar3830 = (forvar3830 + (1'h1)))
        begin
          for (forvar3831 = (1'h0); (forvar3831 < (2'h3)); forvar3831 = (forvar3831 + (1'h1)))
            begin
              reg3832 <= reg3772[(4'hd):(3'h7)];
              reg3833 <= $signed(($unsigned($unsigned($signed(forvar3804))) ?
                  ("YgCeiAk" ^~ reg3822[(5'h11):(5'h10)]) : $unsigned(reg3805[(2'h2):(1'h1)])));
              reg3834 <= {($signed($signed("b1f7q9scuOtuLmOHy7xA")) <<< $unsigned(reg3800[(3'h6):(1'h0)])),
                  (8'hbe)};
              reg3835 = ($signed($signed($unsigned((8'hbc)))) ?
                  {reg3703} : (~^forvar3719));
              reg3836 <= (reg3800[(4'hb):(3'h6)] ?
                  reg3758 : (((-reg3732[(4'ha):(2'h3)]) < "i0csEmeoFxWm") ^ {reg3727[(4'h9):(3'h7)]}));
              for (forvar3837 = (1'h0); (forvar3837 < (2'h3)); forvar3837 = (forvar3837 + (1'h1)))
                begin
                  reg3838 <= $signed((reg3767[(4'ha):(2'h3)] - ({(reg3728 ?
                              reg3759 : reg3792),
                          "vL2SicdOld0mwAJoE"} ?
                      $unsigned((reg3823 >>> reg3782)) : ($signed(forvar3790) | $unsigned(reg3754)))));
                  reg3839 <= $signed($signed((7'h40)));
                  reg3840 = (~reg3780[(1'h0):(1'h0)]);
                  reg3841 <= (~&reg3713);
                  reg3842 <= {("hXFGUS9SO3BMEyOCm2O" ^~ $unsigned(($unsigned(reg3720) * (&forvar3755))))};
                end
            end
          reg3843 <= $signed(reg3788[(4'h8):(3'h4)]);
        end
      for (forvar3844 = (1'h0); (forvar3844 < (3'h4)); forvar3844 = (forvar3844 + (1'h1)))
        begin
          reg3845 <= ($unsigned(forvar3810) ? forvar3728 : $unsigned(reg3725));
          reg3846 <= (!reg3809[(4'hc):(4'h9)]);
          reg3847 <= $signed(($unsigned(reg3778) ^~ reg3824));
        end
      for (forvar3848 = (1'h0); (forvar3848 < (2'h3)); forvar3848 = (forvar3848 + (1'h1)))
        begin
          reg3849 <= {"XqLULG05dug6EyWT4E15R", "UJeJHbNFZpdJ7HJcWVGcvBI"};
        end
      reg3850 <= ($signed("F") == "yE1ZdXeWcEl53LoxLp");
    end
  assign wire3851 = ("Zm0dIPGQpZxROs" ? "Hg" : reg3726[(5'h18):(5'h16)]);
  always
    @(posedge clk) begin
      reg3852 <= $signed({$signed("4trGI7GGF6YsU4ib6GYM4Y8k")});
      reg3853 <= {({reg3768} >> (($unsigned(reg3809) ?
                  (reg3817 ? reg3809 : reg3852) : "YSHun2n1AOiElRTmhcqGsyg") ?
              reg3704 : $signed("Wdfw")))};
      reg3854 <= reg3749;
    end
  assign wire3855 = {"X5hbGAG8nPeOfOI",
                        ($unsigned(reg3788) ?
                            ("TyTqUQkPdopD4kDcOW7aD2" << ({reg3792,
                                reg3772} - (^~wire3699))) : reg3776)};
  always
    @(posedge clk) begin
      for (forvar3856 = (1'h0); (forvar3856 < (1'h0)); forvar3856 = (forvar3856 + (1'h1)))
        begin
          reg3857 <= reg3717;
          reg3858 <= (8'hbf);
          for (forvar3859 = (1'h0); (forvar3859 < (1'h0)); forvar3859 = (forvar3859 + (1'h1)))
            begin
              reg3860 = ($unsigned((8'ha3)) + (^($signed(reg3710) >>> (^(reg3732 | reg3721)))));
              reg3861 <= reg3761;
              reg3862 = $unsigned(({($unsigned(reg3709) && $unsigned(forvar3728))} | $signed({(|wire3699),
                  (forvar3714 == reg3751)})));
              reg3863 <= forvar3794[(5'h1a):(3'h4)];
            end
          reg3864 <= reg3780;
        end
      reg3865 = "oDHy";
      for (forvar3866 = (1'h0); (forvar3866 < (1'h1)); forvar3866 = (forvar3866 + (1'h1)))
        begin
          reg3867 = "QuQciiCBJII1u";
          reg3868 = "EqPlt4HQ0ss0Cs";
          reg3869 <= reg3777[(4'h9):(1'h0)];
          for (forvar3870 = (1'h0); (forvar3870 < (1'h1)); forvar3870 = (forvar3870 + (1'h1)))
            begin
              reg3871 <= $unsigned((+"LNOAi"));
            end
          for (forvar3872 = (1'h0); (forvar3872 < (2'h2)); forvar3872 = (forvar3872 + (1'h1)))
            begin
              reg3873 <= $signed($unsigned(forvar3783[(2'h2):(1'h0)]));
              if (forvar3870[(2'h3):(2'h3)])
                begin
                  reg3874 = {"SX03MfD2gYiJU6kcpP2",
                      (reg3867 + $signed((reg3862 <<< "bLCdxg52g7S31F7m4NkE5")))};
                  reg3875 <= ("3YfgC9Xt7D" >> (reg3704[(3'h5):(1'h1)] >= $unsigned("AQf")));
                  reg3876 = $unsigned(reg3836[(3'h4):(2'h3)]);
                  reg3877 <= reg3812[(3'h5):(2'h3)];
                  reg3878 <= $unsigned((8'hbe));
                  reg3879 <= (reg3707[(4'hb):(3'h7)] || {($signed(reg3759[(1'h1):(1'h1)]) <= ((&reg3717) <<< $signed(reg3741))),
                      (8'ha4)});
                end
              else
                begin
                  reg3874 <= $unsigned((~^$signed($unsigned({reg3752,
                      forvar3730}))));
                  reg3875 <= ($unsigned(((~|$signed(forvar3764)) ?
                      $signed($unsigned(forvar3866)) : ($signed(reg3778) > reg3775))) <= reg3811[(2'h2):(2'h2)]);
                  reg3876 <= reg3734[(3'h6):(2'h2)];
                  reg3877 <= (~|$signed(forvar3796));
                end
              for (forvar3880 = (1'h0); (forvar3880 < (2'h2)); forvar3880 = (forvar3880 + (1'h1)))
                begin
                  reg3881 <= {reg3735};
                end
              reg3882 = {($signed($signed(wire3851[(1'h0):(1'h0)])) ?
                      ($unsigned(forvar3705) ?
                          (7'h46) : reg3759[(2'h2):(1'h1)]) : reg3707[(3'h5):(2'h2)]),
                  $unsigned($unsigned({(^reg3791)}))};
            end
        end
      reg3883 <= $signed(forvar3714[(2'h3):(2'h3)]);
      reg3884 = $unsigned($signed(reg3768[(3'h4):(2'h3)]));
      reg3885 <= reg3839[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg3886 <= $signed(((-reg3881) ?
          $signed(((~&forvar3790) + (reg3874 < reg3874))) : "HYzx4kxllL8JQelrQAs0AU"));
      reg3887 <= ("iMC1mrZa4V5pP0yR97Zxr" > $signed((((^reg3854) ?
          (^~reg3842) : $unsigned(reg3761)) ^ ("AVleAK58SZ4YObh4tXa2TJ8" <= (reg3802 ?
          reg3841 : reg3703)))));
      for (forvar3888 = (1'h0); (forvar3888 < (2'h3)); forvar3888 = (forvar3888 + (1'h1)))
        begin
          reg3889 <= "ht10TZ8BicrcEf0f";
          reg3890 <= $signed({(!$unsigned((7'h40)))});
          for (forvar3891 = (1'h0); (forvar3891 < (3'h5)); forvar3891 = (forvar3891 + (1'h1)))
            begin
              for (forvar3892 = (1'h0); (forvar3892 < (1'h0)); forvar3892 = (forvar3892 + (1'h1)))
                begin
                  reg3893 <= $unsigned(($signed((~^$unsigned((8'hb8)))) ?
                      (^reg3703) : reg3762[(4'ha):(4'ha)]));
                  reg3894 <= (("LMQXGLY4aFZ3cZ" ?
                      forvar3790[(4'h9):(3'h4)] : forvar3714[(2'h2):(1'h0)]) <<< (forvar3892 != ""));
                  reg3895 <= reg3865[(2'h3):(2'h3)];
                  reg3896 <= (~&(-($signed(reg3767[(3'h7):(1'h1)]) | (-(reg3748 < forvar3797)))));
                end
              reg3897 <= $unsigned($signed((~|"WsQGqT9xN9O0B")));
            end
          for (forvar3898 = (1'h0); (forvar3898 < (2'h2)); forvar3898 = (forvar3898 + (1'h1)))
            begin
              reg3899 <= reg3745[(3'h5):(2'h2)];
            end
          for (forvar3900 = (1'h0); (forvar3900 < (2'h2)); forvar3900 = (forvar3900 + (1'h1)))
            begin
              reg3901 <= $unsigned({"d",
                  (reg3702[(4'hb):(3'h5)] >>> "MbmZyxP")});
              reg3902 = (({reg3845} ?
                      $unsigned((forvar3844[(2'h3):(2'h2)] ?
                          $signed(reg3726) : $signed(reg3763))) : forvar3872[(2'h3):(1'h0)]) ?
                  ((~reg3775) ^ "B3Ox") : "EowIHFyyOiyw0Grk8Q45g");
              reg3903 <= "0vXD7dkrS09qn";
            end
          reg3904 <= reg3884[(3'h7):(3'h5)];
        end
      reg3905 <= ((reg3816[(5'h13):(1'h1)] ?
              {(reg3791 ? forvar3844 : $signed(reg3741)),
                  ("9YhEBCivwQxgI5ZwvoJ" ?
                      reg3813[(3'h5):(1'h1)] : $unsigned(reg3786))} : {(~forvar3880[(5'h10):(4'ha)]),
                  $signed("2sugEYzDuOvbfw4Awm2nmyu")}) ?
          (^~reg3853[(3'h7):(2'h2)]) : (8'hab));
    end
  always
    @(posedge clk) begin
      reg3906 <= $signed({reg3807, (7'h44)});
      reg3907 <= ((forvar3898 ?
              $unsigned(reg3768) : (^reg3838[(2'h2):(1'h1)])) ?
          (!(reg3758[(1'h1):(1'h0)] ?
              (reg3889[(1'h0):(1'h0)] < reg3730[(3'h6):(1'h1)]) : {reg3824,
                  (&reg3786)})) : $unsigned($unsigned(reg3879)));
      for (forvar3908 = (1'h0); (forvar3908 < (1'h0)); forvar3908 = (forvar3908 + (1'h1)))
        begin
          reg3909 = (~^$signed((~&reg3786[(2'h2):(1'h1)])));
          reg3910 <= ("uxkVuodN" <<< $signed("Hvl6RUIzM6Pdxz3RF"));
          reg3911 <= ($unsigned(({{forvar3821}, $unsigned(forvar3821)} ?
                  ($signed(reg3786) ?
                      $unsigned((8'hbb)) : "TASuXdr57JdknhwSL6L9kukT2") : $signed($signed(reg3795)))) ?
              reg3771 : reg3769[(1'h1):(1'h0)]);
          reg3912 <= $unsigned({reg3717});
          for (forvar3913 = (1'h0); (forvar3913 < (3'h4)); forvar3913 = (forvar3913 + (1'h1)))
            begin
              reg3914 <= reg3824;
            end
        end
    end
  always
    @(posedge clk) begin
      reg3915 <= (^~"T7tSPY0f");
      reg3916 = $signed(forvar3913[(4'hd):(4'h9)]);
    end
  always
    @(posedge clk) begin
      reg3917 <= ({$unsigned($unsigned($unsigned(reg3867)))} + reg3711);
      for (forvar3918 = (1'h0); (forvar3918 < (3'h4)); forvar3918 = (forvar3918 + (1'h1)))
        begin
          reg3919 <= reg3728;
          reg3920 <= (-"PPYii53NSrl1l2Gr71");
          for (forvar3921 = (1'h0); (forvar3921 < (3'h4)); forvar3921 = (forvar3921 + (1'h1)))
            begin
              reg3922 = (($signed("i") ?
                      $signed((reg3741 ?
                          (reg3799 ? reg3725 : forvar3762) : {reg3871,
                              (8'hb1)})) : (^~{"7KB3DK"})) ?
                  (8'hae) : $unsigned(((reg3784 - $unsigned(reg3776)) ?
                      ($signed(reg3890) ?
                          "h8LhsTTSIWNHV4LNRPG" : ((8'ha7) ?
                              reg3817 : (7'h4c))) : reg3873)));
              for (forvar3923 = (1'h0); (forvar3923 < (3'h5)); forvar3923 = (forvar3923 + (1'h1)))
                begin
                  reg3924 <= "tvH9RWJgADIwD7G5qp";
                end
            end
          for (forvar3925 = (1'h0); (forvar3925 < (1'h1)); forvar3925 = (forvar3925 + (1'h1)))
            begin
              reg3926 <= reg3896;
            end
          reg3927 <= ($signed((reg3834[(1'h1):(1'h1)] == ($signed(reg3850) + $unsigned(reg3791)))) ?
              $unsigned($unsigned("bHMlNlBhR")) : {$signed($signed(reg3907[(3'h7):(2'h2)])),
                  reg3912});
          for (forvar3928 = (1'h0); (forvar3928 < (2'h3)); forvar3928 = (forvar3928 + (1'h1)))
            begin
              for (forvar3929 = (1'h0); (forvar3929 < (2'h2)); forvar3929 = (forvar3929 + (1'h1)))
                begin
                  reg3930 = ($signed(("7RSo6wkzMHMW" < forvar3830[(2'h3):(1'h0)])) || ($signed(reg3717[(1'h1):(1'h1)]) ?
                      "iKOo4oJVW0H" : $signed(forvar3923)));
                  reg3931 <= "yly9Cn2w5xk";
                  reg3932 <= (forvar3783 ? reg3899 : reg3768[(3'h4):(3'h4)]);
                  reg3933 <= reg3858[(4'hd):(3'h6)];
                end
            end
        end
      for (forvar3934 = (1'h0); (forvar3934 < (2'h3)); forvar3934 = (forvar3934 + (1'h1)))
        begin
          reg3935 <= $signed(forvar3719);
          reg3936 <= $signed(((~^forvar3737) ?
              $unsigned(((forvar3764 ?
                  forvar3856 : reg3931) >> "oVSSxXkeotgsxTpHoYoCe")) : {(8'hbb)}));
          reg3937 <= $unsigned((~^$signed(reg3770)));
          reg3938 <= (~|forvar3848[(1'h1):(1'h0)]);
          reg3939 = $unsigned(reg3839[(3'h7):(3'h5)]);
        end
    end
  always
    @(posedge clk) begin
      reg3940 <= (((($unsigned((7'h4d)) != $signed((8'hb0))) ?
              reg3875 : $signed((7'h42))) >> $unsigned(("arsPcEqqCxaMOliSd" ?
              {reg3812} : ((7'h43) ? wire3698 : reg3798)))) ?
          $unsigned("sHYU9v7NqLHTVZOlna") : (~&(((forvar3797 ?
              reg3885 : (8'hbe)) ^ $signed(forvar3796)) ^~ "h2I4zrG123OHet7AwC")));
      for (forvar3941 = (1'h0); (forvar3941 < (3'h5)); forvar3941 = (forvar3941 + (1'h1)))
        begin
          reg3942 <= $signed((forvar3921[(3'h6):(1'h0)] << {$unsigned((^~reg3752))}));
          for (forvar3943 = (1'h0); (forvar3943 < (1'h1)); forvar3943 = (forvar3943 + (1'h1)))
            begin
              for (forvar3944 = (1'h0); (forvar3944 < (3'h4)); forvar3944 = (forvar3944 + (1'h1)))
                begin
                  reg3945 <= $signed("qLpRQoS1zccSPSgbhLMA");
                  reg3946 <= "l";
                  reg3947 <= (-("2NpvGWwWsJ4Tuw" & "7t"));
                  reg3948 <= reg3919;
                  reg3949 <= $signed({{$unsigned($unsigned(forvar3790))},
                      forvar3766[(3'h4):(2'h2)]});
                  reg3950 = (((!forvar3730[(4'hf):(4'h8)]) << $signed(($unsigned(reg3788) ?
                      $signed(reg3850) : (reg3948 >>> (8'h9e))))) ~^ $signed(forvar3929[(5'h15):(4'hb)]));
                end
              for (forvar3951 = (1'h0); (forvar3951 < (2'h2)); forvar3951 = (forvar3951 + (1'h1)))
                begin
                  reg3952 <= reg3879;
                  reg3953 = $signed(((!"0y3H06D3P1") ?
                      ((((8'hb5) >> forvar3925) ?
                              $signed(forvar3762) : reg3757) ?
                          $unsigned("3V1") : (^(^forvar3944))) : "tb2A"));
                  reg3954 = (reg3842[(1'h1):(1'h0)] * $unsigned($unsigned((reg3816 ?
                      $signed((8'hae)) : {reg3763}))));
                  reg3955 <= (|forvar3796[(4'hc):(3'h5)]);
                  reg3956 <= reg3733[(4'he):(4'hc)];
                end
            end
          reg3957 <= $signed({(~(-(reg3899 - reg3767)))});
          reg3958 <= "1Q0bn";
          reg3959 <= (reg3917[(1'h1):(1'h0)] ?
              $signed((reg3769 == forvar3900[(4'h9):(2'h3)])) : reg3955[(4'hd):(2'h2)]);
          for (forvar3960 = (1'h0); (forvar3960 < (3'h5)); forvar3960 = (forvar3960 + (1'h1)))
            begin
              reg3961 <= (reg3897 ? $signed("EmNDhiDKi") : reg3757);
              for (forvar3962 = (1'h0); (forvar3962 < (3'h4)); forvar3962 = (forvar3962 + (1'h1)))
                begin
                  reg3963 <= reg3858[(4'hd):(2'h2)];
                  reg3964 <= (8'hbd);
                  reg3965 = (|$unsigned(forvar3880[(4'hd):(4'hd)]));
                  reg3966 <= reg3835;
                end
              reg3967 <= (+(|"AX6"));
              for (forvar3968 = (1'h0); (forvar3968 < (2'h2)); forvar3968 = (forvar3968 + (1'h1)))
                begin
                  reg3969 <= "hq2S9mW5kxgIfNVSfM";
                end
              for (forvar3970 = (1'h0); (forvar3970 < (1'h0)); forvar3970 = (forvar3970 + (1'h1)))
                begin
                  reg3971 <= $unsigned((reg3730[(3'h6):(1'h1)] - $signed(reg3893)));
                  reg3972 = $signed(reg3839);
                  reg3973 <= "nQC8V";
                  reg3974 <= $unsigned(((forvar3888 ?
                      forvar3892 : (&(reg3708 - reg3752))) != (((+reg3852) == (~^reg3713)) + ((reg3713 ?
                          reg3740 : reg3716) ?
                      forvar3970[(4'hb):(4'h8)] : ""))));
                end
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3638
#( parameter param3692 = ({{(~|(|(8'hb8)))}, (&(((8'h9e) ? (8'hbc) : (7'h4b)) << ((8'hb2) << (7'h45))))} ? (-(^~(7'h40))) : {(((8'hb8) >> ((8'hb5) >= (7'h49))) ? (~&(^~(8'ha5))) : (8'hb5)), {(((8'hbd) * (7'h43)) <= (&(8'h9c))), (((8'hb3) < (8'ha0)) ? ((7'h48) + (8'hac)) : {(8'ha4), (8'hac)})}})
, parameter param3693 = ((((param3692 + (+param3692)) - (param3692 >>> param3692)) + param3692) ? ((~|(((8'hbb) ? param3692 : param3692) ? (7'h42) : (param3692 ^~ (7'h4d)))) ? ((-(param3692 <<< param3692)) ? param3692 : (7'h49)) : (^~{(param3692 ? param3692 : param3692), {param3692}})) : param3692) )
(y, clk, wire3643, wire3642, wire3641, wire3640, wire3639);
  output wire [(32'h279):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire3643;
  input wire [(4'ha):(1'h0)] wire3642;
  input wire signed [(5'h12):(1'h0)] wire3641;
  input wire [(4'hf):(1'h0)] wire3640;
  input wire signed [(2'h2):(1'h0)] wire3639;
  reg [(5'h19):(1'h0)] reg3691 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3690 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3689 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3688 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3687 = (1'h0);
  reg [(4'ha):(1'h0)] reg3686 = (1'h0);
  reg [(5'h15):(1'h0)] reg3685 = (1'h0);
  reg [(5'h17):(1'h0)] reg3684 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3683 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3682 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3681 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3680 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3679 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3678 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3677 = (1'h0);
  reg [(5'h17):(1'h0)] reg3676 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3675 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3674 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3673 = (1'h0);
  reg [(4'hf):(1'h0)] reg3672 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3671 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3670 = (1'h0);
  reg [(4'hc):(1'h0)] reg3669 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3668 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3667 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3666 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar3665 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3664 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3663 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3662 = (1'h0);
  reg [(3'h5):(1'h0)] reg3661 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3660 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3659 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3658 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar3657 = (1'h0);
  reg [(2'h3):(1'h0)] reg3656 = (1'h0);
  reg [(4'hf):(1'h0)] reg3655 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3654 = (1'h0);
  reg [(5'h15):(1'h0)] reg3653 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3652 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3651 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3650 = (1'h0);
  reg [(4'ha):(1'h0)] reg3649 = (1'h0);
  reg [(2'h3):(1'h0)] reg3648 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3647 = (1'h0);
  reg [(5'h17):(1'h0)] reg3646 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire3645;
  wire [(5'h10):(1'h0)] wire3644;
  assign y = {reg3691,
                 reg3690,
                 reg3689,
                 reg3688,
                 reg3687,
                 reg3686,
                 reg3685,
                 reg3684,
                 reg3683,
                 reg3682,
                 forvar3681,
                 reg3680,
                 reg3679,
                 forvar3678,
                 reg3677,
                 reg3676,
                 reg3675,
                 reg3674,
                 reg3673,
                 reg3672,
                 forvar3671,
                 forvar3670,
                 reg3669,
                 reg3668,
                 reg3667,
                 reg3666,
                 forvar3665,
                 reg3664,
                 reg3663,
                 reg3662,
                 reg3661,
                 reg3660,
                 reg3659,
                 reg3658,
                 forvar3657,
                 reg3656,
                 reg3655,
                 forvar3654,
                 reg3653,
                 forvar3652,
                 reg3651,
                 forvar3650,
                 reg3649,
                 reg3648,
                 reg3647,
                 reg3646,
                 wire3645,
                 wire3644,
                 (1'h0)};
  assign wire3644 = $unsigned(wire3642[(3'h7):(2'h3)]);
  assign wire3645 = $unsigned((-wire3642[(3'h4):(2'h2)]));
  always
    @(posedge clk) begin
      reg3646 = (wire3644 * (((~&((8'haf) - wire3644)) < $unsigned($signed(wire3644))) ?
          ($signed({(8'ha5), wire3645}) ?
              $signed(wire3641[(4'h8):(3'h7)]) : $signed(((7'h42) ?
                  wire3641 : wire3641))) : ($unsigned(wire3642) <<< $signed({wire3640,
              wire3639}))));
    end
  always
    @(posedge clk) begin
      reg3647 = {"qsKq13prBEYUoy8XLcHdP", wire3641[(2'h3):(2'h2)]};
      reg3648 <= $signed({wire3641[(4'ha):(2'h3)],
          {((~|wire3641) ?
                  "Uab5pnLrWfsYdw558" : (wire3641 ? (7'h42) : wire3641)),
              ((wire3641 * (8'hbe)) ? wire3641[(4'hd):(2'h2)] : "lc")}});
    end
  always
    @(posedge clk) begin
      reg3649 <= $signed((!$signed((8'h9f))));
    end
  always
    @(posedge clk) begin
      for (forvar3650 = (1'h0); (forvar3650 < (3'h4)); forvar3650 = (forvar3650 + (1'h1)))
        begin
          reg3651 <= "KdaXF8hmGxak4u56OJ";
          for (forvar3652 = (1'h0); (forvar3652 < (1'h0)); forvar3652 = (forvar3652 + (1'h1)))
            begin
              reg3653 = (^((~&"4J46AD5") ?
                  $signed((+reg3649)) : $signed((~$signed(wire3645)))));
              for (forvar3654 = (1'h0); (forvar3654 < (2'h2)); forvar3654 = (forvar3654 + (1'h1)))
                begin
                  reg3655 <= ($signed((((!wire3643) ?
                          (&(7'h42)) : $unsigned(wire3640)) * ((wire3641 >> reg3653) ?
                          "XxH9Bd8lK" : (wire3645 ? wire3641 : wire3639)))) ?
                      $signed(reg3647) : $signed(reg3649[(4'h8):(2'h2)]));
                  reg3656 = ({"pG30mto6OR4NthzNMh6Fy1g44",
                      ($signed(reg3646[(5'h13):(4'h9)]) ?
                          (+reg3651[(4'hd):(4'h8)]) : wire3645[(4'hb):(2'h3)])} * "NTWx");
                end
              for (forvar3657 = (1'h0); (forvar3657 < (3'h5)); forvar3657 = (forvar3657 + (1'h1)))
                begin
                  reg3658 = ("" ^ ($signed("R8TSEClHtDE83Xt8rBllAn8L") ?
                      forvar3654[(2'h3):(2'h2)] : reg3656[(1'h0):(1'h0)]));
                  reg3659 <= (reg3653 ? (~^reg3646) : reg3653);
                  reg3660 <= $unsigned("Mv3DS");
                  reg3661 <= "YNJdZSEJVRF0xme";
                  reg3662 = $unsigned("VuW6IwnduIyv");
                  reg3663 = ($signed("") && "yi3iBtUOrvmd42uYAICzmZtWZ");
                end
              reg3664 = forvar3652[(2'h2):(1'h0)];
              for (forvar3665 = (1'h0); (forvar3665 < (2'h3)); forvar3665 = (forvar3665 + (1'h1)))
                begin
                  reg3666 <= $unsigned(((($unsigned(wire3642) + (|forvar3665)) >= (~&$signed((7'h47)))) * ({$signed((8'hac))} ?
                      reg3647[(4'ha):(3'h7)] : (((7'h4d) ?
                          wire3641 : forvar3652) > {reg3646, reg3656}))));
                  reg3667 = {$unsigned((("PCz00LfU2Ig3rou221Hzq72" ?
                          {reg3664} : "d6kg") ~^ ({reg3662, (8'ha8)} ?
                          reg3666 : (reg3653 != forvar3654)))),
                      $unsigned($signed(($signed(wire3639) ?
                          reg3648[(1'h0):(1'h0)] : "hA9mGFn1SSDK1ABXd")))};
                  reg3668 <= reg3667;
                  reg3669 <= $unsigned(reg3653[(4'he):(4'ha)]);
                end
            end
          for (forvar3670 = (1'h0); (forvar3670 < (1'h1)); forvar3670 = (forvar3670 + (1'h1)))
            begin
              for (forvar3671 = (1'h0); (forvar3671 < (1'h1)); forvar3671 = (forvar3671 + (1'h1)))
                begin
                  reg3672 <= ("Z0vLbXht" ?
                      ("RnI5o5gRUR1" ?
                          $unsigned("GbCLKV5t49b0Z3TKyOJAfpCC") : (^~reg3661[(2'h3):(2'h3)])) : $unsigned("4k"));
                  reg3673 <= $signed(("h2y6e85N1H" <<< "DGwyZmXE"));
                  reg3674 <= (&$signed((($signed(reg3646) ^~ $signed((7'h42))) ?
                      (-(7'h45)) : "e7Mn06kJUryL0p6U")));
                  reg3675 <= reg3673;
                  reg3676 <= $unsigned($unsigned((!(~|forvar3671[(1'h0):(1'h0)]))));
                  reg3677 = (~&((~$signed((^reg3651))) ~^ ($signed((reg3668 ?
                      (8'hac) : reg3674)) << (~|$signed(reg3655)))));
                end
            end
          for (forvar3678 = (1'h0); (forvar3678 < (2'h3)); forvar3678 = (forvar3678 + (1'h1)))
            begin
              reg3679 <= "eSeU0";
              reg3680 = {(8'hab), wire3641[(3'h7):(2'h3)]};
              for (forvar3681 = (1'h0); (forvar3681 < (1'h0)); forvar3681 = (forvar3681 + (1'h1)))
                begin
                  reg3682 <= ((^~(reg3660 ?
                      "" : "y2KD1T94uc1kcixccCMuM")) != "wX7DbxMi");
                  reg3683 <= (^~forvar3665);
                  reg3684 <= (~(forvar3681[(3'h5):(2'h2)] <<< {("" || {forvar3671})}));
                end
            end
          reg3685 <= {"nMedNGlMFmG0US34XrBauDZl", "EuHy2GtKzmtgOaECzQDJhSk"};
          reg3686 = forvar3671;
        end
      reg3687 <= reg3663[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg3688 <= ({("hpzTvuYZQu6oyAvDpr" ?
                  (reg3669[(3'h7):(1'h1)] ?
                      reg3676 : $unsigned(reg3675)) : $unsigned("mdcTVAEwW"))} ?
          wire3643[(4'hb):(1'h0)] : (reg3653[(3'h4):(1'h1)] < ("aY57rnpfwqLY8zabKLxyX" ^ forvar3652[(1'h0):(1'h0)])));
      reg3689 <= (+(wire3645[(2'h3):(1'h1)] ?
          $unsigned("sJ1TPWBtSU") : (~&((~|reg3669) ?
              $signed((8'hbe)) : reg3674))));
      reg3690 = $unsigned("5RaecYPqBZ4UE");
      reg3691 <= (reg3667 >= wire3639[(1'h0):(1'h0)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3568
#( parameter param3635 = (!(((8'ha8) || ({(7'h4b), (7'h41)} ? ((7'h44) ? (8'hbd) : (8'h9c)) : ((7'h4c) ? (8'ha9) : (8'hb9)))) - (((!(7'h4d)) ? {(7'h42)} : ((8'ha3) > (8'haf))) ~^ (^((8'haf) | (7'h42)))))) )
(y, clk, wire3573, wire3572, wire3571, wire3570, wire3569);
  output wire [(32'h356):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire3573;
  input wire [(4'hc):(1'h0)] wire3572;
  input wire [(5'h14):(1'h0)] wire3571;
  input wire signed [(4'h8):(1'h0)] wire3570;
  input wire signed [(3'h4):(1'h0)] wire3569;
  reg signed [(4'h9):(1'h0)] reg3634 = (1'h0);
  reg [(4'hc):(1'h0)] reg3633 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3632 = (1'h0);
  reg [(5'h11):(1'h0)] reg3631 = (1'h0);
  reg [(5'h17):(1'h0)] reg3630 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3629 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire3628;
  reg signed [(5'h12):(1'h0)] reg3627 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3626 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3625 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire3624;
  reg [(5'h10):(1'h0)] reg3623 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3622 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire3621;
  wire [(4'h9):(1'h0)] wire3620;
  reg [(3'h6):(1'h0)] reg3619 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3618 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire3617;
  reg [(3'h4):(1'h0)] reg3616 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3615 = (1'h0);
  reg [(3'h4):(1'h0)] reg3614 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3613 = (1'h0);
  reg [(5'h19):(1'h0)] reg3612 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3611 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3610 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3609 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3608 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3607 = (1'h0);
  reg [(4'h9):(1'h0)] reg3606 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3605 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3604 = (1'h0);
  reg [(5'h12):(1'h0)] reg3603 = (1'h0);
  wire [(5'h11):(1'h0)] wire3602;
  reg [(4'h8):(1'h0)] reg3601 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3600 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3599 = (1'h0);
  reg [(4'h8):(1'h0)] reg3598 = (1'h0);
  reg [(5'h11):(1'h0)] reg3597 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3596 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3595 = (1'h0);
  reg [(5'h14):(1'h0)] forvar3594 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3593 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3592 = (1'h0);
  reg [(3'h4):(1'h0)] reg3591 = (1'h0);
  reg [(5'h19):(1'h0)] reg3590 = (1'h0);
  reg [(2'h3):(1'h0)] reg3589 = (1'h0);
  reg [(3'h5):(1'h0)] reg3588 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar3587 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3586 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3585 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3584 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3583 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3582 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3581 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3580 = (1'h0);
  reg [(4'hf):(1'h0)] reg3579 = (1'h0);
  reg [(5'h16):(1'h0)] reg3578 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3577 = (1'h0);
  reg [(2'h3):(1'h0)] reg3576 = (1'h0);
  wire [(2'h3):(1'h0)] wire3575;
  wire [(4'hd):(1'h0)] wire3574;
  assign y = {reg3634,
                 reg3633,
                 reg3632,
                 reg3631,
                 reg3630,
                 reg3629,
                 wire3628,
                 reg3627,
                 reg3626,
                 reg3625,
                 wire3624,
                 reg3623,
                 reg3622,
                 wire3621,
                 wire3620,
                 reg3619,
                 reg3618,
                 wire3617,
                 reg3616,
                 reg3615,
                 reg3614,
                 reg3613,
                 reg3612,
                 reg3611,
                 forvar3610,
                 reg3609,
                 reg3608,
                 reg3607,
                 reg3606,
                 reg3605,
                 reg3604,
                 reg3603,
                 wire3602,
                 reg3601,
                 reg3600,
                 forvar3599,
                 reg3598,
                 reg3597,
                 reg3596,
                 reg3595,
                 forvar3594,
                 reg3593,
                 reg3592,
                 reg3591,
                 reg3590,
                 reg3589,
                 reg3588,
                 forvar3587,
                 reg3586,
                 reg3585,
                 forvar3584,
                 reg3583,
                 reg3582,
                 forvar3581,
                 reg3580,
                 reg3579,
                 reg3578,
                 forvar3577,
                 reg3576,
                 wire3575,
                 wire3574,
                 (1'h0)};
  assign wire3574 = ("Y5hY1PEHqQiWOJiH" ?
                        (!$signed(wire3569)) : (~|$signed($unsigned(wire3571))));
  assign wire3575 = wire3569;
  always
    @(posedge clk) begin
      reg3576 = (8'hab);
      for (forvar3577 = (1'h0); (forvar3577 < (2'h2)); forvar3577 = (forvar3577 + (1'h1)))
        begin
          reg3578 <= {("3cg42K1QOFVW" < wire3570[(4'h8):(1'h0)]), wire3571};
          reg3579 <= reg3578;
        end
      reg3580 <= ($signed($signed(((~|wire3573) ?
              (~wire3572) : {(7'h4a), reg3576}))) ?
          ({$unsigned({wire3569})} != (+wire3574)) : ((wire3574 ?
              ($unsigned(reg3578) <= (reg3579 <= wire3573)) : ("nGRyCL1Ip" ?
                  $unsigned(wire3572) : (wire3572 || (8'hb9)))) | (^~(^$unsigned(forvar3577)))));
      for (forvar3581 = (1'h0); (forvar3581 < (2'h2)); forvar3581 = (forvar3581 + (1'h1)))
        begin
          reg3582 = $unsigned(wire3574);
          reg3583 <= $signed("uVCNfaneJ6GKc");
          for (forvar3584 = (1'h0); (forvar3584 < (3'h5)); forvar3584 = (forvar3584 + (1'h1)))
            begin
              reg3585 <= "6";
              reg3586 = ((($unsigned((wire3575 ?
                  (7'h42) : wire3569)) ^~ (&(+reg3579))) << forvar3584) > (^~"02mmnabsDkbCFR"));
              for (forvar3587 = (1'h0); (forvar3587 < (1'h0)); forvar3587 = (forvar3587 + (1'h1)))
                begin
                  reg3588 = $signed($signed(wire3571[(3'h7):(3'h5)]));
                  reg3589 <= wire3569[(2'h2):(2'h2)];
                  reg3590 <= $unsigned($signed((((wire3572 >= forvar3587) ?
                          (~&reg3580) : (forvar3581 ^ reg3589)) ?
                      "kt04SASpLdQ4HRy" : "HCr3zq8zXR5QqapD")));
                  reg3591 = "JFwQ";
                  reg3592 = {"s0q"};
                  reg3593 = "YThWHU";
                end
            end
          for (forvar3594 = (1'h0); (forvar3594 < (1'h0)); forvar3594 = (forvar3594 + (1'h1)))
            begin
              reg3595 <= (8'hb1);
              reg3596 <= reg3586[(3'h4):(2'h2)];
            end
          reg3597 <= $signed(((($unsigned(wire3572) >> (8'hbb)) ?
              $unsigned((forvar3587 ^~ forvar3581)) : "ZAnRlh2P4N8KdZo") < reg3578[(5'h15):(5'h13)]));
          reg3598 <= $unsigned(($signed(($signed(reg3591) ?
                  $unsigned(forvar3581) : reg3586)) ?
              ({reg3583, $unsigned(wire3572)} ?
                  reg3597[(3'h6):(1'h1)] : $signed($unsigned(reg3588))) : (~"1kTUMqsYpewERIJQTu")));
        end
      for (forvar3599 = (1'h0); (forvar3599 < (2'h2)); forvar3599 = (forvar3599 + (1'h1)))
        begin
          reg3600 = ($signed("YvmRfoMul5bPIs6dBwGDrK") & ($signed($signed(wire3569)) ?
              reg3592[(5'h11):(4'ha)] : {($unsigned(wire3572) || $signed(wire3569)),
                  {$unsigned((8'h9e)), $signed(wire3571)}}));
          reg3601 = (((^(|reg3576[(2'h3):(1'h0)])) - (8'ha5)) ?
              reg3596[(2'h2):(1'h1)] : wire3570);
        end
    end
  assign wire3602 = {$unsigned($signed(reg3588)),
                        ($signed(wire3572) ?
                            ($signed((reg3582 >> wire3569)) ?
                                ("NRDrmtIkFDiXfpmiQymVQ" >= $unsigned(wire3570)) : {$unsigned(wire3571)}) : $signed(wire3572))};
  always
    @(posedge clk) begin
      reg3603 = ((&(((forvar3587 ? reg3593 : forvar3577) ?
                  (reg3580 >> reg3591) : (wire3575 << wire3574)) ?
              $unsigned((reg3592 + forvar3587)) : "6ylS0bEr7NwBpEcZ452fMyMv")) ?
          ($signed({$unsigned(wire3574), $signed(reg3591)}) ?
              $signed($signed($unsigned(reg3601))) : (~"SlgACkN460Cwo")) : (($signed(wire3602) | (forvar3587 ?
                  wire3602 : (wire3570 ? reg3590 : (8'haa)))) ?
              $unsigned(({reg3601} ? {reg3596} : (~^(8'hb0)))) : wire3569));
      reg3604 <= (~&$unsigned("lDGv"));
      reg3605 <= reg3593[(4'he):(4'he)];
      reg3606 <= $unsigned($unsigned($signed((&"OTPqe"))));
      reg3607 <= (&$unsigned((^$unsigned((+reg3601)))));
    end
  always
    @(posedge clk) begin
      reg3608 <= reg3578[(3'h4):(3'h4)];
      if ($unsigned((~^{wire3573})))
        begin
          reg3609 <= ("zrdZXVFI0vpyGiGdnAOl" ?
              reg3595 : $unsigned($signed(reg3606)));
          for (forvar3610 = (1'h0); (forvar3610 < (3'h4)); forvar3610 = (forvar3610 + (1'h1)))
            begin
              reg3611 <= ("0SIKefbTO8O2v3wgKBN" ?
                  ((^~$signed((+wire3572))) ?
                      (^~"u3uxlPcYeWRa3XGoJkpy") : (wire3602 | (^$signed((8'h9d))))) : (wire3573 + forvar3587));
            end
          reg3612 = "4bqfOWV8outSDPd9raDf6";
        end
      else
        begin
          reg3609 <= reg3588;
        end
    end
  always
    @(posedge clk) begin
      reg3613 <= $unsigned((reg3590 + (forvar3594 + $signed($signed(wire3571)))));
      reg3614 <= reg3605;
      reg3615 <= forvar3599;
    end
  always
    @(posedge clk) begin
      reg3616 <= (wire3573 ^ reg3601);
    end
  assign wire3617 = ({$unsigned($signed("7kL2"))} ?
                        wire3569[(2'h2):(1'h0)] : $signed(reg3615[(5'h11):(3'h6)]));
  always
    @(posedge clk) begin
      reg3618 <= wire3569[(3'h4):(1'h0)];
      reg3619 <= ((~&$unsigned((-$unsigned(reg3616)))) ?
          (|($signed("") == reg3600[(3'h4):(1'h1)])) : {reg3593[(5'h15):(4'ha)]});
    end
  assign wire3620 = (7'h4a);
  assign wire3621 = (8'hae);
  always
    @(posedge clk) begin
      reg3622 <= ((({(^~reg3613)} >= wire3602) ?
          reg3576 : (wire3571 ?
              reg3600[(2'h3):(2'h2)] : reg3583[(4'he):(2'h3)])) | $unsigned($signed(((~|reg3591) == (reg3615 ?
          (8'hb1) : reg3611)))));
      reg3623 <= {(~&{((|wire3572) <<< (~^wire3570)), reg3586[(4'hd):(4'hc)]}),
          (reg3578 * "vvt2n6OkYzt0P")};
    end
  assign wire3624 = {$unsigned($signed($unsigned((wire3620 ?
                            reg3578 : reg3608))))};
  always
    @(posedge clk) begin
      reg3625 <= "WbUdbCyT3Uq0PZ";
      reg3626 <= ("Z7oU5Fq" ?
          ("GOzBOsIqZrdd02aWNi" >> $unsigned(((reg3585 | wire3602) ?
              "Gf1UOMoKxnFaT6ki" : {(7'h40), wire3621}))) : (^~(8'hb6)));
      reg3627 <= reg3591;
    end
  assign wire3628 = {$unsigned($signed(($signed((8'hb7)) ?
                            reg3588[(2'h3):(2'h2)] : {reg3616, reg3590})))};
  always
    @(posedge clk) begin
      reg3629 <= (forvar3577[(2'h3):(1'h1)] ?
          {"sLgDT08SHg", (8'had)} : reg3589);
      reg3630 <= $signed(reg3613);
      reg3631 <= $signed((~$unsigned($signed(reg3578))));
      reg3632 <= {(7'h49)};
      reg3633 <= "Lm0d7EQt3Ruo57kqCOVXcb";
      reg3634 <= (+wire3573[(3'h5):(3'h5)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3450
#( parameter param3565 = ((&{({(7'h45)} ? ((8'haa) ~^ (8'hac)) : (~(8'haa))), (((8'had) ^~ (7'h43)) >= (^(8'hab)))}) * (((^~((8'ha2) | (8'hb5))) | {((8'hb9) ? (8'hb4) : (8'hb5))}) << ({(~&(7'h4b))} >> ((&(8'ha1)) ? ((7'h44) ? (8'haa) : (7'h45)) : ((8'hb7) & (8'hb3)))))) )
(y, clk, wire3455, wire3454, wire3453, wire3452, wire3451);
  output wire [(32'h5e7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire3455;
  input wire [(5'h13):(1'h0)] wire3454;
  input wire [(4'hb):(1'h0)] wire3453;
  input wire signed [(3'h7):(1'h0)] wire3452;
  input wire signed [(3'h5):(1'h0)] wire3451;
  wire signed [(3'h4):(1'h0)] wire3564;
  reg [(3'h6):(1'h0)] reg3563 = (1'h0);
  reg [(5'h19):(1'h0)] forvar3562 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3561 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3560 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3559 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3558 = (1'h0);
  reg [(3'h4):(1'h0)] reg3557 = (1'h0);
  reg [(3'h4):(1'h0)] reg3556 = (1'h0);
  reg [(4'h8):(1'h0)] reg3555 = (1'h0);
  reg [(4'ha):(1'h0)] reg3554 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3553 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3552 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3551 = (1'h0);
  reg [(4'hf):(1'h0)] reg3550 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3549 = (1'h0);
  reg [(5'h15):(1'h0)] reg3548 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3547 = (1'h0);
  reg [(4'he):(1'h0)] forvar3546 = (1'h0);
  reg [(3'h6):(1'h0)] reg3545 = (1'h0);
  reg [(5'h18):(1'h0)] reg3544 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3543 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3542 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3541 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3540 = (1'h0);
  reg [(5'h10):(1'h0)] reg3539 = (1'h0);
  reg [(5'h11):(1'h0)] reg3538 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3537 = (1'h0);
  reg [(4'hc):(1'h0)] reg3536 = (1'h0);
  reg [(5'h18):(1'h0)] reg3535 = (1'h0);
  reg [(4'hb):(1'h0)] reg3534 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3533 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3532 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3531 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3530 = (1'h0);
  reg [(5'h10):(1'h0)] reg3529 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3528 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire3527;
  reg signed [(2'h2):(1'h0)] reg3526 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3525 = (1'h0);
  reg [(4'hf):(1'h0)] reg3524 = (1'h0);
  reg [(5'h10):(1'h0)] reg3523 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3522 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar3521 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3520 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3519 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3518 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3517 = (1'h0);
  reg [(5'h19):(1'h0)] reg3516 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3515 = (1'h0);
  reg [(5'h16):(1'h0)] reg3514 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3513 = (1'h0);
  reg [(4'ha):(1'h0)] reg3512 = (1'h0);
  reg [(4'ha):(1'h0)] reg3511 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3510 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3509 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3508 = (1'h0);
  reg [(5'h19):(1'h0)] reg3507 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3506 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3505 = (1'h0);
  reg [(3'h6):(1'h0)] reg3504 = (1'h0);
  reg [(3'h6):(1'h0)] reg3503 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3502 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar3501 = (1'h0);
  reg [(5'h15):(1'h0)] reg3500 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3499 = (1'h0);
  reg [(5'h16):(1'h0)] reg3498 = (1'h0);
  reg [(4'hf):(1'h0)] reg3497 = (1'h0);
  reg [(5'h14):(1'h0)] reg3496 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3495 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3494 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3493 = (1'h0);
  reg [(4'hb):(1'h0)] reg3492 = (1'h0);
  reg [(4'h8):(1'h0)] reg3491 = (1'h0);
  reg [(5'h14):(1'h0)] reg3490 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3489 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3488 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3487 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3486 = (1'h0);
  reg [(4'h8):(1'h0)] reg3485 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3484 = (1'h0);
  reg [(4'h9):(1'h0)] reg3483 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3482 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3481 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3480 = (1'h0);
  reg [(5'h15):(1'h0)] forvar3479 = (1'h0);
  reg [(4'h9):(1'h0)] reg3478 = (1'h0);
  reg [(4'hd):(1'h0)] reg3477 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3476 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3475 = (1'h0);
  reg [(4'he):(1'h0)] reg3474 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3473 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3472 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3471 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3470 = (1'h0);
  reg [(5'h12):(1'h0)] reg3469 = (1'h0);
  reg [(4'h8):(1'h0)] reg3468 = (1'h0);
  wire [(4'hf):(1'h0)] wire3467;
  reg [(3'h6):(1'h0)] reg3466 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3465 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3464 = (1'h0);
  reg [(4'hf):(1'h0)] reg3463 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3462 = (1'h0);
  reg [(5'h17):(1'h0)] reg3461 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire3460;
  reg [(2'h2):(1'h0)] reg3459 = (1'h0);
  reg [(5'h13):(1'h0)] reg3458 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3457 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3456 = (1'h0);
  assign y = {wire3564,
                 reg3563,
                 forvar3562,
                 reg3561,
                 reg3560,
                 reg3559,
                 forvar3558,
                 reg3557,
                 reg3556,
                 reg3555,
                 reg3554,
                 reg3553,
                 reg3552,
                 forvar3551,
                 reg3550,
                 reg3549,
                 reg3548,
                 reg3547,
                 forvar3546,
                 reg3545,
                 reg3544,
                 reg3543,
                 forvar3542,
                 reg3541,
                 reg3540,
                 reg3539,
                 reg3538,
                 forvar3537,
                 reg3536,
                 reg3535,
                 reg3534,
                 forvar3533,
                 reg3532,
                 reg3531,
                 reg3530,
                 reg3529,
                 forvar3528,
                 wire3527,
                 reg3526,
                 reg3525,
                 reg3524,
                 reg3523,
                 reg3522,
                 forvar3521,
                 reg3520,
                 reg3519,
                 reg3518,
                 reg3517,
                 reg3516,
                 reg3515,
                 reg3514,
                 forvar3513,
                 reg3512,
                 reg3511,
                 reg3510,
                 reg3509,
                 reg3508,
                 reg3507,
                 reg3506,
                 reg3505,
                 reg3504,
                 reg3503,
                 reg3502,
                 forvar3501,
                 reg3500,
                 forvar3499,
                 reg3498,
                 reg3497,
                 reg3496,
                 reg3495,
                 reg3494,
                 reg3493,
                 reg3492,
                 reg3491,
                 reg3490,
                 reg3489,
                 forvar3488,
                 forvar3487,
                 forvar3486,
                 reg3485,
                 reg3484,
                 reg3483,
                 reg3482,
                 reg3481,
                 reg3480,
                 forvar3479,
                 reg3478,
                 reg3477,
                 forvar3476,
                 reg3475,
                 reg3474,
                 reg3473,
                 reg3472,
                 reg3471,
                 forvar3470,
                 reg3469,
                 reg3468,
                 wire3467,
                 reg3466,
                 reg3465,
                 reg3464,
                 reg3463,
                 reg3462,
                 reg3461,
                 wire3460,
                 reg3459,
                 reg3458,
                 reg3457,
                 reg3456,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg3456 <= "PxgUQNegYKUMzCt5NR";
      reg3457 <= wire3451;
      reg3458 <= "7urr";
      reg3459 <= "PMYb1tZ6YNgp8iMT";
    end
  assign wire3460 = reg3456;
  always
    @(posedge clk) begin
      reg3461 <= {(^(&$unsigned("qtrpp7")))};
    end
  always
    @(posedge clk) begin
      reg3462 = $signed(reg3461[(5'h15):(5'h11)]);
      reg3463 <= wire3451;
    end
  always
    @(posedge clk) begin
      reg3464 <= $unsigned(("K1NwpSI5X88E" >> $unsigned(((wire3454 ?
          reg3456 : (8'hb8)) | wire3452))));
      reg3465 <= (-$signed((+(reg3461 ? wire3453 : "pFp0Ltvwt1"))));
      reg3466 <= reg3464;
    end
  assign wire3467 = $signed(reg3463);
  always
    @(posedge clk) begin
      reg3468 <= wire3452[(1'h1):(1'h0)];
      reg3469 <= $signed(reg3456[(2'h3):(1'h0)]);
    end
  always
    @(posedge clk) begin
      for (forvar3470 = (1'h0); (forvar3470 < (1'h1)); forvar3470 = (forvar3470 + (1'h1)))
        begin
          reg3471 <= "K7hbSNw4RRd4AS4rZY4popv";
          reg3472 <= "Gcma4pFTsFWLfBNO93A";
          reg3473 = $unsigned((!{"E4L7BeUGHlH0", ""}));
          reg3474 <= ("e6WcI" ?
              wire3451[(2'h3):(2'h2)] : ((7'h4e) ~^ wire3451[(2'h2):(1'h0)]));
        end
      reg3475 = (7'h4a);
      for (forvar3476 = (1'h0); (forvar3476 < (3'h5)); forvar3476 = (forvar3476 + (1'h1)))
        begin
          reg3477 = forvar3476;
          reg3478 <= (("6nwyBBWxNAzMo5za7n" && "r3RhwZnKXRHapOtZlS1") ?
              $signed(((~$unsigned(wire3467)) ?
                  reg3468 : $unsigned((reg3457 ?
                      reg3456 : reg3475)))) : $signed("cnbLObQeRxWvergMteN8f8"));
          for (forvar3479 = (1'h0); (forvar3479 < (2'h2)); forvar3479 = (forvar3479 + (1'h1)))
            begin
              reg3480 = ($signed("QZaFk7wmTVsoTBPOF1") <<< $signed((~^wire3452[(3'h6):(2'h3)])));
              reg3481 = ($signed({forvar3470}) >>> (wire3452 ?
                  "qODm2BbKz6ogp" : (-"")));
              reg3482 <= reg3469;
              reg3483 = ((~^reg3475) ? (~(8'had)) : reg3472[(2'h3):(2'h3)]);
            end
          reg3484 <= (((reg3481 <= ($signed(wire3451) << "mgXYLkA53tBg4KtxY4IM")) ?
                  ("ranaA" || "") : {(reg3459 >= (reg3456 - reg3471))}) ?
              reg3472 : ({((~|reg3475) | (reg3462 * reg3483))} <= $unsigned(((wire3467 ?
                      wire3467 : reg3465) ?
                  (reg3462 != wire3453) : $unsigned(forvar3479)))));
        end
      reg3485 <= {{$unsigned($signed((7'h44)))}};
      for (forvar3486 = (1'h0); (forvar3486 < (1'h1)); forvar3486 = (forvar3486 + (1'h1)))
        begin
          for (forvar3487 = (1'h0); (forvar3487 < (3'h4)); forvar3487 = (forvar3487 + (1'h1)))
            begin
              for (forvar3488 = (1'h0); (forvar3488 < (2'h2)); forvar3488 = (forvar3488 + (1'h1)))
                begin
                  reg3489 <= reg3469;
                  reg3490 = forvar3488;
                  reg3491 = wire3467[(2'h3):(2'h2)];
                end
              reg3492 <= "tPdDe9c";
              reg3493 = (~|(+(~&reg3461[(2'h3):(2'h3)])));
              reg3494 <= $unsigned($unsigned(reg3493[(2'h3):(1'h0)]));
            end
          reg3495 <= {((((reg3456 ? (8'hba) : reg3475) ?
                      {forvar3488} : (reg3489 ?
                          reg3484 : wire3455)) || "UoLg2XQMuslepmsQ") ?
                  ((~|wire3452[(3'h6):(2'h2)]) ?
                      "XBDEq" : ((7'h41) ?
                          "" : (forvar3486 ?
                              reg3471 : reg3494))) : $signed((((8'ha5) ?
                      reg3490 : wire3460) ^ $signed(reg3466))))};
          reg3496 <= (~$signed((forvar3486 ^ "9f9p")));
          reg3497 <= ((&(~|$signed("eggWMAQ"))) < $unsigned({($unsigned(reg3474) <<< $unsigned(reg3465)),
              "4VTn26t"}));
          reg3498 <= $signed((!"4gHq45TYbiUJ"));
        end
    end
  always
    @(posedge clk) begin
      for (forvar3499 = (1'h0); (forvar3499 < (2'h2)); forvar3499 = (forvar3499 + (1'h1)))
        begin
          reg3500 <= {$signed({$unsigned(reg3456[(2'h2):(2'h2)]),
                  {$unsigned((7'h47))}})};
          for (forvar3501 = (1'h0); (forvar3501 < (2'h2)); forvar3501 = (forvar3501 + (1'h1)))
            begin
              reg3502 <= (($signed(($unsigned(reg3498) ?
                      "UnYanMW8X" : (reg3459 ^~ (7'h4d)))) ?
                  "plQXQA" : $signed("cm")) ^ reg3498[(4'hf):(3'h4)]);
              if (((~|"K4h0m96DNXOtA6Tpiz0qrTTO") == $unsigned($unsigned((~^{reg3484,
                  reg3493})))))
                begin
                  reg3503 <= (reg3462 ?
                      ({forvar3476[(2'h2):(1'h1)],
                              $signed(reg3497[(3'h5):(1'h1)])} ?
                          (({reg3472} ?
                              $signed(reg3456) : "aTK") << reg3489[(4'hd):(4'hb)]) : "zP1oonJ3myecn3AveIWn") : "FgncWm");
                  reg3504 <= {($unsigned({$unsigned(reg3462),
                          $unsigned(reg3496)}) ^~ (reg3475[(5'h11):(4'h9)] ?
                          wire3452 : $signed(reg3466[(1'h0):(1'h0)]))),
                      $unsigned(reg3472)};
                  reg3505 = $signed("RPh5vYa0B0Sr4YU1");
                  reg3506 <= "cN3AG8hXNQKBF";
                  reg3507 <= (&$unsigned($unsigned($signed($signed(reg3457)))));
                  reg3508 <= reg3506[(1'h1):(1'h0)];
                end
              else
                begin
                  reg3503 <= reg3507[(5'h15):(5'h13)];
                  reg3504 <= reg3457[(3'h7):(3'h7)];
                  reg3505 <= {{reg3468}};
                  reg3506 = $signed("");
                  reg3507 <= reg3502[(3'h4):(1'h1)];
                end
            end
          reg3509 <= $signed(wire3451[(3'h5):(3'h5)]);
          reg3510 <= ("2V5Vd2bNWVnINepsE" ?
              reg3490 : $signed((~|(~&(!reg3474)))));
        end
      reg3511 <= "LgnQ";
      reg3512 = reg3500[(5'h15):(4'he)];
      for (forvar3513 = (1'h0); (forvar3513 < (3'h5)); forvar3513 = (forvar3513 + (1'h1)))
        begin
          reg3514 <= $signed("YEFdBi0FlqB");
          reg3515 = ($unsigned(((reg3511 ^~ (~&(7'h45))) < ("esJYyZV1NegpksVUfI" ?
                  "tIGFgztLuvwuc5CBqtL5sKlT2" : reg3481))) ?
              (&$signed({(reg3514 - (7'h4c))})) : reg3504[(2'h3):(1'h1)]);
          reg3516 <= (($unsigned((~|(reg3490 == reg3483))) ^ forvar3488) ?
              ($signed(((7'h47) - reg3506[(3'h4):(2'h2)])) > (!{reg3506[(5'h12):(4'hf)],
                  $unsigned(reg3505)})) : ((wire3454[(3'h5):(3'h4)] ?
                  reg3511 : (~&(8'hb6))) <= {$signed(forvar3486), reg3514}));
          reg3517 <= (&(reg3471 >>> (wire3467 ?
              $unsigned($signed(reg3505)) : "9Hs")));
          reg3518 <= (reg3508 ?
              (~^"HGgkIqscJgfbBGPr0G8ile78V") : (|$unsigned(reg3498[(4'h9):(4'h8)])));
        end
    end
  always
    @(posedge clk) begin
      reg3519 <= $unsigned(("k0iEVeDWERl41B" ?
          $unsigned(reg3461[(4'hd):(4'ha)]) : ("K" + $signed((8'had)))));
      reg3520 <= $unsigned((-(^~$unsigned($signed(reg3516)))));
      for (forvar3521 = (1'h0); (forvar3521 < (2'h3)); forvar3521 = (forvar3521 + (1'h1)))
        begin
          reg3522 <= $unsigned(forvar3499[(3'h4):(1'h1)]);
          reg3523 <= reg3468[(2'h3):(2'h3)];
          reg3524 <= (&({(+(reg3504 + reg3474))} ?
              {$unsigned($unsigned((7'h4d)))} : $unsigned($unsigned(reg3483[(1'h1):(1'h0)]))));
          reg3525 <= (~{forvar3476});
        end
      reg3526 = (8'hb8);
    end
  assign wire3527 = (($unsigned($signed({(7'h49)})) ?
                            $unsigned({""}) : {($signed((8'ha5)) * (forvar3479 <= wire3453))}) ?
                        {{forvar3521[(5'h12):(4'h9)],
                                (reg3519[(5'h10):(4'hc)] ?
                                    {reg3465} : "dQqA5mR1K6el")},
                            "cIahq3"} : $signed($unsigned(("khOHtLe" || "AKA6vssEwKJ5FSa"))));
  always
    @(posedge clk) begin
      for (forvar3528 = (1'h0); (forvar3528 < (2'h3)); forvar3528 = (forvar3528 + (1'h1)))
        begin
          reg3529 <= forvar3487[(3'h5):(2'h3)];
        end
      reg3530 <= (~^("4XOguzW1WuybK1Vkm6" ? reg3522 : "bPC0J0EHH5ug5ykbLApp"));
    end
  always
    @(posedge clk) begin
      reg3531 <= reg3474[(3'h6):(3'h4)];
      reg3532 <= "ex9VO2HOTbwCbQLD";
      for (forvar3533 = (1'h0); (forvar3533 < (3'h5)); forvar3533 = (forvar3533 + (1'h1)))
        begin
          reg3534 <= $signed((({(reg3502 ? reg3498 : reg3473),
                      $unsigned((7'h4e))} ?
                  reg3480[(1'h0):(1'h0)] : reg3464[(2'h2):(1'h0)]) ?
              reg3524 : $signed(((reg3508 ? reg3500 : wire3454) ?
                  reg3492 : reg3459))));
          reg3535 <= ($unsigned((("AFusVpYnB36ma" || reg3482[(3'h6):(1'h1)]) | reg3531)) ?
              ((~reg3525) ?
                  $signed($signed((~^(7'h45)))) : "CqXc7oeqKTfYA") : "rolCKSovlh1YkhL1UHL");
        end
      reg3536 <= (~&{($signed(wire3451[(3'h5):(2'h2)]) * reg3478[(2'h3):(2'h3)]),
          ("bPUYd3pZBdi55C4Ti" ?
              $unsigned(((8'hb9) ? reg3457 : reg3518)) : $unsigned(reg3510))});
      for (forvar3537 = (1'h0); (forvar3537 < (2'h2)); forvar3537 = (forvar3537 + (1'h1)))
        begin
          reg3538 <= $unsigned($signed(("biXaV6pGY" ?
              $unsigned({reg3525}) : ($signed(forvar3513) ~^ "IILnC4WFnVTd"))));
          reg3539 <= (reg3461[(4'hb):(4'h9)] | reg3511[(4'h9):(3'h4)]);
          reg3540 <= (+$unsigned((-reg3471)));
          reg3541 <= reg3456[(3'h6):(1'h1)];
          for (forvar3542 = (1'h0); (forvar3542 < (1'h0)); forvar3542 = (forvar3542 + (1'h1)))
            begin
              reg3543 = {{reg3464, (^$signed(reg3478))}, ""};
              reg3544 = {$signed(($signed((reg3536 + reg3505)) >>> "Uf3x3I8OcMkptN1"))};
              reg3545 = (reg3523[(3'h7):(2'h2)] || $signed($unsigned({reg3472,
                  reg3478})));
              for (forvar3546 = (1'h0); (forvar3546 < (2'h3)); forvar3546 = (forvar3546 + (1'h1)))
                begin
                  reg3547 <= (reg3478 << $signed($unsigned((7'h42))));
                  reg3548 <= ((~|$signed(forvar3513[(3'h7):(3'h6)])) << {(reg3505 ?
                          {reg3477[(2'h2):(1'h0)],
                              "YKCYSqKvBfSi"} : (forvar3537 ?
                              "75CrE9PaJf7PAJcZt2" : (~|wire3454))),
                      "2le2Txyv5d"});
                  reg3549 = (((((&reg3530) && (reg3473 ?
                          forvar3542 : reg3511)) <= "xx") != (forvar3487[(4'ha):(2'h2)] & "")) ?
                      {reg3498[(5'h13):(5'h12)],
                          ((-reg3507[(3'h4):(2'h2)]) << (!{reg3484}))} : {reg3530[(2'h2):(1'h1)],
                          (((8'h9d) * forvar3470) ~^ $unsigned("RI50Ef94bWuNtsaIeH2Z"))});
                  reg3550 = (((~|((+reg3463) < (!reg3480))) ?
                      "eRNRzWiabY" : {reg3524,
                          ("UGqhGDvmO" ?
                              $signed(reg3524) : $unsigned((8'h9e)))}) * "");
                end
              for (forvar3551 = (1'h0); (forvar3551 < (3'h5)); forvar3551 = (forvar3551 + (1'h1)))
                begin
                  reg3552 <= (($signed((wire3451[(3'h4):(2'h3)] ?
                          {reg3520, reg3491} : reg3504[(3'h5):(2'h2)])) ?
                      ($unsigned($signed(forvar3551)) + (((8'hb1) <= reg3468) ?
                          ((8'ha9) ?
                              reg3510 : reg3541) : reg3484[(2'h3):(2'h3)])) : reg3520[(3'h4):(2'h2)]) * (~reg3506[(4'he):(2'h2)]));
                  reg3553 <= (~|$signed((8'haf)));
                  reg3554 <= (!$unsigned(((-$unsigned(reg3539)) ?
                      $unsigned({reg3532}) : reg3465[(1'h1):(1'h1)])));
                  reg3555 <= wire3527;
                  reg3556 <= ("LWSex" ? {"7cDOfa"} : $unsigned(reg3552));
                  reg3557 <= (+(forvar3513[(4'h8):(4'h8)] ?
                      "w1k23fEg5JB0Nzs5F6T" : $unsigned(forvar3476[(1'h1):(1'h0)])));
                end
              for (forvar3558 = (1'h0); (forvar3558 < (2'h2)); forvar3558 = (forvar3558 + (1'h1)))
                begin
                  reg3559 = {(8'h9d), reg3484};
                  reg3560 <= forvar3521[(3'h4):(2'h2)];
                end
            end
          reg3561 <= "et904hmRpJsFXCkxS7XVF";
        end
      for (forvar3562 = (1'h0); (forvar3562 < (2'h2)); forvar3562 = (forvar3562 + (1'h1)))
        begin
          reg3563 = forvar3533[(4'hc):(4'ha)];
        end
    end
  assign wire3564 = $signed("VTRY");
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3401
#( parameter param3445 = (|{((~^{(8'ha8), (8'ha4)}) >>> (~((8'haf) || (8'hb8))))})
, parameter param3446 = (((|(~&param3445)) ? {param3445} : {param3445, {(^~(8'haa))}}) << ({param3445} ? {(8'hb8), {(param3445 ? param3445 : param3445), (+param3445)}} : (~{(8'hb3)}))) )
(y, clk, wire3406, wire3405, wire3404, wire3403, wire3402);
  output wire [(32'h216):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire3406;
  input wire signed [(5'h15):(1'h0)] wire3405;
  input wire signed [(4'hb):(1'h0)] wire3404;
  input wire signed [(5'h15):(1'h0)] wire3403;
  input wire [(4'h8):(1'h0)] wire3402;
  reg signed [(4'h9):(1'h0)] reg3444 = (1'h0);
  reg [(5'h13):(1'h0)] reg3443 = (1'h0);
  reg [(4'he):(1'h0)] reg3442 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3441 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3440 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3439 = (1'h0);
  reg [(4'hd):(1'h0)] reg3438 = (1'h0);
  reg [(5'h15):(1'h0)] forvar3437 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3436 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3435 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3434 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3433 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3432 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3431 = (1'h0);
  reg [(3'h6):(1'h0)] reg3430 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3429 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3428 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3427 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3426 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3425 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3424 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3423 = (1'h0);
  reg [(3'h7):(1'h0)] reg3422 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar3421 = (1'h0);
  reg [(2'h2):(1'h0)] reg3420 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3419 = (1'h0);
  reg [(3'h6):(1'h0)] reg3418 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3417 = (1'h0);
  reg [(5'h14):(1'h0)] forvar3416 = (1'h0);
  reg [(5'h19):(1'h0)] reg3415 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar3414 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3413 = (1'h0);
  wire signed [(5'h1a):(1'h0)] wire3412;
  wire signed [(5'h1a):(1'h0)] wire3411;
  reg signed [(2'h3):(1'h0)] reg3410 = (1'h0);
  reg [(3'h6):(1'h0)] reg3409 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3408 = (1'h0);
  reg [(2'h2):(1'h0)] reg3407 = (1'h0);
  assign y = {reg3444,
                 reg3443,
                 reg3442,
                 reg3441,
                 reg3440,
                 reg3439,
                 reg3438,
                 forvar3437,
                 reg3436,
                 reg3435,
                 reg3434,
                 reg3433,
                 reg3432,
                 reg3431,
                 reg3430,
                 forvar3429,
                 reg3428,
                 reg3427,
                 reg3426,
                 forvar3425,
                 reg3424,
                 forvar3423,
                 reg3422,
                 forvar3421,
                 reg3420,
                 reg3419,
                 reg3418,
                 reg3417,
                 forvar3416,
                 reg3415,
                 forvar3414,
                 reg3413,
                 wire3412,
                 wire3411,
                 reg3410,
                 reg3409,
                 reg3408,
                 reg3407,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg3407 <= (({wire3406,
              ($signed((8'ha0)) ? wire3403 : (wire3402 * wire3405))} ?
          (wire3405[(4'ha):(2'h3)] ?
              (8'hb8) : ((~&wire3402) ?
                  $signed(wire3406) : (wire3406 ?
                      wire3402 : (7'h40)))) : ($unsigned((~|wire3404)) ?
              ((wire3402 ?
                  wire3403 : wire3403) == ((8'hab) << wire3405)) : $unsigned("kVRrVDAQ2eA"))) <<< wire3406[(2'h2):(1'h1)]);
      reg3408 <= "tfsBBnVh";
      reg3409 <= $unsigned((8'haf));
      reg3410 <= (($signed((reg3407 ?
              $unsigned(wire3404) : (wire3404 ^~ wire3404))) * reg3407[(2'h2):(1'h0)]) ?
          wire3406 : (8'ha1));
    end
  assign wire3411 = wire3405;
  assign wire3412 = {$signed($unsigned($unsigned($unsigned(reg3409))))};
  always
    @(posedge clk) begin
      reg3413 <= "8MfCdQZeTICi";
      for (forvar3414 = (1'h0); (forvar3414 < (3'h4)); forvar3414 = (forvar3414 + (1'h1)))
        begin
          reg3415 = $signed((("h3" ?
              (wire3406 > (reg3408 ?
                  reg3407 : (7'h42))) : "cadeLObuHFEQelrvWdOFe") * ($signed(wire3402[(1'h1):(1'h1)]) ?
              wire3406 : "")));
          for (forvar3416 = (1'h0); (forvar3416 < (1'h1)); forvar3416 = (forvar3416 + (1'h1)))
            begin
              reg3417 = reg3410;
              reg3418 <= {reg3409[(1'h1):(1'h1)],
                  ((&wire3405) >>> reg3410[(2'h3):(2'h3)])};
              reg3419 <= $unsigned(reg3407[(1'h0):(1'h0)]);
              reg3420 <= wire3412[(5'h1a):(3'h6)];
            end
          for (forvar3421 = (1'h0); (forvar3421 < (1'h0)); forvar3421 = (forvar3421 + (1'h1)))
            begin
              reg3422 <= $signed((reg3410 + reg3419));
            end
          for (forvar3423 = (1'h0); (forvar3423 < (3'h4)); forvar3423 = (forvar3423 + (1'h1)))
            begin
              reg3424 <= "xFU7345F1k4bonifW";
              for (forvar3425 = (1'h0); (forvar3425 < (3'h5)); forvar3425 = (forvar3425 + (1'h1)))
                begin
                  reg3426 = forvar3414;
                  reg3427 <= forvar3425;
                  reg3428 <= wire3406[(3'h5):(2'h3)];
                end
              for (forvar3429 = (1'h0); (forvar3429 < (3'h4)); forvar3429 = (forvar3429 + (1'h1)))
                begin
                  reg3430 = reg3415;
                  reg3431 <= $unsigned(forvar3416);
                end
              reg3432 <= $unsigned($unsigned(($unsigned($unsigned(reg3430)) <= $unsigned({forvar3421,
                  reg3418}))));
              reg3433 <= "7ZrKbk0avqdK";
              reg3434 <= ({((&{reg3415}) - ($signed(reg3420) ?
                      reg3431 : reg3418[(1'h0):(1'h0)]))} - (~|reg3415[(5'h16):(5'h16)]));
            end
          reg3435 <= (+($unsigned("XdRZZTnS3J5cRPPuGVxI") & ("ftTf7tAbUDLisknW28KY3R" ?
              ($unsigned(reg3417) ?
                  "tWBbn0zE7JlV4" : $unsigned(forvar3425)) : ((&reg3424) >= reg3422))));
          reg3436 = {{{$unsigned((wire3404 > reg3415))}}};
        end
      for (forvar3437 = (1'h0); (forvar3437 < (3'h5)); forvar3437 = (forvar3437 + (1'h1)))
        begin
          reg3438 <= "vfx";
          reg3439 = (~^forvar3416);
          reg3440 = ($unsigned((forvar3425[(2'h3):(2'h2)] & $unsigned((~^forvar3425)))) <= $unsigned((forvar3437 || reg3417)));
        end
      reg3441 <= wire3412;
    end
  always
    @(posedge clk) begin
      reg3442 <= (((((~|(8'hba)) ?
              {(8'hbd)} : $unsigned(reg3422)) >>> forvar3414) ^~ (("iFLiIWZZelHhqyvSvu" < $signed(forvar3437)) ?
              reg3419 : wire3411)) ?
          $unsigned(reg3410) : "PRyqX");
      reg3443 <= (|(|((~^wire3402) ?
          {forvar3423} : ("LEkuNoCZ0ODepFPVN7pN7Y" >> forvar3416[(3'h4):(2'h3)]))));
      reg3444 <= reg3422[(3'h4):(2'h3)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3204
#( parameter param3397 = (|((({(8'hb1)} ? ((7'h41) ? (8'hb2) : (8'hb2)) : ((7'h49) ? (8'ha8) : (8'had))) ? {((7'h41) ? (8'hbf) : (8'hac))} : ((~&(8'hb4)) ? {(8'ha7), (7'h40)} : (&(8'hbd)))) ? ((|((7'h47) ? (7'h47) : (8'hbe))) ^ (+(&(7'h4c)))) : ((((7'h43) < (8'haa)) ? ((8'haa) || (8'hbb)) : ((7'h49) ? (8'hbd) : (7'h44))) ? (((7'h42) ? (8'hb7) : (8'had)) >>> ((7'h46) >>> (7'h40))) : (~|(&(8'hb6))))))
, parameter param3398 = (((param3397 ? (|(param3397 ? param3397 : param3397)) : ({param3397, param3397} ? (param3397 + param3397) : param3397)) ? (7'h44) : (((~&param3397) ? param3397 : (param3397 ^~ param3397)) != (~|(param3397 << param3397)))) ^~ ((~^param3397) != {(~^(param3397 ? (8'haf) : param3397)), ((param3397 ? param3397 : param3397) ? ((8'hb1) - param3397) : (^param3397))})) )
(y, clk, wire3208, wire3207, wire3206, wire3205);
  output wire [(32'ha2e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire3208;
  input wire signed [(5'h19):(1'h0)] wire3207;
  input wire signed [(4'h8):(1'h0)] wire3206;
  input wire signed [(5'h17):(1'h0)] wire3205;
  wire signed [(4'hc):(1'h0)] wire3396;
  reg signed [(4'hd):(1'h0)] reg3395 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3394 = (1'h0);
  reg [(4'he):(1'h0)] reg3393 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3392 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3391 = (1'h0);
  reg [(5'h15):(1'h0)] reg3390 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3389 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3388 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3387 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3386 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3385 = (1'h0);
  reg [(5'h10):(1'h0)] reg3384 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3383 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3382 = (1'h0);
  reg [(5'h18):(1'h0)] reg3381 = (1'h0);
  reg [(5'h13):(1'h0)] reg3380 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar3379 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3378 = (1'h0);
  reg [(5'h18):(1'h0)] forvar3377 = (1'h0);
  reg [(4'ha):(1'h0)] reg3376 = (1'h0);
  reg [(4'h8):(1'h0)] reg3375 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3374 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3373 = (1'h0);
  reg [(2'h2):(1'h0)] reg3372 = (1'h0);
  reg [(5'h18):(1'h0)] reg3371 = (1'h0);
  reg [(3'h6):(1'h0)] reg3370 = (1'h0);
  reg [(4'he):(1'h0)] reg3369 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3368 = (1'h0);
  reg [(3'h4):(1'h0)] reg3367 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3366 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3365 = (1'h0);
  reg [(4'ha):(1'h0)] reg3364 = (1'h0);
  reg [(5'h16):(1'h0)] reg3363 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3362 = (1'h0);
  wire signed [(5'h19):(1'h0)] wire3361;
  reg [(3'h5):(1'h0)] reg3360 = (1'h0);
  reg [(3'h4):(1'h0)] reg3359 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3358 = (1'h0);
  reg [(5'h10):(1'h0)] reg3357 = (1'h0);
  reg [(4'hc):(1'h0)] reg3356 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3355 = (1'h0);
  reg [(4'hd):(1'h0)] reg3354 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3353 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3352 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3351 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3350 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar3349 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3348 = (1'h0);
  reg [(5'h14):(1'h0)] forvar3347 = (1'h0);
  reg [(5'h12):(1'h0)] reg3346 = (1'h0);
  reg [(3'h4):(1'h0)] reg3345 = (1'h0);
  reg [(4'hb):(1'h0)] reg3344 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3343 = (1'h0);
  reg [(5'h11):(1'h0)] reg3342 = (1'h0);
  reg [(4'ha):(1'h0)] reg3341 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3340 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3339 = (1'h0);
  reg [(5'h13):(1'h0)] reg3338 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3337 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3336 = (1'h0);
  reg [(2'h2):(1'h0)] reg3335 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3334 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3333 = (1'h0);
  reg [(4'ha):(1'h0)] reg3332 = (1'h0);
  reg [(4'hf):(1'h0)] reg3331 = (1'h0);
  reg [(5'h10):(1'h0)] reg3330 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3329 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3328 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3327 = (1'h0);
  reg [(5'h10):(1'h0)] reg3326 = (1'h0);
  reg [(5'h18):(1'h0)] forvar3325 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3324 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3323 = (1'h0);
  reg [(2'h2):(1'h0)] reg3322 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3321 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar3320 = (1'h0);
  reg [(4'he):(1'h0)] reg3319 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3318 = (1'h0);
  reg [(2'h2):(1'h0)] reg3317 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3316 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3315 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3314 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3313 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3312 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3311 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3310 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar3309 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire3308;
  reg signed [(5'h12):(1'h0)] reg3307 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3306 = (1'h0);
  reg [(4'hf):(1'h0)] reg3305 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3304 = (1'h0);
  reg [(5'h17):(1'h0)] reg3303 = (1'h0);
  reg [(5'h17):(1'h0)] reg3302 = (1'h0);
  reg [(3'h6):(1'h0)] reg3301 = (1'h0);
  reg [(3'h5):(1'h0)] reg3300 = (1'h0);
  reg [(2'h2):(1'h0)] reg3299 = (1'h0);
  reg [(4'ha):(1'h0)] reg3298 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3297 = (1'h0);
  reg [(5'h10):(1'h0)] reg3296 = (1'h0);
  reg [(5'h17):(1'h0)] forvar3295 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3294 = (1'h0);
  reg [(5'h10):(1'h0)] reg3293 = (1'h0);
  reg [(4'he):(1'h0)] reg3280 = (1'h0);
  reg [(4'hd):(1'h0)] reg3292 = (1'h0);
  reg [(4'h8):(1'h0)] reg3291 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3290 = (1'h0);
  reg [(5'h16):(1'h0)] reg3289 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3288 = (1'h0);
  reg [(5'h14):(1'h0)] reg3287 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3286 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3285 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3284 = (1'h0);
  reg [(5'h14):(1'h0)] reg3283 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3282 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3281 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar3280 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3279 = (1'h0);
  reg [(3'h4):(1'h0)] reg3278 = (1'h0);
  reg [(5'h14):(1'h0)] forvar3277 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3276 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3275 = (1'h0);
  reg [(5'h12):(1'h0)] forvar3274 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3273 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3272 = (1'h0);
  reg [(4'he):(1'h0)] reg3271 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3270 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3269 = (1'h0);
  reg [(5'h15):(1'h0)] forvar3268 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3267 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3266 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3265 = (1'h0);
  reg [(5'h11):(1'h0)] reg3264 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3263 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3262 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3261 = (1'h0);
  reg [(5'h11):(1'h0)] reg3260 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3259 = (1'h0);
  reg [(4'hd):(1'h0)] reg3258 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3257 = (1'h0);
  reg [(4'he):(1'h0)] reg3256 = (1'h0);
  reg [(5'h11):(1'h0)] reg3255 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3254 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar3253 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3252 = (1'h0);
  reg [(3'h4):(1'h0)] reg3251 = (1'h0);
  reg [(5'h16):(1'h0)] forvar3250 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3249 = (1'h0);
  reg [(5'h17):(1'h0)] reg3248 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3247 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3246 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3245 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3244 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3243 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3242 = (1'h0);
  reg [(3'h6):(1'h0)] reg3241 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3240 = (1'h0);
  reg [(5'h11):(1'h0)] reg3239 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3238 = (1'h0);
  reg [(5'h14):(1'h0)] forvar3237 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3236 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3235 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3234 = (1'h0);
  reg [(2'h2):(1'h0)] reg3233 = (1'h0);
  reg [(5'h18):(1'h0)] reg3232 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3231 = (1'h0);
  reg [(4'he):(1'h0)] forvar3230 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar3229 = (1'h0);
  reg [(2'h3):(1'h0)] reg3228 = (1'h0);
  reg [(3'h6):(1'h0)] reg3227 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3226 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar3225 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3224 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar3223 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar3222 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire3221;
  wire signed [(5'h12):(1'h0)] wire3220;
  reg [(3'h6):(1'h0)] reg3219 = (1'h0);
  reg [(3'h6):(1'h0)] reg3218 = (1'h0);
  reg [(3'h7):(1'h0)] reg3217 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3216 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3215 = (1'h0);
  reg [(3'h7):(1'h0)] reg3214 = (1'h0);
  reg [(4'hd):(1'h0)] reg3213 = (1'h0);
  reg [(5'h11):(1'h0)] forvar3212 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3211 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3210 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar3209 = (1'h0);
  assign y = {wire3396,
                 reg3395,
                 reg3394,
                 reg3393,
                 reg3392,
                 forvar3391,
                 reg3390,
                 reg3389,
                 reg3388,
                 reg3387,
                 reg3386,
                 reg3385,
                 reg3384,
                 reg3383,
                 reg3382,
                 reg3381,
                 reg3380,
                 forvar3379,
                 reg3378,
                 forvar3377,
                 reg3376,
                 reg3375,
                 forvar3374,
                 reg3373,
                 reg3372,
                 reg3371,
                 reg3370,
                 reg3369,
                 reg3368,
                 reg3367,
                 reg3366,
                 forvar3365,
                 reg3364,
                 reg3363,
                 forvar3362,
                 wire3361,
                 reg3360,
                 reg3359,
                 reg3358,
                 reg3357,
                 reg3356,
                 reg3355,
                 reg3354,
                 reg3353,
                 reg3352,
                 reg3351,
                 reg3350,
                 forvar3349,
                 reg3348,
                 forvar3347,
                 reg3346,
                 reg3345,
                 reg3344,
                 reg3343,
                 reg3342,
                 reg3341,
                 reg3340,
                 reg3339,
                 reg3338,
                 forvar3337,
                 forvar3336,
                 reg3335,
                 reg3334,
                 forvar3333,
                 reg3332,
                 reg3331,
                 reg3330,
                 reg3329,
                 reg3328,
                 reg3327,
                 reg3326,
                 forvar3325,
                 forvar3324,
                 reg3323,
                 reg3322,
                 reg3321,
                 forvar3320,
                 reg3319,
                 reg3318,
                 reg3317,
                 reg3316,
                 reg3315,
                 reg3314,
                 reg3313,
                 reg3312,
                 reg3311,
                 reg3310,
                 forvar3309,
                 wire3308,
                 reg3307,
                 reg3306,
                 reg3305,
                 reg3304,
                 reg3303,
                 reg3302,
                 reg3301,
                 reg3300,
                 reg3299,
                 reg3298,
                 forvar3297,
                 reg3296,
                 forvar3295,
                 forvar3294,
                 reg3293,
                 reg3280,
                 reg3292,
                 reg3291,
                 reg3290,
                 reg3289,
                 reg3288,
                 reg3287,
                 reg3286,
                 forvar3285,
                 reg3284,
                 reg3283,
                 reg3282,
                 reg3281,
                 forvar3280,
                 reg3279,
                 reg3278,
                 forvar3277,
                 reg3276,
                 reg3275,
                 forvar3274,
                 reg3273,
                 reg3272,
                 reg3271,
                 reg3270,
                 forvar3269,
                 forvar3268,
                 reg3267,
                 reg3266,
                 reg3265,
                 reg3264,
                 reg3263,
                 reg3262,
                 reg3261,
                 reg3260,
                 reg3259,
                 reg3258,
                 reg3257,
                 reg3256,
                 reg3255,
                 reg3254,
                 forvar3253,
                 reg3252,
                 reg3251,
                 forvar3250,
                 reg3249,
                 reg3248,
                 reg3247,
                 reg3246,
                 reg3245,
                 forvar3244,
                 forvar3243,
                 reg3242,
                 reg3241,
                 reg3240,
                 reg3239,
                 reg3238,
                 forvar3237,
                 reg3236,
                 reg3235,
                 reg3234,
                 reg3233,
                 reg3232,
                 reg3231,
                 forvar3230,
                 forvar3229,
                 reg3228,
                 reg3227,
                 reg3226,
                 forvar3225,
                 reg3224,
                 forvar3223,
                 forvar3222,
                 wire3221,
                 wire3220,
                 reg3219,
                 reg3218,
                 reg3217,
                 reg3216,
                 reg3215,
                 reg3214,
                 reg3213,
                 forvar3212,
                 reg3211,
                 reg3210,
                 forvar3209,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar3209 = (1'h0); (forvar3209 < (1'h1)); forvar3209 = (forvar3209 + (1'h1)))
        begin
          reg3210 = (wire3207 <= $signed($unsigned(wire3206)));
          reg3211 <= (|(^~$signed((wire3208[(4'he):(4'hb)] * wire3207))));
          for (forvar3212 = (1'h0); (forvar3212 < (3'h4)); forvar3212 = (forvar3212 + (1'h1)))
            begin
              reg3213 <= {(8'hab)};
              reg3214 = $signed(forvar3209[(3'h4):(2'h3)]);
              reg3215 <= wire3207;
              reg3216 <= ((reg3213[(1'h1):(1'h0)] != "W") < forvar3209[(3'h4):(1'h0)]);
            end
        end
      reg3217 <= $unsigned(((+reg3214[(3'h4):(1'h0)]) ?
          wire3206[(2'h3):(1'h0)] : $signed((forvar3212[(3'h7):(1'h0)] ?
              "Q5" : (reg3214 ? (8'hb9) : wire3205)))));
      reg3218 <= $unsigned((^~$unsigned($signed(reg3215[(1'h0):(1'h0)]))));
      reg3219 <= $unsigned(($signed(reg3210[(5'h12):(3'h6)]) ?
          ((+wire3205) ?
              (forvar3212[(5'h11):(4'h9)] ?
                  (~&reg3213) : reg3218) : wire3208) : ((~|(reg3215 ?
              reg3216 : wire3208)) << $signed({reg3215, reg3217}))));
    end
  assign wire3220 = wire3207;
  assign wire3221 = (|(8'hac));
  always
    @(posedge clk) begin
      for (forvar3222 = (1'h0); (forvar3222 < (3'h4)); forvar3222 = (forvar3222 + (1'h1)))
        begin
          for (forvar3223 = (1'h0); (forvar3223 < (3'h5)); forvar3223 = (forvar3223 + (1'h1)))
            begin
              reg3224 <= wire3206;
              for (forvar3225 = (1'h0); (forvar3225 < (1'h0)); forvar3225 = (forvar3225 + (1'h1)))
                begin
                  reg3226 = (((((reg3214 >> reg3210) ?
                          forvar3223 : $unsigned(forvar3225)) ^ ((|forvar3222) ?
                          $signed(wire3208) : "4cvPVnJzgUPE72O4ZMZZLx9Gk")) >> (~wire3208)) ?
                      reg3215[(2'h3):(1'h1)] : (^forvar3225[(4'hc):(4'h9)]));
                  reg3227 = wire3205[(4'hd):(4'hb)];
                end
            end
          reg3228 <= (wire3220 ? $unsigned($unsigned("fFqPB5sPz2oT8ME")) : "M");
          for (forvar3229 = (1'h0); (forvar3229 < (3'h4)); forvar3229 = (forvar3229 + (1'h1)))
            begin
              for (forvar3230 = (1'h0); (forvar3230 < (1'h0)); forvar3230 = (forvar3230 + (1'h1)))
                begin
                  reg3231 <= reg3218;
                  reg3232 <= reg3226;
                  reg3233 <= (~&("Qv8y6twecrN1" != (((~^reg3227) & {reg3218}) * ($unsigned(wire3221) >>> reg3210))));
                  reg3234 = ((8'ha2) == (~&$unsigned(reg3213[(2'h3):(2'h2)])));
                  reg3235 = (^~$signed(($signed($unsigned(reg3224)) ?
                      reg3216 : ($signed(reg3210) ?
                          ((7'h40) ?
                              reg3213 : wire3206) : $unsigned(reg3213)))));
                  reg3236 = $signed((+reg3232[(3'h6):(1'h0)]));
                end
              for (forvar3237 = (1'h0); (forvar3237 < (3'h4)); forvar3237 = (forvar3237 + (1'h1)))
                begin
                  reg3238 <= forvar3225;
                  reg3239 <= $signed(reg3213);
                  reg3240 <= reg3231[(4'hd):(3'h4)];
                  reg3241 <= $unsigned(((|((wire3208 ? wire3220 : reg3235) ?
                          $signed(reg3217) : "mg8o")) ?
                      (forvar3212[(4'hd):(2'h2)] ?
                          reg3213[(3'h6):(3'h6)] : $unsigned($unsigned(reg3219))) : reg3236));
                  reg3242 <= {($unsigned($signed(reg3211)) * reg3224[(2'h3):(2'h3)])};
                end
            end
        end
      for (forvar3243 = (1'h0); (forvar3243 < (3'h5)); forvar3243 = (forvar3243 + (1'h1)))
        begin
          for (forvar3244 = (1'h0); (forvar3244 < (3'h4)); forvar3244 = (forvar3244 + (1'h1)))
            begin
              reg3245 <= reg3226;
              reg3246 <= (($unsigned(forvar3225[(1'h0):(1'h0)]) ^~ (~^(!forvar3229))) ?
                  (($unsigned(wire3205) - reg3226[(2'h3):(1'h0)]) + (-"Ta6R7zM")) : reg3245[(1'h1):(1'h1)]);
              reg3247 <= forvar3230;
              reg3248 = $unsigned((reg3245[(1'h0):(1'h0)] ?
                  {"rNw2z6x2wnxKY9",
                      reg3219} : ("KaO2OiMmxrzmcoUIa3Z9" <<< "Z9UMKdDq5rlqPguMbtXJYLFn")));
            end
          reg3249 <= $unsigned(reg3226);
          for (forvar3250 = (1'h0); (forvar3250 < (3'h5)); forvar3250 = (forvar3250 + (1'h1)))
            begin
              reg3251 <= (~^$signed((reg3246 ? "GxkNpvVWYHf" : (8'hbf))));
              reg3252 = {(forvar3225[(3'h7):(1'h1)] || $unsigned(((forvar3209 < wire3220) ?
                      $unsigned(reg3233) : reg3217[(1'h0):(1'h0)])))};
              for (forvar3253 = (1'h0); (forvar3253 < (3'h5)); forvar3253 = (forvar3253 + (1'h1)))
                begin
                  reg3254 <= "mHNHf28KgQat";
                  reg3255 = reg3233;
                  reg3256 = reg3228;
                  reg3257 <= ($signed((~forvar3209)) ^ ((^~reg3238) < $signed((~^$unsigned(reg3245)))));
                  reg3258 <= (-"wdcPk");
                end
              reg3259 <= reg3231[(4'ha):(2'h3)];
            end
          reg3260 <= (&"1ZXN");
          reg3261 <= $signed("0");
        end
      reg3262 <= (7'h40);
      reg3263 <= $unsigned(("sf" ? "viJf" : reg3252));
      reg3264 <= forvar3225[(3'h5):(2'h3)];
      reg3265 <= $unsigned($signed({(&(8'hba)), {(!reg3214)}}));
    end
  always
    @(posedge clk) begin
      reg3266 <= reg3231;
      reg3267 = reg3232;
      for (forvar3268 = (1'h0); (forvar3268 < (2'h2)); forvar3268 = (forvar3268 + (1'h1)))
        begin
          for (forvar3269 = (1'h0); (forvar3269 < (2'h3)); forvar3269 = (forvar3269 + (1'h1)))
            begin
              reg3270 <= reg3239[(4'ha):(4'h8)];
            end
          reg3271 <= {($unsigned($signed((&reg3235))) ?
                  (forvar3225 ?
                      reg3265[(1'h1):(1'h0)] : forvar3212[(3'h4):(3'h4)]) : (|{{reg3249},
                      (8'hbc)}))};
        end
      reg3272 <= (wire3206[(3'h4):(2'h3)] ?
          "dp21V5g0agf3Dzmp0e" : (wire3220 ?
              "ooRGm7cAWaUeAW2dn" : (-(|(reg3231 <<< reg3267)))));
      reg3273 <= ($unsigned("i3Jzd8NMVGclJshv") * $signed((reg3247[(3'h4):(3'h4)] ?
          $unsigned((^~forvar3244)) : reg3261[(3'h7):(1'h0)])));
    end
  always
    @(posedge clk) begin
      for (forvar3274 = (1'h0); (forvar3274 < (1'h0)); forvar3274 = (forvar3274 + (1'h1)))
        begin
          reg3275 <= ($signed($signed((|reg3254[(3'h7):(3'h7)]))) ^~ reg3266[(1'h0):(1'h0)]);
          reg3276 = reg3267;
        end
      for (forvar3277 = (1'h0); (forvar3277 < (2'h2)); forvar3277 = (forvar3277 + (1'h1)))
        begin
          reg3278 <= $signed(forvar3225[(4'hc):(4'h9)]);
          if ((^$unsigned(((reg3211[(5'h14):(3'h5)] ? (~reg3260) : {reg3246}) ?
              ({reg3259} == (~&(8'ha4))) : reg3262))))
            begin
              reg3279 <= ($unsigned({$unsigned($signed(forvar3250))}) ^ $signed(reg3276[(4'hd):(4'hc)]));
              for (forvar3280 = (1'h0); (forvar3280 < (1'h1)); forvar3280 = (forvar3280 + (1'h1)))
                begin
                  reg3281 = "OeVc8GusIr";
                  reg3282 = $signed((~|$unsigned({(reg3247 ?
                          (8'hac) : reg3249)})));
                  reg3283 = wire3208;
                  reg3284 = (~|(+(("m9hiE5FZxkYURHGJR" | (^~(7'h4c))) ?
                      (reg3226[(3'h4):(1'h0)] <<< reg3233) : (-reg3255[(4'hd):(4'h9)]))));
                end
              for (forvar3285 = (1'h0); (forvar3285 < (2'h3)); forvar3285 = (forvar3285 + (1'h1)))
                begin
                  reg3286 = $unsigned((forvar3243 ?
                      "J2vc8LAgqBwy" : $signed(((~&reg3259) == forvar3253[(2'h2):(1'h1)]))));
                  reg3287 <= $unsigned($unsigned("KGQD9LGmNGTcs"));
                  reg3288 <= (8'hb0);
                  reg3289 <= $unsigned(((({reg3282, reg3257} ?
                          (reg3217 ? forvar3222 : wire3206) : forvar3223) ?
                      (^~$unsigned(forvar3268)) : reg3227) != (reg3262[(4'ha):(2'h2)] ?
                      ("ZgDHanF4Wal2" & "YELzKLf") : reg3284[(4'hb):(4'hb)])));
                  reg3290 <= $signed($unsigned(({((8'h9f) ?
                              wire3220 : (7'h4a))} ?
                      (~(-reg3271)) : (~reg3226[(4'ha):(3'h4)]))));
                end
              reg3291 <= (|("mbMhoV" <<< "cqFfbFuXGqVtq"));
              reg3292 <= "Tx";
            end
          else
            begin
              reg3279 <= {(8'ha1)};
              reg3280 <= reg3256;
            end
        end
      reg3293 = (!$unsigned(reg3288));
      for (forvar3294 = (1'h0); (forvar3294 < (2'h2)); forvar3294 = (forvar3294 + (1'h1)))
        begin
          for (forvar3295 = (1'h0); (forvar3295 < (2'h2)); forvar3295 = (forvar3295 + (1'h1)))
            begin
              reg3296 <= (reg3211[(3'h5):(2'h2)] ^ (($signed("Mdp4Sc") != forvar3268[(2'h3):(1'h1)]) == $signed("X3XfILv3")));
              for (forvar3297 = (1'h0); (forvar3297 < (2'h2)); forvar3297 = (forvar3297 + (1'h1)))
                begin
                  reg3298 <= reg3224[(3'h6):(3'h5)];
                  reg3299 <= (~$unsigned((~&{"QIXxb"})));
                  reg3300 = (+(reg3283[(4'hc):(2'h3)] ?
                      wire3207 : reg3242[(1'h0):(1'h0)]));
                end
              reg3301 <= ((&$unsigned(reg3300)) < $unsigned(forvar3280[(4'he):(3'h7)]));
              reg3302 <= (7'h48);
              reg3303 <= forvar3229;
              reg3304 <= (reg3256[(3'h4):(2'h3)] >>> {$signed(reg3242)});
            end
          reg3305 = ((wire3208[(2'h2):(1'h1)] ?
              {reg3234,
                  forvar3297[(1'h1):(1'h1)]} : wire3207[(4'ha):(1'h1)]) - ("yt3VZJt2Z6f" ?
              "qy1IigpTFkynlnsJynmO" : {"iGxnYRswuSaysyJ8osrDaU"}));
          reg3306 <= reg3266[(2'h3):(2'h2)];
        end
      reg3307 <= $signed(forvar3225[(3'h4):(2'h2)]);
    end
  assign wire3308 = $signed((+"w5E3P"));
  always
    @(posedge clk) begin
      for (forvar3309 = (1'h0); (forvar3309 < (2'h2)); forvar3309 = (forvar3309 + (1'h1)))
        begin
          reg3310 <= (reg3267 << {"OO7mQDFgQWGSVzMkY0uaMLcMr"});
          reg3311 <= "bL";
          reg3312 <= $unsigned((~^((~$signed(forvar3294)) ?
              (~&$unsigned((8'hb4))) : (-reg3307[(4'hb):(2'h3)]))));
          reg3313 <= {"mhB0Z0lym8vvBlUlSO"};
          reg3314 <= {(reg3271 ?
                  $signed($unsigned(((8'haf) ?
                      reg3300 : reg3265))) : $signed((~|(reg3291 ?
                      reg3215 : reg3235)))),
              reg3313};
        end
    end
  always
    @(posedge clk) begin
      reg3315 <= forvar3285;
      reg3316 <= (-("ifPCVSbxCR" ?
          ($signed($unsigned(wire3208)) ?
              {reg3314[(4'h8):(3'h4)],
                  $signed((7'h4d))} : ((forvar3274 >>> reg3226) + "xBgQXnnXHCOdwTJzX9pE")) : ($unsigned(reg3279[(4'h9):(1'h0)]) ~^ reg3216)));
      reg3317 <= forvar3280[(5'h11):(3'h6)];
      reg3318 <= (forvar3244[(4'hc):(1'h0)] ?
          $unsigned("YwiNFub1LK6YxlckV") : (~&forvar3250[(5'h11):(4'h9)]));
    end
  always
    @(posedge clk) begin
      reg3319 = (forvar3209 ^ reg3210[(5'h14):(5'h10)]);
      for (forvar3320 = (1'h0); (forvar3320 < (3'h4)); forvar3320 = (forvar3320 + (1'h1)))
        begin
          reg3321 = $unsigned((|$signed(wire3206)));
          reg3322 <= {(reg3275 ^~ {"0oBMteZytzQU2N",
                  ((reg3264 ? reg3241 : reg3238) ?
                      (|(7'h49)) : reg3282[(5'h15):(5'h14)])}),
              $unsigned(({(^reg3231),
                  (reg3242 ? reg3228 : (7'h41))} ^~ {$signed(forvar3223)}))};
          reg3323 <= forvar3320;
          for (forvar3324 = (1'h0); (forvar3324 < (2'h2)); forvar3324 = (forvar3324 + (1'h1)))
            begin
              for (forvar3325 = (1'h0); (forvar3325 < (2'h2)); forvar3325 = (forvar3325 + (1'h1)))
                begin
                  reg3326 <= ($unsigned({"3WKqlGENmX2AOi2cRo"}) ?
                      $unsigned(reg3239) : "DKiGfDkgu");
                  reg3327 <= {"8p4gs5"};
                end
              reg3328 <= $unsigned(reg3310[(4'h8):(3'h5)]);
            end
          reg3329 <= (8'hb1);
        end
      reg3330 <= wire3208;
      reg3331 <= reg3288;
      reg3332 <= (~^$unsigned((~|forvar3285)));
    end
  always
    @(posedge clk) begin
      for (forvar3333 = (1'h0); (forvar3333 < (3'h5)); forvar3333 = (forvar3333 + (1'h1)))
        begin
          reg3334 <= ($signed(($unsigned($unsigned(reg3234)) ?
              wire3220 : "pPgpaGFfCni3RNLnT8")) + (^~(reg3264 > reg3322[(1'h0):(1'h0)])));
        end
      reg3335 <= "B0H9ArJ8NXAL3iRZ6dh7C";
      for (forvar3336 = (1'h0); (forvar3336 < (2'h3)); forvar3336 = (forvar3336 + (1'h1)))
        begin
          for (forvar3337 = (1'h0); (forvar3337 < (1'h0)); forvar3337 = (forvar3337 + (1'h1)))
            begin
              reg3338 <= reg3213[(4'hd):(4'hb)];
              reg3339 <= "5efzwBcUkA4cZ";
              reg3340 <= $unsigned(($unsigned($unsigned($signed(reg3236))) ?
                  $unsigned(((~|(7'h42)) == reg3255[(3'h5):(1'h1)])) : $signed({$signed(reg3224)})));
            end
          reg3341 <= forvar3250[(4'hc):(1'h1)];
          reg3342 <= $unsigned(forvar3297);
          reg3343 <= "Qlr5JIPvY";
          reg3344 <= ((~^$signed(("qnP" <<< (|reg3249)))) || "B25rKFu4bMxcRJisMl");
        end
      reg3345 <= $unsigned($signed(reg3286));
    end
  always
    @(posedge clk) begin
      reg3346 = {reg3328, reg3310};
      for (forvar3347 = (1'h0); (forvar3347 < (3'h5)); forvar3347 = (forvar3347 + (1'h1)))
        begin
          reg3348 <= ($unsigned($signed(forvar3269[(3'h5):(3'h5)])) & (+((forvar3250[(3'h6):(1'h0)] && $unsigned(reg3326)) ?
              (7'h41) : reg3303)));
          for (forvar3349 = (1'h0); (forvar3349 < (1'h1)); forvar3349 = (forvar3349 + (1'h1)))
            begin
              reg3350 = $unsigned((reg3344[(3'h4):(1'h1)] ?
                  ((reg3275[(1'h1):(1'h1)] ? $unsigned(reg3259) : reg3335) ?
                      reg3267 : ((reg3338 <<< reg3346) - (forvar3225 ?
                          reg3228 : reg3267))) : "beRkYU63478JXvzU"));
              reg3351 <= reg3249;
              reg3352 = reg3245;
            end
        end
      reg3353 = (reg3232[(4'hc):(2'h2)] ?
          forvar3347[(4'hd):(4'h9)] : "fVUGH75DrYGoFp");
      reg3354 <= reg3278[(2'h2):(1'h0)];
      reg3355 <= "sQxsgESvE7pci";
      reg3356 = ({"Nc1z"} * (reg3331 ^ reg3241));
    end
  always
    @(posedge clk) begin
      reg3357 <= ((reg3302 & $unsigned(($unsigned((8'hbf)) ?
          reg3279[(5'h10):(4'he)] : ((7'h47) ?
              forvar3320 : reg3245)))) > forvar3253);
      reg3358 <= reg3258;
      reg3359 <= ({(~^"ISwMTUyq7qTqBivF")} <= forvar3209[(4'hc):(3'h4)]);
      reg3360 <= ("a7Quh" ?
          "lEYipwlZnLQyIPtpFLdTnACVO" : $unsigned(reg3281[(4'hc):(1'h1)]));
    end
  assign wire3361 = ((reg3339 >> $signed((~&{forvar3277}))) ~^ (!({reg3258[(3'h7):(2'h3)]} ?
                        ("OGHvMqUTwvQn19sdee0lD" * reg3355[(4'he):(3'h7)]) : "Fr")));
  always
    @(posedge clk) begin
      for (forvar3362 = (1'h0); (forvar3362 < (1'h0)); forvar3362 = (forvar3362 + (1'h1)))
        begin
          reg3363 <= $signed((^~"a"));
          reg3364 <= (-$unsigned((reg3266[(3'h7):(2'h3)] == $signed((reg3342 ?
              reg3278 : reg3327)))));
          for (forvar3365 = (1'h0); (forvar3365 < (2'h2)); forvar3365 = (forvar3365 + (1'h1)))
            begin
              reg3366 <= reg3357[(4'hf):(3'h5)];
              reg3367 <= $signed("NP0HQyfeXWJqPw");
              reg3368 <= forvar3336[(1'h1):(1'h1)];
              reg3369 <= $signed($unsigned((^"2aucwDBNhm9c")));
            end
          reg3370 <= ((|$unsigned(("" && "4v54mVytnEzPy6"))) * reg3300[(1'h1):(1'h1)]);
          reg3371 = $signed($unsigned(reg3366));
        end
      reg3372 = ((|reg3307) != $signed(forvar3268[(5'h10):(3'h4)]));
      reg3373 = forvar3250[(4'hc):(4'hb)];
      for (forvar3374 = (1'h0); (forvar3374 < (3'h4)); forvar3374 = (forvar3374 + (1'h1)))
        begin
          reg3375 <= (8'hba);
          reg3376 <= {forvar3309};
        end
      for (forvar3377 = (1'h0); (forvar3377 < (1'h1)); forvar3377 = (forvar3377 + (1'h1)))
        begin
          reg3378 <= "scD";
        end
    end
  always
    @(posedge clk) begin
      for (forvar3379 = (1'h0); (forvar3379 < (2'h2)); forvar3379 = (forvar3379 + (1'h1)))
        begin
          reg3380 <= $signed($signed({$signed((forvar3253 ?
                  reg3296 : forvar3229))}));
          reg3381 <= reg3264[(1'h1):(1'h0)];
          reg3382 <= $unsigned((&$signed("rNGYgXmNOoYdEcB")));
          reg3383 <= reg3380;
        end
      reg3384 <= ((($unsigned($signed(forvar3337)) ?
              ("BGbmlRn6WXy12fKIEzY" ? reg3364 : (^forvar3333)) : ((^reg3343) ?
                  (-reg3334) : "1hbe6p32zpqek5zwx7GxS")) + reg3371) ?
          $signed((reg3246[(1'h0):(1'h0)] != ($unsigned((7'h44)) * $unsigned(forvar3277)))) : $unsigned((((reg3213 ?
                      (8'hbb) : forvar3244) ?
                  $signed(reg3331) : {reg3292, reg3271}) ?
              ((reg3278 ? reg3239 : reg3239) ?
                  (forvar3244 ?
                      reg3381 : reg3215) : (|reg3215)) : (&$unsigned(reg3314)))));
      reg3385 <= "4Us";
      reg3386 <= {(~&reg3270[(5'h10):(3'h6)]), (+$unsigned("qvyaHZfehJRD9Aa"))};
    end
  always
    @(posedge clk) begin
      reg3387 = reg3316[(2'h3):(2'h3)];
      reg3388 = ((~^reg3386[(2'h2):(1'h0)]) != reg3385);
      reg3389 = reg3251;
      reg3390 <= reg3257[(5'h13):(1'h0)];
      for (forvar3391 = (1'h0); (forvar3391 < (3'h4)); forvar3391 = (forvar3391 + (1'h1)))
        begin
          reg3392 <= $signed(((~|reg3267) ?
              reg3367 : (forvar3237[(5'h14):(4'h9)] ?
                  ($signed(wire3207) ?
                      (forvar3269 ? reg3210 : reg3330) : wire3308) : "")));
          reg3393 <= $signed($signed($signed(forvar3223)));
          reg3394 <= reg3266[(3'h7):(2'h3)];
        end
      reg3395 <= reg3328;
    end
  assign wire3396 = (((~|$signed($signed(forvar3295))) < $unsigned(wire3205[(5'h16):(3'h6)])) ?
                        ($signed($signed((reg3224 ?
                            reg3307 : forvar3244))) ^~ reg3224) : ($unsigned(((forvar3297 | reg3342) ?
                            ((8'h9d) ^~ reg3265) : forvar3285[(2'h3):(2'h2)])) <= (($unsigned(reg3344) ?
                                (!(8'ha1)) : $unsigned(forvar3347)) ?
                            ((reg3341 & reg3283) << reg3378) : reg3375)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3068
#( parameter param3200 = (!(((~&((8'hb5) - (8'h9f))) | ({(7'h4d)} ? (^(7'h47)) : ((8'h9c) <= (8'hb1)))) == {(((8'ha3) ? (8'h9c) : (8'hac)) ? ((8'h9d) || (7'h4c)) : ((8'hbc) <= (8'hb7)))}))
, parameter param3201 = {((7'h49) ? param3200 : (~param3200))} )
(y, clk, wire3072, wire3071, wire3070, wire3069);
  output wire [(32'h77d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire3072;
  input wire [(5'h16):(1'h0)] wire3071;
  input wire [(5'h16):(1'h0)] wire3070;
  input wire signed [(4'hd):(1'h0)] wire3069;
  wire signed [(5'h12):(1'h0)] wire3199;
  wire signed [(2'h2):(1'h0)] wire3198;
  wire signed [(5'h12):(1'h0)] wire3197;
  wire [(5'h19):(1'h0)] wire3196;
  reg signed [(5'h11):(1'h0)] reg3195 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3194 = (1'h0);
  reg [(5'h16):(1'h0)] reg3193 = (1'h0);
  reg [(4'h9):(1'h0)] reg3192 = (1'h0);
  reg [(5'h15):(1'h0)] reg3191 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3190 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar3186 = (1'h0);
  reg [(4'hc):(1'h0)] reg3183 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3189 = (1'h0);
  reg [(5'h14):(1'h0)] reg3188 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3187 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3186 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3185 = (1'h0);
  reg [(5'h13):(1'h0)] reg3184 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar3183 = (1'h0);
  reg [(2'h3):(1'h0)] reg3182 = (1'h0);
  reg [(5'h18):(1'h0)] reg3181 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3180 = (1'h0);
  reg [(4'hc):(1'h0)] reg3179 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3178 = (1'h0);
  reg [(2'h2):(1'h0)] reg3177 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3176 = (1'h0);
  reg [(4'he):(1'h0)] reg3175 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3174 = (1'h0);
  reg [(5'h19):(1'h0)] forvar3173 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3172 = (1'h0);
  reg [(3'h6):(1'h0)] reg3171 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3170 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3169 = (1'h0);
  wire signed [(5'h19):(1'h0)] wire3168;
  reg signed [(5'h13):(1'h0)] reg3167 = (1'h0);
  reg [(5'h19):(1'h0)] reg3166 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3165 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3164 = (1'h0);
  reg [(4'h9):(1'h0)] reg3163 = (1'h0);
  reg [(3'h6):(1'h0)] reg3150 = (1'h0);
  reg [(3'h6):(1'h0)] reg3162 = (1'h0);
  reg [(3'h6):(1'h0)] reg3161 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3160 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3159 = (1'h0);
  reg [(2'h3):(1'h0)] reg3158 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3157 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3156 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3155 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3154 = (1'h0);
  reg [(5'h14):(1'h0)] reg3153 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3152 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3151 = (1'h0);
  reg [(5'h15):(1'h0)] forvar3150 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3149 = (1'h0);
  reg [(4'h9):(1'h0)] reg3148 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3147 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire3146;
  wire signed [(5'h11):(1'h0)] wire3145;
  wire signed [(5'h16):(1'h0)] wire3144;
  reg signed [(5'h18):(1'h0)] reg3143 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3142 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3141 = (1'h0);
  reg [(4'hb):(1'h0)] reg3140 = (1'h0);
  reg [(2'h2):(1'h0)] reg3139 = (1'h0);
  reg [(5'h10):(1'h0)] reg3138 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3137 = (1'h0);
  reg [(2'h2):(1'h0)] reg3136 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3135 = (1'h0);
  reg [(5'h15):(1'h0)] reg3134 = (1'h0);
  reg [(4'hc):(1'h0)] reg3133 = (1'h0);
  reg [(4'he):(1'h0)] reg3132 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3131 = (1'h0);
  reg [(5'h17):(1'h0)] reg3130 = (1'h0);
  reg [(2'h3):(1'h0)] reg3129 = (1'h0);
  wire [(4'ha):(1'h0)] wire3128;
  reg [(5'h17):(1'h0)] reg3127 = (1'h0);
  reg [(4'h9):(1'h0)] reg3126 = (1'h0);
  reg [(4'ha):(1'h0)] reg3125 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3124 = (1'h0);
  reg [(5'h12):(1'h0)] forvar3123 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3122 = (1'h0);
  wire signed [(5'h1a):(1'h0)] wire3121;
  reg signed [(3'h6):(1'h0)] reg3120 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3119 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3118 = (1'h0);
  reg [(4'h9):(1'h0)] reg3117 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3116 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar3115 = (1'h0);
  reg [(3'h6):(1'h0)] reg3114 = (1'h0);
  reg [(3'h7):(1'h0)] reg3113 = (1'h0);
  reg [(2'h3):(1'h0)] reg3112 = (1'h0);
  reg [(3'h4):(1'h0)] reg3111 = (1'h0);
  reg [(3'h4):(1'h0)] reg3110 = (1'h0);
  reg [(3'h5):(1'h0)] reg3109 = (1'h0);
  reg [(5'h16):(1'h0)] reg3108 = (1'h0);
  reg [(5'h17):(1'h0)] reg3107 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3106 = (1'h0);
  reg [(5'h13):(1'h0)] reg3105 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3104 = (1'h0);
  reg [(5'h17):(1'h0)] reg3103 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3102 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3101 = (1'h0);
  reg [(5'h10):(1'h0)] reg3100 = (1'h0);
  reg [(5'h16):(1'h0)] reg3099 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3098 = (1'h0);
  reg [(5'h11):(1'h0)] forvar3097 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3096 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3095 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3094 = (1'h0);
  reg [(4'hc):(1'h0)] reg3093 = (1'h0);
  reg [(5'h18):(1'h0)] reg3092 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3091 = (1'h0);
  reg [(5'h14):(1'h0)] reg3090 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3089 = (1'h0);
  reg [(5'h15):(1'h0)] reg3088 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3087 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3086 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3085 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3084 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3083 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3082 = (1'h0);
  reg [(5'h18):(1'h0)] reg3081 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3080 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3079 = (1'h0);
  reg [(5'h19):(1'h0)] forvar3078 = (1'h0);
  wire [(5'h1a):(1'h0)] wire3077;
  wire [(5'h15):(1'h0)] wire3076;
  reg signed [(5'h19):(1'h0)] reg3075 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3074 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3073 = (1'h0);
  assign y = {wire3199,
                 wire3198,
                 wire3197,
                 wire3196,
                 reg3195,
                 reg3194,
                 reg3193,
                 reg3192,
                 reg3191,
                 reg3190,
                 forvar3186,
                 reg3183,
                 reg3189,
                 reg3188,
                 reg3187,
                 reg3186,
                 reg3185,
                 reg3184,
                 forvar3183,
                 reg3182,
                 reg3181,
                 forvar3180,
                 reg3179,
                 reg3178,
                 reg3177,
                 reg3176,
                 reg3175,
                 forvar3174,
                 forvar3173,
                 forvar3172,
                 reg3171,
                 reg3170,
                 forvar3169,
                 wire3168,
                 reg3167,
                 reg3166,
                 reg3165,
                 forvar3164,
                 reg3163,
                 reg3150,
                 reg3162,
                 reg3161,
                 reg3160,
                 reg3159,
                 reg3158,
                 reg3157,
                 reg3156,
                 reg3155,
                 reg3154,
                 reg3153,
                 reg3152,
                 forvar3151,
                 forvar3150,
                 reg3149,
                 reg3148,
                 reg3147,
                 wire3146,
                 wire3145,
                 wire3144,
                 reg3143,
                 reg3142,
                 reg3141,
                 reg3140,
                 reg3139,
                 reg3138,
                 forvar3137,
                 reg3136,
                 forvar3135,
                 reg3134,
                 reg3133,
                 reg3132,
                 reg3131,
                 reg3130,
                 reg3129,
                 wire3128,
                 reg3127,
                 reg3126,
                 reg3125,
                 reg3124,
                 forvar3123,
                 reg3122,
                 wire3121,
                 reg3120,
                 reg3119,
                 reg3118,
                 reg3117,
                 reg3116,
                 forvar3115,
                 reg3114,
                 reg3113,
                 reg3112,
                 reg3111,
                 reg3110,
                 reg3109,
                 reg3108,
                 reg3107,
                 reg3106,
                 reg3105,
                 reg3104,
                 reg3103,
                 reg3102,
                 forvar3101,
                 reg3100,
                 reg3099,
                 reg3098,
                 forvar3097,
                 reg3096,
                 reg3095,
                 forvar3094,
                 reg3093,
                 reg3092,
                 reg3091,
                 reg3090,
                 reg3089,
                 reg3088,
                 reg3087,
                 forvar3086,
                 reg3085,
                 reg3084,
                 reg3083,
                 reg3082,
                 reg3081,
                 reg3080,
                 reg3079,
                 forvar3078,
                 wire3077,
                 wire3076,
                 reg3075,
                 reg3074,
                 reg3073,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg3073 <= (wire3071[(2'h3):(1'h0)] << $signed($unsigned(wire3069)));
      reg3074 <= ("84GYUKg0zMlcWnmewa" | ((-((-reg3073) & "zcLkY")) != (wire3070[(5'h14):(4'hb)] ^ wire3071)));
      reg3075 <= ("KtKih2OC" ? (7'h4b) : wire3070[(4'he):(3'h4)]);
    end
  assign wire3076 = $signed((^~(8'ha8)));
  assign wire3077 = $signed((wire3076 ?
                        (reg3073[(1'h0):(1'h0)] ?
                            ((^~reg3074) < (+wire3069)) : reg3075[(5'h15):(4'ha)]) : reg3074));
  always
    @(posedge clk) begin
      for (forvar3078 = (1'h0); (forvar3078 < (3'h5)); forvar3078 = (forvar3078 + (1'h1)))
        begin
          reg3079 <= "";
          reg3080 <= $unsigned((^~(|"f")));
          reg3081 <= wire3076;
        end
      reg3082 = wire3077;
      reg3083 = ((($signed(reg3073[(1'h1):(1'h1)]) ?
          reg3081 : "zgFYZnro7g3VVz6UCpyC4K") - $signed($unsigned($unsigned(wire3071)))) != "BRo3C8cdQlI3veoOQW");
      reg3084 <= $signed($signed((reg3073 ?
          {(^reg3083)} : {reg3080, (^wire3071)})));
      if ((("Ma0yZAvsBOSLSNLVC7w" ?
          reg3083[(2'h2):(2'h2)] : (~&("v5n" ?
              $unsigned(reg3081) : (reg3079 ?
                  (8'hba) : (8'hb8))))) - (~^$unsigned("lGLM"))))
        begin
          reg3085 <= (&reg3079);
          for (forvar3086 = (1'h0); (forvar3086 < (2'h3)); forvar3086 = (forvar3086 + (1'h1)))
            begin
              reg3087 <= forvar3086;
            end
          reg3088 <= forvar3086;
          reg3089 <= reg3079;
          reg3090 <= {(8'ha0)};
        end
      else
        begin
          reg3085 <= reg3087[(1'h0):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      reg3091 <= forvar3078[(5'h16):(4'h9)];
      reg3092 <= $signed((~^(+$signed($unsigned(forvar3078)))));
      reg3093 <= wire3069;
      for (forvar3094 = (1'h0); (forvar3094 < (1'h1)); forvar3094 = (forvar3094 + (1'h1)))
        begin
          reg3095 <= wire3070;
        end
    end
  always
    @(posedge clk) begin
      reg3096 <= ($signed($signed(reg3080)) - {(+reg3093[(1'h0):(1'h0)])});
      for (forvar3097 = (1'h0); (forvar3097 < (2'h2)); forvar3097 = (forvar3097 + (1'h1)))
        begin
          reg3098 <= ((~|"") ?
              wire3076[(1'h1):(1'h1)] : ($unsigned(reg3090[(3'h6):(1'h1)]) > ($unsigned(reg3079) ?
                  $unsigned((wire3077 ? reg3087 : reg3083)) : reg3095)));
          reg3099 = $unsigned(($unsigned(reg3088) ?
              {((wire3077 == wire3069) ?
                      "C9Gpv4S1bwiuNlqaG" : "8JNKAwYLKXdC9Qma1p6BqLg")} : (&$unsigned((reg3081 <= wire3076)))));
          reg3100 <= $signed("rmZYyAukS4W4EAYBRcIA9Ep");
          for (forvar3101 = (1'h0); (forvar3101 < (3'h5)); forvar3101 = (forvar3101 + (1'h1)))
            begin
              reg3102 <= "ORlHPnhOuRzztFq0Y0RIto0v";
              reg3103 <= $unsigned($signed(reg3089[(3'h7):(1'h1)]));
              reg3104 <= $unsigned(($unsigned($signed((wire3076 >= reg3092))) ?
                  reg3096[(2'h2):(1'h0)] : reg3091));
            end
          reg3105 = (forvar3094[(1'h1):(1'h1)] ?
              ({{$signed(reg3075), {reg3103, reg3089}},
                  (|(reg3088 ? reg3080 : wire3076))} + (("4OYKzMopinui6fKo" ?
                  reg3074 : {reg3073,
                      reg3102}) * (~$signed(reg3102)))) : {(~&$signed("FWk5zaInm"))});
        end
    end
  always
    @(posedge clk) begin
      reg3106 = $unsigned("U");
      reg3107 = forvar3101[(4'hd):(3'h6)];
      if ($unsigned((~&$unsigned({(8'hb4)}))))
        begin
          reg3108 <= ("eu" ? ((7'h4a) && {(7'h48), "KegAe1Bmc"}) : reg3083);
        end
      else
        begin
          reg3108 <= forvar3094[(2'h2):(2'h2)];
          reg3109 <= $unsigned("Yh");
          reg3110 <= (reg3098[(3'h7):(3'h6)] >> reg3085);
          reg3111 <= (|("dmbaHsUZnJu3t7r" ?
              {(~^{reg3079, reg3093}),
                  ((reg3074 >>> reg3100) ?
                      (reg3087 || reg3079) : {reg3104,
                          reg3079})} : (((|forvar3094) <<< (~(8'hb2))) + (7'h45))));
          reg3112 <= $unsigned(((~$unsigned($signed(wire3072))) ?
              forvar3086[(2'h2):(2'h2)] : $signed($unsigned("G6T7ExRRRZ649Unw"))));
          reg3113 <= "JuYHnCC8yLAgJghZh1";
        end
    end
  always
    @(posedge clk) begin
      reg3114 <= $signed((reg3103[(4'hf):(2'h3)] != $unsigned(({reg3081} ?
          (reg3080 ? reg3107 : reg3111) : {wire3077}))));
      for (forvar3115 = (1'h0); (forvar3115 < (3'h4)); forvar3115 = (forvar3115 + (1'h1)))
        begin
          reg3116 <= (reg3084 ?
              (|($signed(wire3070) & ((-wire3071) << reg3073[(1'h1):(1'h1)]))) : (-forvar3078[(4'ha):(4'h9)]));
          reg3117 <= (^~(~(reg3112[(2'h3):(1'h0)] ?
              (-(forvar3094 ? reg3106 : (7'h46))) : {(!reg3102)})));
          reg3118 <= (((wire3071 ?
              ((^~reg3099) + reg3089) : (+$unsigned(forvar3078))) ^ (+((+reg3112) ?
              (reg3099 ? reg3073 : reg3096) : (reg3089 ?
                  wire3077 : reg3109)))) <= reg3113[(3'h5):(3'h5)]);
          reg3119 = $unsigned(($signed(("odLbAgFu3dg" >>> (~|reg3106))) ?
              $signed(reg3088) : ($signed((reg3091 ? reg3105 : (8'ha9))) ?
                  $signed(wire3072) : reg3092)));
        end
      reg3120 <= "g7nMwhRK6hHQEHIS";
    end
  assign wire3121 = $signed(reg3075[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg3122 <= (~&"72ykT");
      for (forvar3123 = (1'h0); (forvar3123 < (2'h2)); forvar3123 = (forvar3123 + (1'h1)))
        begin
          reg3124 <= {reg3098};
          reg3125 <= (|reg3109[(3'h4):(2'h3)]);
          reg3126 <= reg3093;
        end
      reg3127 = reg3079;
    end
  assign wire3128 = (~reg3108[(3'h7):(3'h5)]);
  always
    @(posedge clk) begin
      reg3129 <= reg3112[(1'h1):(1'h1)];
      reg3130 <= "AU46YN";
      reg3131 <= $unsigned(reg3108[(3'h5):(1'h0)]);
      reg3132 <= (^(forvar3101 < $unsigned(forvar3078[(5'h11):(5'h10)])));
      reg3133 = (("Z5YrDhJ" <<< $signed(((reg3124 ? reg3095 : (8'hb4)) ?
          (reg3093 ? (8'h9e) : wire3121) : (reg3088 ?
              wire3076 : reg3098)))) & reg3118);
    end
  always
    @(posedge clk) begin
      reg3134 <= (~&$unsigned(({(reg3082 ? wire3121 : reg3118),
          reg3131} != (~^reg3091))));
      for (forvar3135 = (1'h0); (forvar3135 < (1'h0)); forvar3135 = (forvar3135 + (1'h1)))
        begin
          reg3136 <= (8'ha4);
          for (forvar3137 = (1'h0); (forvar3137 < (3'h4)); forvar3137 = (forvar3137 + (1'h1)))
            begin
              reg3138 <= "51UbW";
              reg3139 <= $signed($unsigned($signed($unsigned($signed((7'h42))))));
              reg3140 = (^~"");
              reg3141 <= reg3132;
            end
          reg3142 <= $signed(reg3083[(2'h3):(2'h2)]);
          reg3143 <= reg3089[(4'he):(4'ha)];
        end
    end
  assign wire3144 = {((forvar3123 + reg3083[(2'h3):(1'h0)]) ?
                            reg3130 : reg3118),
                        forvar3101};
  assign wire3145 = $unsigned({$signed(((~^(8'ha0)) ?
                            $unsigned(reg3092) : "mbiDepoZFJ2sGOFvClz"))});
  assign wire3146 = (reg3131 < $signed("TdKyfy0"));
  always
    @(posedge clk) begin
      reg3147 <= wire3077[(4'hc):(2'h2)];
      reg3148 = (wire3128[(1'h1):(1'h1)] ?
          (8'ha8) : ({reg3129[(2'h3):(1'h0)],
                  ((wire3145 >= reg3098) * $unsigned(forvar3115))} ?
              wire3069[(4'hd):(4'hb)] : "nxtRHWiQ0hnocy9kTm"));
      if (reg3133[(3'h5):(2'h2)])
        begin
          reg3149 <= ($signed(((reg3100[(4'h9):(1'h0)] + reg3106[(1'h0):(1'h0)]) ^~ $unsigned(forvar3123))) ^ "7iN");
          for (forvar3150 = (1'h0); (forvar3150 < (3'h4)); forvar3150 = (forvar3150 + (1'h1)))
            begin
              for (forvar3151 = (1'h0); (forvar3151 < (1'h1)); forvar3151 = (forvar3151 + (1'h1)))
                begin
                  reg3152 <= "CCNgWqmH47iL";
                  reg3153 <= wire3076[(5'h10):(4'hb)];
                  reg3154 <= reg3119[(3'h7):(2'h3)];
                  reg3155 = $signed((("OwRegHIkt9hFx084acU" ?
                      "CZZyYkLwpoJy3ivMV49WYWv" : {((8'h9e) - reg3129)}) < (-("aF0ZSG" ?
                      $unsigned((7'h41)) : wire3072))));
                  reg3156 <= forvar3151[(1'h0):(1'h0)];
                end
              reg3157 <= forvar3135[(2'h3):(1'h1)];
              reg3158 <= ((!(8'hba)) * ($unsigned((~(~^reg3083))) ?
                  $signed({(reg3119 ?
                          reg3107 : reg3099)}) : forvar3086[(2'h3):(1'h0)]));
              reg3159 <= reg3140[(4'h9):(3'h4)];
            end
          reg3160 <= reg3155[(4'he):(4'h9)];
          reg3161 = ($signed((^~(8'h9e))) ~^ {(8'ha1)});
          reg3162 <= $unsigned(((reg3131[(4'h9):(3'h7)] > forvar3086) ?
              ("PZcxsElPFYB" ?
                  (~(8'ha0)) : reg3085[(2'h2):(2'h2)]) : (^~(&(forvar3135 ^ wire3069)))));
        end
      else
        begin
          reg3149 <= "vDXiIZuGUP848T0mlC9DM";
          reg3150 <= ($signed("SeNHKMMnMun7JRl") < $unsigned(wire3072));
          for (forvar3151 = (1'h0); (forvar3151 < (3'h5)); forvar3151 = (forvar3151 + (1'h1)))
            begin
              reg3152 <= "UfX79OGx3fwoyLBBMgAeHEW";
              reg3153 = (8'hb7);
              reg3154 <= {($unsigned($unsigned($unsigned(forvar3101))) ?
                      $signed(($unsigned(reg3143) ?
                          $signed(reg3104) : (reg3105 > forvar3150))) : "Rh"),
                  "4nwxNIXnate3BGO7SwhvC6"};
            end
          reg3155 <= ("AzQA3muH6nTOiIXV" ?
              ($signed(((forvar3115 & reg3088) ?
                  (^wire3145) : $signed(reg3114))) >= ((reg3134[(5'h13):(4'h8)] ?
                  reg3075 : $unsigned(reg3162)) && (!"iuKr5rnUXd06n"))) : (reg3161[(1'h0):(1'h0)] ^~ ("DxpqGv6tUW4N10" ?
                  "PH" : reg3129)));
        end
    end
  always
    @(posedge clk) begin
      reg3163 <= "mQJVio8ns";
      for (forvar3164 = (1'h0); (forvar3164 < (2'h3)); forvar3164 = (forvar3164 + (1'h1)))
        begin
          reg3165 <= $signed($unsigned((8'ha7)));
          reg3166 = forvar3078;
          reg3167 = ($signed($signed($unsigned(reg3133))) ~^ (reg3093[(2'h3):(1'h1)] ^ (wire3076[(3'h7):(3'h6)] || ((8'ha3) ^ reg3119[(4'hd):(3'h5)]))));
        end
    end
  assign wire3168 = (8'h9e);
  always
    @(posedge clk) begin
      for (forvar3169 = (1'h0); (forvar3169 < (2'h2)); forvar3169 = (forvar3169 + (1'h1)))
        begin
          reg3170 <= (&$unsigned(reg3153[(3'h4):(2'h3)]));
        end
      reg3171 <= forvar3150;
      for (forvar3172 = (1'h0); (forvar3172 < (2'h3)); forvar3172 = (forvar3172 + (1'h1)))
        begin
          for (forvar3173 = (1'h0); (forvar3173 < (2'h2)); forvar3173 = (forvar3173 + (1'h1)))
            begin
              for (forvar3174 = (1'h0); (forvar3174 < (2'h2)); forvar3174 = (forvar3174 + (1'h1)))
                begin
                  reg3175 <= $unsigned(((forvar3137 ?
                          $signed("fCxzBeK9Fb5OMGWKWl1B45yBB") : {$signed(reg3171),
                              (~reg3074)}) ?
                      reg3091 : forvar3123[(1'h0):(1'h0)]));
                  reg3176 <= reg3160[(2'h3):(2'h3)];
                end
              reg3177 = $signed("EmWC6ycSqJFEBcn");
              reg3178 <= ($unsigned($unsigned({(~&reg3110)})) ?
                  $unsigned(reg3153) : {reg3170[(2'h3):(1'h0)],
                      (("" >>> ((8'hbd) ? reg3120 : reg3170)) ?
                          (~reg3083[(2'h3):(1'h1)]) : ({reg3073} ?
                              {reg3165} : (~&reg3161)))});
              reg3179 <= ((~&reg3103[(5'h14):(3'h6)]) != {(~&$signed({reg3167,
                      wire3076})),
                  (^~{"wB"})});
              for (forvar3180 = (1'h0); (forvar3180 < (2'h3)); forvar3180 = (forvar3180 + (1'h1)))
                begin
                  reg3181 = $unsigned(reg3074[(3'h4):(1'h1)]);
                  reg3182 <= (~^($unsigned((8'h9e)) ?
                      (($signed(reg3122) ?
                          reg3139 : $signed(forvar3094)) >= "PKE5qTBPos1oCTLIJLCubGTIb") : reg3124));
                end
            end
          if (reg3110[(1'h1):(1'h0)])
            begin
              for (forvar3183 = (1'h0); (forvar3183 < (2'h2)); forvar3183 = (forvar3183 + (1'h1)))
                begin
                  reg3184 <= {$unsigned(reg3153[(5'h10):(4'hd)]), "I729X32"};
                  reg3185 <= wire3071;
                  reg3186 = reg3159;
                  reg3187 <= ($unsigned("ayChG6C0xyz") + "");
                  reg3188 <= (reg3150[(2'h2):(1'h0)] ? "7catv1G" : reg3175);
                  reg3189 = reg3141[(4'hd):(3'h4)];
                end
            end
          else
            begin
              reg3183 <= reg3141[(5'h16):(3'h7)];
              reg3184 <= {("X" ?
                      "sgWs4Ped4Rh8JkJXfLw" : $unsigned(wire3077[(1'h0):(1'h0)]))};
              reg3185 = reg3132[(4'hc):(2'h2)];
              for (forvar3186 = (1'h0); (forvar3186 < (3'h4)); forvar3186 = (forvar3186 + (1'h1)))
                begin
                  reg3187 <= $unsigned(((8'ha1) < $unsigned($unsigned((reg3161 ?
                      (8'hb4) : reg3100)))));
                  reg3188 <= (^~$unsigned($unsigned("yNuIgdgu")));
                  reg3189 <= $unsigned(forvar3101);
                  reg3190 = "x2kteOCHvxcRv5zDy9c";
                end
              reg3191 <= (reg3127 ?
                  {reg3095,
                      $unsigned("TlckPbD")} : "xAWX8Kalapt59WUZwWyiT0GH6");
              reg3192 <= reg3091[(3'h4):(1'h0)];
            end
          reg3193 = wire3128[(4'ha):(3'h4)];
        end
      reg3194 = {$signed($signed((!{(8'hb1)})))};
      reg3195 <= reg3127;
    end
  assign wire3196 = "f2NUD";
  assign wire3197 = $signed(("nL0gA0yQSV" + (((|reg3183) ?
                        (forvar3123 >= wire3168) : (+reg3120)) ^ ((reg3147 ?
                        wire3146 : reg3108) >>> (reg3098 ?
                        forvar3186 : (7'h49))))));
  assign wire3198 = "DnTflYJzwQ7uw8n1z7lWrK";
  assign wire3199 = $unsigned("f52PT2w9S9RpcxF");
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3018  (y, clk, wire3023, wire3022, wire3021, wire3020, wire3019);
  output wire [(32'h22f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire3023;
  input wire signed [(3'h4):(1'h0)] wire3022;
  input wire [(5'h17):(1'h0)] wire3021;
  input wire [(5'h14):(1'h0)] wire3020;
  input wire signed [(4'he):(1'h0)] wire3019;
  wire signed [(3'h4):(1'h0)] wire3065;
  reg signed [(4'ha):(1'h0)] reg3064 = (1'h0);
  reg [(4'ha):(1'h0)] reg3063 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3062 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3061 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3060 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3059 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3058 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3057 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3056 = (1'h0);
  reg [(4'h8):(1'h0)] reg3055 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3054 = (1'h0);
  reg [(4'h9):(1'h0)] reg3053 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3052 = (1'h0);
  reg [(4'hf):(1'h0)] reg3051 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3050 = (1'h0);
  reg [(5'h14):(1'h0)] reg3049 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar3048 = (1'h0);
  wire signed [(5'h19):(1'h0)] wire3047;
  reg signed [(3'h5):(1'h0)] reg3046 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3045 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire3044;
  reg [(3'h5):(1'h0)] reg3043 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3042 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3041 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3040 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3039 = (1'h0);
  reg [(4'he):(1'h0)] reg3038 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3037 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3036 = (1'h0);
  reg [(4'hb):(1'h0)] reg3035 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3034 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3033 = (1'h0);
  reg [(4'hd):(1'h0)] reg3032 = (1'h0);
  reg [(4'h9):(1'h0)] reg3031 = (1'h0);
  reg [(4'hb):(1'h0)] reg3030 = (1'h0);
  reg [(4'ha):(1'h0)] reg3029 = (1'h0);
  reg [(4'hd):(1'h0)] reg3028 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3027 = (1'h0);
  reg [(4'hd):(1'h0)] reg3026 = (1'h0);
  wire [(3'h4):(1'h0)] wire3025;
  wire [(5'h1a):(1'h0)] wire3024;
  assign y = {wire3065,
                 reg3064,
                 reg3063,
                 reg3062,
                 reg3061,
                 reg3060,
                 reg3059,
                 reg3058,
                 reg3057,
                 forvar3056,
                 reg3055,
                 reg3054,
                 reg3053,
                 reg3052,
                 reg3051,
                 forvar3050,
                 reg3049,
                 forvar3048,
                 wire3047,
                 reg3046,
                 reg3045,
                 wire3044,
                 reg3043,
                 reg3042,
                 reg3041,
                 reg3040,
                 forvar3039,
                 reg3038,
                 reg3037,
                 reg3036,
                 reg3035,
                 reg3034,
                 reg3033,
                 reg3032,
                 reg3031,
                 reg3030,
                 reg3029,
                 reg3028,
                 reg3027,
                 reg3026,
                 wire3025,
                 wire3024,
                 (1'h0)};
  assign wire3024 = (&{wire3019[(4'hb):(1'h0)],
                        ($unsigned((wire3021 ?
                            wire3020 : wire3021)) - (~^$signed(wire3021)))});
  assign wire3025 = ((((-wire3022) || wire3019[(4'hc):(3'h4)]) | ((|(~|wire3024)) >> ((~wire3020) & wire3021))) && $unsigned(((+wire3024) ?
                        ((wire3024 < (7'h45)) ?
                            $signed(wire3022) : (wire3023 ?
                                wire3019 : wire3019)) : (wire3020 * (wire3023 ?
                            wire3020 : wire3023)))));
  always
    @(posedge clk) begin
      reg3026 <= ("sKNyb1H" ~^ ((wire3022 ?
              (((8'h9d) != wire3023) ?
                  (!wire3023) : (~^(8'haa))) : ($signed((8'hbe)) ~^ wire3024)) ?
          "GwWpxBuSyNTxAU8b2XqnLPb" : "OkzBo7e7K"));
      reg3027 = (+wire3023);
      reg3028 <= wire3024;
      reg3029 = $unsigned(wire3020);
      reg3030 = wire3019[(4'hb):(1'h1)];
      reg3031 <= (8'hab);
    end
  always
    @(posedge clk) begin
      reg3032 <= $unsigned((-wire3022));
      reg3033 <= $signed({$unsigned((~|$unsigned(wire3025)))});
    end
  always
    @(posedge clk) begin
      reg3034 <= $unsigned(wire3025);
      reg3035 <= $unsigned("zg1SG1");
      reg3036 <= ((~^wire3019) ?
          "M4Rx4AzLsN2VJ6Mvm" : ({{(wire3023 ^~ reg3028)},
              wire3021[(3'h5):(2'h2)]} - (~&"HqP")));
    end
  always
    @(posedge clk) begin
      reg3037 <= ((-(+$unsigned("sZTyOSh6OQ"))) ~^ {$signed((-(reg3030 + wire3019)))});
      reg3038 <= {{"GksGWnFWY",
              ((!wire3025[(3'h4):(2'h3)]) ?
                  wire3021[(4'hf):(3'h5)] : (^~wire3023[(4'hf):(4'ha)]))},
          {(reg3033[(5'h14):(4'h9)] ?
                  $unsigned(((8'hb3) == reg3034)) : wire3023),
              ($unsigned($unsigned(reg3032)) ~^ ((reg3037 > wire3021) ?
                  $signed(wire3022) : $signed(reg3037)))}};
      for (forvar3039 = (1'h0); (forvar3039 < (3'h5)); forvar3039 = (forvar3039 + (1'h1)))
        begin
          reg3040 <= ({reg3033} * wire3019[(4'h8):(1'h1)]);
        end
      reg3041 = ($unsigned(forvar3039) == "3vZqIhGf43uCSCfWAoH");
      reg3042 = {forvar3039,
          $unsigned((("w" ?
                  (wire3025 ? reg3030 : reg3027) : (reg3037 - (8'ha6))) ?
              $signed((reg3040 >>> reg3030)) : $unsigned(reg3036)))};
      reg3043 <= (~^reg3036[(3'h4):(3'h4)]);
    end
  assign wire3044 = (~$signed({reg3034[(2'h2):(2'h2)]}));
  always
    @(posedge clk) begin
      reg3045 <= $unsigned((((&(^reg3032)) ?
          (~$unsigned(reg3032)) : (~&(~&reg3036))) - (-wire3021[(1'h1):(1'h1)])));
      reg3046 <= $signed($signed($signed((8'hba))));
    end
  assign wire3047 = ((^(|$signed({(8'ha2),
                        reg3041}))) << {(~&reg3030[(4'ha):(1'h1)])});
  always
    @(posedge clk) begin
      for (forvar3048 = (1'h0); (forvar3048 < (3'h4)); forvar3048 = (forvar3048 + (1'h1)))
        begin
          reg3049 <= $unsigned(forvar3048[(1'h0):(1'h0)]);
        end
      for (forvar3050 = (1'h0); (forvar3050 < (3'h4)); forvar3050 = (forvar3050 + (1'h1)))
        begin
          reg3051 <= "qfNJkyyYAKhJewfRVaEs";
          reg3052 = reg3051;
          reg3053 <= (reg3043 ?
              ((~(reg3043[(3'h4):(1'h0)] ?
                  $unsigned(reg3049) : reg3042)) || (($unsigned(reg3029) ?
                  $unsigned((7'h42)) : reg3034) <= reg3049)) : $unsigned($signed($signed((reg3051 ?
                  reg3027 : reg3029)))));
          reg3054 <= $signed({$signed($signed($signed(wire3021))),
              reg3026[(3'h4):(1'h0)]});
          reg3055 <= ((wire3024 - reg3038[(4'ha):(4'h8)]) - $signed((-wire3023[(4'hd):(4'hd)])));
          for (forvar3056 = (1'h0); (forvar3056 < (3'h4)); forvar3056 = (forvar3056 + (1'h1)))
            begin
              reg3057 <= reg3046[(1'h0):(1'h0)];
              reg3058 <= {reg3026,
                  {(~|$signed((&reg3029))),
                      (reg3030[(4'h9):(4'h9)] >= $unsigned(wire3021))}};
              reg3059 <= reg3051[(3'h6):(1'h0)];
              reg3060 <= $unsigned("y2eey2xQmcJlW7B");
              reg3061 <= reg3034;
              reg3062 <= {$signed($unsigned({$signed((7'h46))}))};
            end
        end
      reg3063 <= $unsigned(reg3028[(4'hd):(3'h5)]);
      reg3064 <= ("wbwV2" - ($signed(wire3047[(5'h13):(4'hf)]) * $signed(($signed(reg3052) != ((8'ha8) ?
          reg3053 : (8'ha7))))));
    end
  assign wire3065 = (~$signed(wire3023));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2841  (y, clk, wire2846, wire2845, wire2844, wire2843, wire2842);
  output wire [(32'h79b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire2846;
  input wire signed [(4'h8):(1'h0)] wire2845;
  input wire [(5'h16):(1'h0)] wire2844;
  input wire [(5'h1a):(1'h0)] wire2843;
  input wire [(2'h2):(1'h0)] wire2842;
  wire signed [(5'h10):(1'h0)] wire2981;
  reg [(2'h2):(1'h0)] reg2980 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2979 = (1'h0);
  reg [(2'h3):(1'h0)] reg2978 = (1'h0);
  reg [(3'h4):(1'h0)] reg2977 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2976 = (1'h0);
  reg [(5'h12):(1'h0)] reg2975 = (1'h0);
  reg [(4'hc):(1'h0)] reg2974 = (1'h0);
  reg [(5'h13):(1'h0)] reg2973 = (1'h0);
  reg [(4'hf):(1'h0)] reg2972 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2971 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2970 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2969 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2968 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2967 = (1'h0);
  reg [(4'hd):(1'h0)] reg2966 = (1'h0);
  reg [(5'h12):(1'h0)] reg2965 = (1'h0);
  reg [(5'h18):(1'h0)] reg2964 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2963 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2962 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2961 = (1'h0);
  reg [(5'h13):(1'h0)] reg2961 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2960 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2959 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2958 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2957 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2956 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire2955;
  reg signed [(2'h3):(1'h0)] reg2954 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2953 = (1'h0);
  reg [(5'h18):(1'h0)] reg2952 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2951 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2950 = (1'h0);
  reg [(5'h10):(1'h0)] reg2949 = (1'h0);
  reg [(5'h14):(1'h0)] reg2948 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2947 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2946 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2945 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2944 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2943 = (1'h0);
  reg [(4'hc):(1'h0)] reg2942 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2941 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2938 = (1'h0);
  reg [(4'ha):(1'h0)] reg2940 = (1'h0);
  reg [(5'h15):(1'h0)] reg2939 = (1'h0);
  reg [(5'h18):(1'h0)] reg2938 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2937 = (1'h0);
  reg [(5'h14):(1'h0)] reg2936 = (1'h0);
  reg [(4'he):(1'h0)] reg2935 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2934 = (1'h0);
  reg [(2'h2):(1'h0)] reg2933 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2932 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2931 = (1'h0);
  reg [(5'h17):(1'h0)] reg2930 = (1'h0);
  reg [(4'he):(1'h0)] reg2929 = (1'h0);
  reg [(4'ha):(1'h0)] reg2928 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2927 = (1'h0);
  reg [(4'hd):(1'h0)] reg2926 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2925 = (1'h0);
  reg [(5'h19):(1'h0)] reg2924 = (1'h0);
  reg [(4'h8):(1'h0)] reg2923 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar2922 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2921 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2920 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2919 = (1'h0);
  reg [(5'h16):(1'h0)] reg2918 = (1'h0);
  reg [(4'hc):(1'h0)] reg2917 = (1'h0);
  reg [(4'h8):(1'h0)] reg2916 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2915 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2914 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2913 = (1'h0);
  reg [(5'h13):(1'h0)] reg2912 = (1'h0);
  reg [(2'h2):(1'h0)] reg2911 = (1'h0);
  reg [(3'h6):(1'h0)] reg2910 = (1'h0);
  reg [(5'h14):(1'h0)] reg2909 = (1'h0);
  reg [(5'h17):(1'h0)] reg2908 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2907 = (1'h0);
  reg [(4'ha):(1'h0)] reg2906 = (1'h0);
  reg [(3'h5):(1'h0)] reg2905 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2904 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar2902 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2899 = (1'h0);
  reg [(4'h9):(1'h0)] reg2903 = (1'h0);
  reg [(5'h16):(1'h0)] reg2902 = (1'h0);
  reg [(4'hf):(1'h0)] reg2901 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2900 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2899 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2898 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2897 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2896 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2895 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2894 = (1'h0);
  reg [(4'ha):(1'h0)] reg2893 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2892 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2891 = (1'h0);
  wire [(5'h17):(1'h0)] wire2890;
  reg signed [(3'h4):(1'h0)] reg2889 = (1'h0);
  reg [(5'h10):(1'h0)] reg2888 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2887 = (1'h0);
  reg [(2'h3):(1'h0)] reg2886 = (1'h0);
  reg [(4'hf):(1'h0)] reg2885 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2884 = (1'h0);
  reg [(4'h9):(1'h0)] reg2883 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2882 = (1'h0);
  reg [(2'h3):(1'h0)] reg2881 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2880 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2879 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2878 = (1'h0);
  reg [(4'h8):(1'h0)] reg2877 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2876 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2875 = (1'h0);
  reg [(5'h17):(1'h0)] reg2874 = (1'h0);
  reg [(5'h16):(1'h0)] forvar2873 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2872 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2871 = (1'h0);
  reg [(4'h9):(1'h0)] reg2870 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2869 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2868 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2867 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2866 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2865 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2864 = (1'h0);
  reg [(4'ha):(1'h0)] reg2863 = (1'h0);
  reg [(4'hb):(1'h0)] reg2862 = (1'h0);
  reg [(3'h5):(1'h0)] reg2861 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2860 = (1'h0);
  reg [(5'h15):(1'h0)] reg2859 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2858 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2857 = (1'h0);
  reg [(5'h14):(1'h0)] reg2856 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar2855 = (1'h0);
  reg [(3'h5):(1'h0)] reg2854 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2853 = (1'h0);
  reg [(5'h13):(1'h0)] reg2852 = (1'h0);
  reg [(4'hf):(1'h0)] reg2851 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2850 = (1'h0);
  reg [(5'h19):(1'h0)] reg2849 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2848 = (1'h0);
  reg [(2'h2):(1'h0)] reg2847 = (1'h0);
  assign y = {wire2981,
                 reg2980,
                 reg2979,
                 reg2978,
                 reg2977,
                 reg2976,
                 reg2975,
                 reg2974,
                 reg2973,
                 reg2972,
                 forvar2971,
                 forvar2970,
                 reg2969,
                 reg2968,
                 reg2967,
                 reg2966,
                 reg2965,
                 reg2964,
                 reg2963,
                 reg2962,
                 forvar2961,
                 reg2961,
                 reg2960,
                 forvar2959,
                 reg2958,
                 reg2957,
                 reg2956,
                 wire2955,
                 reg2954,
                 reg2953,
                 reg2952,
                 reg2951,
                 reg2950,
                 reg2949,
                 reg2948,
                 forvar2947,
                 reg2946,
                 forvar2945,
                 reg2944,
                 reg2943,
                 reg2942,
                 reg2941,
                 forvar2938,
                 reg2940,
                 reg2939,
                 reg2938,
                 reg2937,
                 reg2936,
                 reg2935,
                 reg2934,
                 reg2933,
                 reg2932,
                 reg2931,
                 reg2930,
                 reg2929,
                 reg2928,
                 reg2927,
                 reg2926,
                 forvar2925,
                 reg2924,
                 reg2923,
                 forvar2922,
                 reg2921,
                 reg2920,
                 reg2919,
                 reg2918,
                 reg2917,
                 reg2916,
                 reg2915,
                 reg2914,
                 reg2913,
                 reg2912,
                 reg2911,
                 reg2910,
                 reg2909,
                 reg2908,
                 forvar2907,
                 reg2906,
                 reg2905,
                 reg2904,
                 forvar2902,
                 forvar2899,
                 reg2903,
                 reg2902,
                 reg2901,
                 reg2900,
                 reg2899,
                 reg2898,
                 reg2897,
                 reg2896,
                 reg2895,
                 forvar2894,
                 reg2893,
                 reg2892,
                 reg2891,
                 wire2890,
                 reg2889,
                 reg2888,
                 reg2887,
                 reg2886,
                 reg2885,
                 forvar2884,
                 reg2883,
                 reg2882,
                 reg2881,
                 forvar2880,
                 reg2879,
                 reg2878,
                 reg2877,
                 reg2876,
                 reg2875,
                 reg2874,
                 forvar2873,
                 reg2872,
                 reg2871,
                 reg2870,
                 forvar2869,
                 forvar2868,
                 reg2867,
                 reg2866,
                 reg2865,
                 reg2864,
                 reg2863,
                 reg2862,
                 reg2861,
                 forvar2860,
                 reg2859,
                 reg2858,
                 reg2857,
                 reg2856,
                 forvar2855,
                 reg2854,
                 forvar2853,
                 reg2852,
                 reg2851,
                 reg2850,
                 reg2849,
                 forvar2848,
                 reg2847,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg2847 <= $unsigned(("OcGODM2nQBlgJI" << $unsigned(($signed(wire2846) >>> wire2843))));
    end
  always
    @(posedge clk) begin
      for (forvar2848 = (1'h0); (forvar2848 < (1'h0)); forvar2848 = (forvar2848 + (1'h1)))
        begin
          reg2849 = forvar2848[(1'h1):(1'h0)];
          reg2850 <= (reg2849[(4'h9):(3'h5)] ?
              $unsigned((($signed(wire2844) * reg2849) ?
                  (8'hb4) : (wire2843 ?
                      {reg2849} : $signed(wire2842)))) : reg2849[(5'h13):(4'hb)]);
          reg2851 <= ($unsigned(forvar2848[(1'h0):(1'h0)]) & $unsigned("xmpU"));
          reg2852 <= (!forvar2848);
        end
      for (forvar2853 = (1'h0); (forvar2853 < (3'h5)); forvar2853 = (forvar2853 + (1'h1)))
        begin
          if ((~^(wire2843 ? "T1HW" : (^$unsigned((wire2843 & reg2850))))))
            begin
              reg2854 <= (~reg2851);
              for (forvar2855 = (1'h0); (forvar2855 < (3'h4)); forvar2855 = (forvar2855 + (1'h1)))
                begin
                  reg2856 <= (^~"9");
                end
            end
          else
            begin
              reg2854 = "uFBCJ";
            end
          reg2857 <= $signed($signed("U0OJXuu5983XM"));
          reg2858 <= $signed(reg2847);
          reg2859 <= reg2849;
          for (forvar2860 = (1'h0); (forvar2860 < (2'h2)); forvar2860 = (forvar2860 + (1'h1)))
            begin
              reg2861 = "vuT07H3m49bIQLPvw";
              reg2862 <= $signed($signed($signed((((7'h4d) ?
                      wire2843 : reg2847) ?
                  wire2842 : $unsigned(reg2850)))));
              reg2863 <= ($signed(((!$unsigned((8'ha6))) ?
                      {reg2851} : ((forvar2855 <<< forvar2855) ?
                          "axiW2PBUwJx9URPtDFV5xUx" : $signed(reg2849)))) ?
                  $unsigned($signed("OCmzqQqJtGUNZ1ZW")) : "8O");
              reg2864 <= (reg2852[(5'h12):(1'h1)] > $unsigned("XZ5Lkf"));
            end
        end
      reg2865 <= (($unsigned($signed(reg2847[(1'h0):(1'h0)])) ?
          ($unsigned($signed(forvar2848)) ?
              $signed((~^forvar2853)) : $signed((reg2862 & reg2852))) : ({(^reg2851)} ?
              (^~(-reg2861)) : (-$signed(forvar2853)))) << (forvar2853[(3'h5):(1'h0)] ?
          "A45bmgm3YNkuM9RE5" : $signed(("84uVDt2" + wire2845[(3'h5):(3'h4)]))));
      reg2866 <= $unsigned((reg2847 ^ reg2857[(4'hb):(4'h8)]));
      reg2867 <= $signed({(&wire2843[(4'hc):(3'h7)]), reg2851[(2'h2):(1'h1)]});
      for (forvar2868 = (1'h0); (forvar2868 < (3'h4)); forvar2868 = (forvar2868 + (1'h1)))
        begin
          for (forvar2869 = (1'h0); (forvar2869 < (3'h5)); forvar2869 = (forvar2869 + (1'h1)))
            begin
              reg2870 <= (reg2847 ?
                  forvar2853[(3'h4):(1'h0)] : $unsigned($unsigned((&reg2863[(4'h8):(3'h4)]))));
              reg2871 <= ($signed((reg2849 ?
                      reg2851 : ($signed(reg2859) != "KWx0E8g"))) ?
                  wire2843 : $unsigned(reg2856[(5'h11):(3'h4)]));
              reg2872 = {$unsigned((reg2864[(1'h1):(1'h1)] ?
                      $signed((~reg2867)) : reg2862)),
                  ($signed("e4XFiZAMHdawxRwx3tPRgAGa") | ((reg2861[(1'h0):(1'h0)] ?
                      {wire2843} : $signed(reg2858)) <<< ("bSOtVLKTIhyeXgWKRd4la3w" << reg2850)))};
              for (forvar2873 = (1'h0); (forvar2873 < (1'h1)); forvar2873 = (forvar2873 + (1'h1)))
                begin
                  reg2874 <= (forvar2869[(3'h4):(3'h4)] ?
                      ({$signed("duqsvPyIBKBODztSlPoEQyc5"),
                              forvar2853[(3'h4):(3'h4)]} ?
                          ("EtG2" ^~ (~&$signed(reg2859))) : "dtW0KkS") : $signed(reg2866));
                  reg2875 <= ($signed("V6lwEOsZl13HN9Tb") < {$unsigned((&(reg2863 + reg2858)))});
                  reg2876 <= (+"gmDZADZAg8bZIQPm5J6dvg5");
                  reg2877 = "26pyMD9zixkoCx0DRy3H8";
                  reg2878 <= {(($unsigned($unsigned(forvar2869)) ^ "yw6") * (~&reg2858[(1'h0):(1'h0)])),
                      $signed((~{(wire2843 >>> forvar2855)}))};
                end
            end
          reg2879 <= $unsigned(wire2843[(4'hb):(4'hb)]);
          for (forvar2880 = (1'h0); (forvar2880 < (1'h0)); forvar2880 = (forvar2880 + (1'h1)))
            begin
              reg2881 <= "AcTtWMuPF";
            end
          reg2882 = $unsigned($signed((|$signed($unsigned(reg2859)))));
          reg2883 = "3lWOyWDLDtb0rXr81ldckt8p";
          for (forvar2884 = (1'h0); (forvar2884 < (1'h0)); forvar2884 = (forvar2884 + (1'h1)))
            begin
              reg2885 = forvar2873[(3'h5):(3'h5)];
              reg2886 = (reg2876[(3'h4):(2'h2)] ?
                  $signed("7HRshVI53huiVk1Mcd") : $signed($unsigned(reg2867[(3'h5):(1'h1)])));
              reg2887 <= {$unsigned("Zwq0gmiVOg")};
              reg2888 <= reg2863[(3'h7):(2'h3)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg2889 <= (reg2883 ?
          $unsigned("dloU4R1zqmmegwM") : $signed($unsigned((^~forvar2853[(4'h8):(1'h1)]))));
    end
  assign wire2890 = "mLUo55qn";
  always
    @(posedge clk) begin
      reg2891 <= (reg2870[(4'h8):(3'h5)] ^ $unsigned(reg2852[(2'h2):(1'h0)]));
      reg2892 = "oydhGVM4prflo";
      reg2893 = reg2865;
      for (forvar2894 = (1'h0); (forvar2894 < (3'h5)); forvar2894 = (forvar2894 + (1'h1)))
        begin
          reg2895 = ((($signed($unsigned((7'h48))) << $signed((!(8'hb4)))) ?
                  (~$signed((wire2845 ?
                      reg2859 : reg2882))) : (+$unsigned("Ke1m5"))) ?
              (reg2863[(3'h6):(2'h3)] >= {"t9JANtZ8UNP",
                  reg2863[(2'h3):(1'h0)]}) : {("m" >= (|(!(8'h9e))))});
          reg2896 <= reg2862[(4'h8):(1'h0)];
          reg2897 <= "QqUnMrd";
          reg2898 <= (~(!"iJueVnLPuBey"));
        end
      if ($unsigned({$unsigned($signed((!forvar2853))), $unsigned(reg2856)}))
        begin
          reg2899 <= (8'ha0);
          reg2900 <= $unsigned("8fsOTfrSU67L4");
          reg2901 <= ((reg2889 ?
                  ($unsigned(forvar2860[(5'h13):(5'h12)]) | ((reg2889 ?
                          reg2878 : reg2863) ?
                      $signed(forvar2869) : (forvar2873 << reg2872))) : ({"IHK64lZm581FvhSlJWeqx",
                      "gUnGCFJEnGBv"} == reg2864)) ?
              forvar2848[(3'h4):(1'h1)] : reg2883);
          reg2902 <= {{(($signed(forvar2873) ?
                          $unsigned(reg2883) : $unsigned(reg2852)) ?
                      $unsigned($unsigned(reg2858)) : reg2874)},
              ($signed(reg2870) ?
                  reg2858[(3'h4):(2'h3)] : ($signed((reg2889 >>> reg2893)) || reg2883))};
          reg2903 <= $unsigned(({$signed($signed((7'h47))),
              ($unsigned(wire2844) ?
                  $unsigned((7'h44)) : {reg2866,
                      reg2892})} - ($signed(reg2877) ?
              {(7'h4d)} : $signed((^(8'hab))))));
        end
      else
        begin
          for (forvar2899 = (1'h0); (forvar2899 < (3'h5)); forvar2899 = (forvar2899 + (1'h1)))
            begin
              reg2900 = reg2885;
              reg2901 = forvar2868[(3'h4):(1'h1)];
              for (forvar2902 = (1'h0); (forvar2902 < (2'h2)); forvar2902 = (forvar2902 + (1'h1)))
                begin
                  reg2903 <= $unsigned("8qZs9g7yfH1v");
                end
              reg2904 <= "YXd49HW2GtC";
              reg2905 <= ((!(!("WPo49SOBzls3gZKl8ZXI6o" ?
                      reg2849 : ((8'hb5) ? forvar2880 : (7'h43))))) ?
                  (reg2886 ?
                      forvar2899[(2'h2):(1'h0)] : (^$unsigned({reg2867,
                          reg2879}))) : (8'hbf));
              reg2906 <= "fOTaGYbQ8AI0wW";
            end
          for (forvar2907 = (1'h0); (forvar2907 < (1'h0)); forvar2907 = (forvar2907 + (1'h1)))
            begin
              if ($signed("QkwckQr8fwqYe"))
                begin
                  reg2908 <= $unsigned(reg2885[(3'h5):(1'h1)]);
                  reg2909 <= "wtn";
                  reg2910 <= reg2864[(1'h0):(1'h0)];
                  reg2911 = {$signed(forvar2899), $signed((~^{"2"}))};
                  reg2912 <= (8'h9e);
                  reg2913 <= ($signed((8'ha4)) & $unsigned($unsigned($signed(forvar2853))));
                end
              else
                begin
                  reg2908 <= ({("k0Ntam9wTz6m" || $unsigned($unsigned(reg2886))),
                      reg2911[(2'h2):(1'h0)]} >= "YnBK");
                  reg2909 = wire2845[(3'h4):(3'h4)];
                  reg2910 <= $unsigned((($unsigned((forvar2848 >>> reg2849)) ?
                          {((7'h4d) <= forvar2880),
                              "Z"} : $unsigned((forvar2848 && (7'h4d)))) ?
                      $signed((!reg2887[(1'h1):(1'h0)])) : ((-$signed((8'hba))) ?
                          reg2887 : (^reg2852))));
                  reg2911 <= reg2909[(2'h2):(1'h0)];
                end
              reg2914 = (reg2852[(4'hb):(1'h0)] >>> $unsigned((8'hb5)));
              reg2915 <= $unsigned($unsigned((~&$signed(reg2854))));
              reg2916 <= $signed(reg2856);
              reg2917 <= ($unsigned((((forvar2853 * wire2890) ?
                      reg2891 : $signed(reg2891)) - reg2915)) ?
                  (~&($signed({reg2859, reg2866}) ?
                      reg2849 : "dGwpXHSsLYQ4OsHoSxdUhVA")) : forvar2902[(4'hd):(4'h9)]);
              reg2918 = reg2905[(2'h3):(2'h2)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg2919 <= $signed((reg2899 * $signed(($signed(reg2854) + $unsigned(wire2846)))));
      reg2920 <= (8'hbd);
      reg2921 <= (((((reg2885 && (8'hb4)) ? {forvar2884} : "8o") ?
          $signed((wire2846 <= reg2871)) : ((reg2854 && reg2916) >> (-reg2886))) == $unsigned(reg2901)) < "oT01YdwChgSVVt");
      for (forvar2922 = (1'h0); (forvar2922 < (3'h4)); forvar2922 = (forvar2922 + (1'h1)))
        begin
          reg2923 <= ((({{reg2866}} >>> (~&(reg2912 ? forvar2880 : reg2850))) ?
                  reg2877[(1'h0):(1'h0)] : (~|"")) ?
              $signed((8'hb3)) : $unsigned("kOZr"));
          reg2924 <= (8'haf);
          for (forvar2925 = (1'h0); (forvar2925 < (2'h3)); forvar2925 = (forvar2925 + (1'h1)))
            begin
              reg2926 <= ($unsigned(reg2852) ?
                  (|"QypnNYlsQ5NhT") : "fTfD1y1kDMbN");
              reg2927 <= ("FWt68rhRlPgC9k9vSDinrMq" == forvar2925[(4'hf):(3'h4)]);
              reg2928 <= {($unsigned(($unsigned(reg2900) > (~^reg2874))) <= "Uc62zNwL")};
              reg2929 <= "UVA8mgEYGnkGSVgvqk";
              reg2930 = $unsigned((~^reg2897[(3'h7):(2'h3)]));
              if ((~|(($signed((reg2905 <<< (8'hae))) ?
                  reg2904[(3'h5):(2'h2)] : $signed("ER0ODT3xhqxsBaVUX")) <= (^~(~$unsigned(forvar2880))))))
                begin
                  reg2931 <= (~$signed((!$signed(reg2859[(3'h4):(3'h4)]))));
                end
              else
                begin
                  reg2931 <= forvar2869[(4'hd):(4'hd)];
                  reg2932 <= (reg2851[(1'h0):(1'h0)] ?
                      ($unsigned(reg2865) ?
                          $unsigned(forvar2907[(2'h3):(2'h2)]) : "lYKzwrFJ") : (&(wire2845[(2'h2):(1'h1)] && "OPm")));
                  reg2933 = ((&(reg2896[(2'h3):(2'h2)] ?
                      ((reg2885 - reg2924) + "cpaiawIGQb") : $unsigned((reg2857 ?
                          forvar2855 : wire2842)))) <= (&((&reg2910) ?
                      "Dd4Fewuu" : forvar2869)));
                  reg2934 <= "PsDHr";
                  reg2935 <= "UO2f0hJX";
                  reg2936 <= reg2916[(4'h8):(2'h2)];
                end
            end
          reg2937 <= "9Y0oNC";
          if (reg2924)
            begin
              reg2938 <= (wire2890 ?
                  ($signed((+(+forvar2868))) ?
                      ("RiQ3EDEU49kx" ?
                          reg2914[(5'h17):(1'h0)] : reg2896) : {(~(|forvar2894)),
                          $signed("be1yuwHn5eMN")}) : $signed(forvar2848));
              reg2939 = (7'h42);
              reg2940 <= reg2864[(1'h0):(1'h0)];
            end
          else
            begin
              for (forvar2938 = (1'h0); (forvar2938 < (3'h4)); forvar2938 = (forvar2938 + (1'h1)))
                begin
                  reg2939 = reg2902[(1'h1):(1'h1)];
                  reg2940 <= (|$unsigned(forvar2873));
                  reg2941 = $signed($unsigned(reg2898));
                  reg2942 = $unsigned($signed(($unsigned(reg2857) != ((reg2899 || reg2926) ?
                      reg2906 : {(7'h4a), reg2933}))));
                  reg2943 <= (-((^~(reg2940 || reg2917)) != $signed((^reg2849))));
                end
              reg2944 <= $signed($unsigned(reg2864[(1'h0):(1'h0)]));
              for (forvar2945 = (1'h0); (forvar2945 < (1'h1)); forvar2945 = (forvar2945 + (1'h1)))
                begin
                  reg2946 <= $signed((("hhPuOPTqSZz9tRebRyBXDovEX" ?
                          reg2864[(1'h1):(1'h1)] : ($unsigned(forvar2873) ~^ "bHOCnay9mD")) ?
                      (^~(reg2901 ?
                          (reg2912 ?
                              reg2875 : reg2930) : reg2917[(4'ha):(3'h6)])) : (reg2913[(1'h0):(1'h0)] <= (~|$signed(reg2903)))));
                end
              for (forvar2947 = (1'h0); (forvar2947 < (1'h1)); forvar2947 = (forvar2947 + (1'h1)))
                begin
                  reg2948 <= "x325pdQvUKziZ";
                  reg2949 <= "hdvVcxWQAYImNr";
                  reg2950 <= (((((reg2905 >= reg2910) == $signed(reg2943)) ?
                      (reg2946 != ((8'hae) ?
                          reg2891 : (7'h4a))) : $signed("GRefP3rsgNlWIL7sMURzBDOC")) <<< $signed($signed($signed(reg2901)))) - $signed(reg2889[(3'h4):(2'h2)]));
                  reg2951 <= reg2914[(5'h10):(4'hf)];
                  reg2952 = (~^"PYceSfV4v1H3EN0zqfi");
                  reg2953 <= $signed("5DJK6b1N7QpNHXooom6rN9");
                end
            end
        end
      reg2954 <= {$signed(reg2934)};
    end
  assign wire2955 = (|(8'had));
  always
    @(posedge clk) begin
      reg2956 = "vgd5SPh1VHkc84nDfsa902q";
      reg2957 <= (($unsigned("UnVPU2gPW") + (forvar2947[(4'he):(1'h0)] > ($unsigned(reg2920) < (reg2850 == reg2913)))) != forvar2945);
      reg2958 <= (reg2929 < (^~(reg2881 <= "e")));
      for (forvar2959 = (1'h0); (forvar2959 < (2'h3)); forvar2959 = (forvar2959 + (1'h1)))
        begin
          reg2960 <= (8'hac);
          if ((($signed(({forvar2907} ? (!reg2930) : (^~(8'hba)))) ?
                  {wire2844} : $signed((-(&reg2886)))) ?
              {(&$unsigned((wire2955 ?
                      (8'ha9) : forvar2868)))} : (|((^reg2895[(4'h9):(3'h7)]) ?
                  $signed({reg2902}) : (reg2856 < (reg2878 ?
                      reg2920 : (8'ha8)))))))
            begin
              reg2961 <= $signed($unsigned((forvar2894 ?
                  "NKCe0CaNbdBe" : reg2954[(1'h1):(1'h1)])));
            end
          else
            begin
              for (forvar2961 = (1'h0); (forvar2961 < (1'h1)); forvar2961 = (forvar2961 + (1'h1)))
                begin
                  reg2962 <= {$signed((wire2955[(5'h11):(4'h9)] ^ $signed("0hWDR3Q18dZN5UQ8gOEn"))),
                      "SbvuUDIT"};
                  reg2963 <= forvar2945[(4'ha):(3'h5)];
                end
              reg2964 = (reg2861 - (8'h9d));
            end
          reg2965 <= $unsigned(((reg2948 ?
                  reg2877[(4'h8):(2'h2)] : $unsigned($signed(wire2845))) ?
              $unsigned(($signed((8'h9e)) | $unsigned(reg2940))) : "tlSwvOCvXriTCOX"));
          reg2966 <= (~(8'hb5));
        end
      reg2967 = ($signed((($signed(reg2948) ?
          reg2852[(1'h0):(1'h0)] : reg2949[(1'h1):(1'h1)]) <= $unsigned($signed((7'h49))))) & wire2846[(2'h2):(1'h1)]);
      reg2968 <= forvar2961;
    end
  always
    @(posedge clk) begin
      reg2969 <= (^(forvar2947 == $signed(((forvar2884 ? wire2844 : reg2951) ?
          (~|forvar2902) : (reg2949 ? reg2905 : reg2856)))));
      for (forvar2970 = (1'h0); (forvar2970 < (1'h0)); forvar2970 = (forvar2970 + (1'h1)))
        begin
          for (forvar2971 = (1'h0); (forvar2971 < (1'h1)); forvar2971 = (forvar2971 + (1'h1)))
            begin
              reg2972 <= $signed(((reg2870[(3'h6):(2'h3)] ?
                      $signed((!reg2899)) : {"wBy"}) ?
                  $signed($signed(((7'h42) ?
                      reg2924 : forvar2880))) : $unsigned((reg2921[(4'hb):(4'h9)] >>> (reg2924 != reg2927)))));
              reg2973 = (^reg2886[(1'h1):(1'h1)]);
              reg2974 = $unsigned({{reg2867[(2'h3):(2'h2)], (7'h48)}});
              reg2975 <= $signed(reg2909);
              reg2976 <= forvar2907;
              reg2977 <= (^~reg2899);
            end
        end
      reg2978 = (~$signed("TgRI1ZJIyQzg25366rJf"));
      reg2979 <= $signed(reg2911);
    end
  always
    @(posedge clk) begin
      reg2980 <= ((~|{$unsigned(reg2963[(2'h3):(2'h2)]),
              (reg2877[(1'h0):(1'h0)] - "PluK36YvikGEsHYqB9D5T")}) ?
          reg2891 : ((reg2857 ~^ forvar2894) ?
              reg2954[(2'h3):(1'h0)] : (("O2ZxNbErbxD" ?
                      reg2847[(1'h0):(1'h0)] : "wcrB5WOar") ?
                  $signed(reg2976[(2'h3):(1'h0)]) : (^"EZrvMaFl5qVuI4CH"))));
    end
  assign wire2981 = {reg2866[(4'hc):(1'h1)]};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2781  (y, clk, wire2785, wire2784, wire2783, wire2782);
  output wire [(32'h2f2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h18):(1'h0)] wire2785;
  input wire [(5'h1a):(1'h0)] wire2784;
  input wire [(5'h18):(1'h0)] wire2783;
  input wire signed [(5'h13):(1'h0)] wire2782;
  reg [(2'h3):(1'h0)] reg2838 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2837 = (1'h0);
  reg [(4'hb):(1'h0)] reg2836 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2835 = (1'h0);
  reg [(2'h3):(1'h0)] reg2834 = (1'h0);
  reg [(4'he):(1'h0)] reg2833 = (1'h0);
  reg [(5'h17):(1'h0)] reg2832 = (1'h0);
  reg [(4'h9):(1'h0)] reg2831 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2830 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2829 = (1'h0);
  reg [(3'h6):(1'h0)] reg2828 = (1'h0);
  reg [(4'h8):(1'h0)] reg2827 = (1'h0);
  reg [(5'h14):(1'h0)] reg2826 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2825 = (1'h0);
  reg [(4'h9):(1'h0)] reg2820 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2818 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2824 = (1'h0);
  reg [(5'h15):(1'h0)] reg2823 = (1'h0);
  reg [(5'h10):(1'h0)] reg2822 = (1'h0);
  reg [(2'h3):(1'h0)] reg2821 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2820 = (1'h0);
  reg [(5'h12):(1'h0)] reg2819 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2818 = (1'h0);
  reg [(4'ha):(1'h0)] reg2817 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2816 = (1'h0);
  wire [(4'hb):(1'h0)] wire2815;
  wire signed [(5'h19):(1'h0)] wire2814;
  reg signed [(5'h19):(1'h0)] reg2813 = (1'h0);
  reg [(3'h6):(1'h0)] reg2812 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2811 = (1'h0);
  wire [(3'h6):(1'h0)] wire2810;
  reg [(4'hb):(1'h0)] reg2809 = (1'h0);
  reg [(5'h15):(1'h0)] reg2808 = (1'h0);
  reg [(5'h17):(1'h0)] reg2807 = (1'h0);
  reg [(4'hc):(1'h0)] reg2806 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2805 = (1'h0);
  reg [(2'h3):(1'h0)] reg2804 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2803 = (1'h0);
  reg [(5'h16):(1'h0)] reg2802 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2801 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2800 = (1'h0);
  reg [(5'h18):(1'h0)] reg2799 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2798 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2797 = (1'h0);
  reg [(3'h5):(1'h0)] reg2796 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2795 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2794 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2793 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2792 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2791 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2790 = (1'h0);
  reg [(5'h12):(1'h0)] reg2789 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2788 = (1'h0);
  reg [(5'h19):(1'h0)] reg2787 = (1'h0);
  reg [(3'h6):(1'h0)] reg2786 = (1'h0);
  assign y = {reg2838,
                 reg2837,
                 reg2836,
                 reg2835,
                 reg2834,
                 reg2833,
                 reg2832,
                 reg2831,
                 reg2830,
                 reg2829,
                 reg2828,
                 reg2827,
                 reg2826,
                 forvar2825,
                 reg2820,
                 forvar2818,
                 reg2824,
                 reg2823,
                 reg2822,
                 reg2821,
                 forvar2820,
                 reg2819,
                 reg2818,
                 reg2817,
                 forvar2816,
                 wire2815,
                 wire2814,
                 reg2813,
                 reg2812,
                 reg2811,
                 wire2810,
                 reg2809,
                 reg2808,
                 reg2807,
                 reg2806,
                 reg2805,
                 reg2804,
                 reg2803,
                 reg2802,
                 forvar2801,
                 reg2800,
                 reg2799,
                 reg2798,
                 forvar2797,
                 reg2796,
                 forvar2795,
                 reg2794,
                 reg2793,
                 reg2792,
                 forvar2791,
                 reg2790,
                 reg2789,
                 reg2788,
                 reg2787,
                 reg2786,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg2786 <= (!wire2785);
      reg2787 = (|($signed(wire2783[(4'ha):(4'ha)]) ?
          (($unsigned(reg2786) ?
              (reg2786 ?
                  wire2783 : wire2784) : $signed(wire2785)) ^ $signed(wire2784[(5'h18):(5'h18)])) : $signed($signed($signed(wire2783)))));
      reg2788 = wire2785[(5'h13):(4'hd)];
      reg2789 <= "4YLzZsDEnoam0DYcJ";
      reg2790 <= (|reg2788[(5'h13):(5'h12)]);
    end
  always
    @(posedge clk) begin
      for (forvar2791 = (1'h0); (forvar2791 < (2'h3)); forvar2791 = (forvar2791 + (1'h1)))
        begin
          reg2792 <= (+(wire2782 << wire2782));
          reg2793 <= (("P3VJNIzbESQbfexVbg3" <= $signed($signed((~&(8'h9d))))) >> ((+((reg2789 + reg2792) || $unsigned(wire2785))) && reg2792[(4'hd):(4'hc)]));
          reg2794 = (!({(^(+(8'hbc)))} ?
              reg2793 : (reg2787[(3'h7):(3'h7)] ?
                  "5To1XOe80i" : $unsigned($unsigned(reg2793)))));
          for (forvar2795 = (1'h0); (forvar2795 < (3'h4)); forvar2795 = (forvar2795 + (1'h1)))
            begin
              reg2796 <= reg2793;
              for (forvar2797 = (1'h0); (forvar2797 < (2'h3)); forvar2797 = (forvar2797 + (1'h1)))
                begin
                  reg2798 = $unsigned(("zZlkcKUzGzkGC6UMS" ?
                      $unsigned(reg2788[(5'h10):(4'hf)]) : ("B4BC88dPQbZx" << $signed({(8'ha3)}))));
                  reg2799 <= $unsigned((reg2798[(4'hc):(3'h6)] ~^ ((^~wire2783) ?
                      ("OTENT4NlfUD" ?
                          {reg2786} : reg2796[(3'h5):(3'h5)]) : (reg2792 ?
                          "FVU7hBtBz" : (reg2792 <<< reg2790)))));
                end
              reg2800 <= $unsigned($signed((~{$unsigned(reg2796)})));
              for (forvar2801 = (1'h0); (forvar2801 < (1'h0)); forvar2801 = (forvar2801 + (1'h1)))
                begin
                  reg2802 <= ((reg2794[(1'h1):(1'h1)] * (~&($signed(reg2800) >>> $signed(reg2789)))) << (~wire2782));
                  reg2803 <= $signed($signed(reg2788[(5'h15):(4'h9)]));
                  reg2804 = $unsigned(reg2793[(4'hf):(4'hd)]);
                end
            end
          reg2805 = (wire2783 ?
              forvar2791 : ($unsigned((reg2800 - $unsigned(reg2802))) ?
                  (~"hUMedlLRaWLo") : reg2793[(4'h8):(3'h6)]));
        end
      reg2806 <= $signed((reg2804[(1'h1):(1'h0)] ~^ (&({reg2786} ~^ "qmr55Po"))));
      reg2807 <= ($unsigned((~&wire2782)) ?
          $signed($unsigned((^$unsigned(reg2802)))) : ({(reg2790[(5'h15):(4'h8)] < $unsigned(reg2802)),
                  $signed({reg2786, reg2800})} ?
              (reg2799[(5'h12):(2'h3)] ?
                  $signed(wire2782) : (+reg2796)) : reg2790));
      reg2808 <= wire2784;
      reg2809 <= (~|(reg2808[(4'he):(4'h8)] ?
          {($signed(reg2790) | $unsigned(reg2799)),
              $signed((~|reg2800))} : $unsigned((((8'ha3) ? reg2793 : reg2796) ?
              $signed(wire2782) : {(7'h49)}))));
    end
  assign wire2810 = {(reg2803 ? (!$unsigned(forvar2801)) : {forvar2797}),
                        forvar2801};
  always
    @(posedge clk) begin
      reg2811 <= reg2799[(5'h17):(4'hd)];
      reg2812 = reg2809[(4'ha):(3'h7)];
      reg2813 <= "HhBKhLKXEZ89qBCGQVmSwsrU";
    end
  assign wire2814 = reg2788;
  assign wire2815 = $signed(wire2810[(2'h2):(2'h2)]);
  always
    @(posedge clk) begin
      for (forvar2816 = (1'h0); (forvar2816 < (3'h5)); forvar2816 = (forvar2816 + (1'h1)))
        begin
          if (($signed((!reg2794[(4'h8):(4'h8)])) ?
              (forvar2791 ?
                  "" : (reg2787 <= wire2815[(4'h9):(3'h6)])) : "nck6gcVQtPM2wWa8dzUQJvVS"))
            begin
              reg2817 = forvar2791[(2'h2):(1'h1)];
              reg2818 = "hrRur9gvAP";
              reg2819 <= (^~reg2809[(2'h3):(2'h2)]);
              for (forvar2820 = (1'h0); (forvar2820 < (2'h3)); forvar2820 = (forvar2820 + (1'h1)))
                begin
                  reg2821 <= (&reg2792[(4'hf):(2'h3)]);
                  reg2822 = "zYaqW2QHsE0ZCz";
                  reg2823 = ($signed($unsigned({$signed(reg2786)})) ^~ {wire2784,
                      wire2784[(5'h19):(5'h13)]});
                end
              reg2824 <= {"ONqUOKBqQK"};
            end
          else
            begin
              reg2817 <= (reg2794 ? "dVQtfQ5kL" : reg2821);
              for (forvar2818 = (1'h0); (forvar2818 < (3'h5)); forvar2818 = (forvar2818 + (1'h1)))
                begin
                  reg2819 <= $signed((~wire2815[(4'h9):(4'h9)]));
                  reg2820 <= reg2794;
                  reg2821 <= reg2794[(4'h9):(1'h0)];
                  reg2822 <= $signed($signed((~&$unsigned(((8'ha6) && forvar2818)))));
                  reg2823 = reg2804;
                  reg2824 <= (reg2817 ?
                      reg2805[(3'h5):(1'h1)] : ($signed(((reg2821 ?
                              reg2808 : forvar2820) ?
                          $unsigned(reg2821) : $unsigned(forvar2820))) << (($signed(reg2790) ?
                              forvar2816[(2'h2):(1'h0)] : (~^reg2803)) ?
                          ((^~(8'ha2)) ^ (~|reg2818)) : "boDKT")));
                end
              for (forvar2825 = (1'h0); (forvar2825 < (3'h4)); forvar2825 = (forvar2825 + (1'h1)))
                begin
                  reg2826 <= (~&wire2785[(2'h3):(2'h2)]);
                  reg2827 <= (forvar2797[(1'h0):(1'h0)] ?
                      "" : ((reg2800[(3'h4):(2'h2)] ?
                          reg2798 : "15nPrGE6") && reg2800));
                  reg2828 <= ((reg2817 ?
                      (~^($unsigned(reg2803) >= (~^reg2817))) : ($signed($signed(reg2788)) ^ (-$unsigned(forvar2820)))) >> ($signed(((~wire2783) != (~^reg2812))) ?
                      reg2813 : $signed({((8'haa) ? (7'h42) : wire2784)})));
                  reg2829 <= (~"OWX7Uiyi");
                  reg2830 <= (($signed((^~(reg2818 >>> reg2807))) || ((8'hbf) & {(reg2788 ?
                          (7'h40) : (8'hbe))})) | reg2794[(3'h5):(3'h5)]);
                end
            end
          reg2831 = (reg2830[(3'h5):(3'h4)] || {(~$signed($unsigned(wire2782)))});
        end
      reg2832 <= $signed($unsigned("P0BD"));
      reg2833 <= (~^$unsigned($signed(reg2787)));
      reg2834 <= wire2814;
    end
  always
    @(posedge clk) begin
      reg2835 <= (reg2830 | wire2815[(1'h1):(1'h0)]);
      reg2836 = (^~reg2800);
      reg2837 <= forvar2791[(4'h8):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg2838 <= ("abe7bSPxHnEeYHwwb" != ((!reg2796[(2'h2):(2'h2)]) != ($signed(reg2828[(3'h6):(1'h0)]) ?
          ((reg2790 ? reg2836 : reg2836) | $unsigned((8'h9e))) : "Go")));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2696
#( parameter param2766 = (~(((((8'hac) ? (8'ha6) : (8'ha5)) ? (+(8'ha6)) : ((7'h47) ? (7'h46) : (7'h4d))) == ((~|(7'h41)) & {(7'h4b), (8'ha7)})) ? (((-(8'ha8)) || ((8'h9f) | (8'hae))) && ((&(7'h4d)) < {(8'hb8)})) : ((+((8'hac) && (8'ha4))) ? (((8'h9e) ? (8'h9e) : (8'hac)) ? ((8'h9e) ? (7'h42) : (8'hab)) : (+(7'h47))) : (&((7'h48) ? (7'h4d) : (8'hb4)))))) )
(y, clk, wire2700, wire2699, wire2698, wire2697);
  output wire [(32'h381):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire2700;
  input wire [(4'h8):(1'h0)] wire2699;
  input wire signed [(5'h14):(1'h0)] wire2698;
  input wire [(5'h15):(1'h0)] wire2697;
  wire [(3'h5):(1'h0)] wire2765;
  reg signed [(5'h15):(1'h0)] reg2764 = (1'h0);
  reg [(5'h18):(1'h0)] reg2763 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2762 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2761 = (1'h0);
  reg [(5'h19):(1'h0)] reg2760 = (1'h0);
  reg [(4'h8):(1'h0)] reg2759 = (1'h0);
  reg [(3'h4):(1'h0)] reg2758 = (1'h0);
  reg [(4'hb):(1'h0)] reg2757 = (1'h0);
  reg [(4'h9):(1'h0)] reg2756 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2755 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2754 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2753 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2752 = (1'h0);
  reg [(3'h5):(1'h0)] reg2751 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2750 = (1'h0);
  reg [(3'h7):(1'h0)] reg2749 = (1'h0);
  reg [(5'h10):(1'h0)] reg2748 = (1'h0);
  reg [(4'hd):(1'h0)] reg2747 = (1'h0);
  reg [(5'h15):(1'h0)] reg2746 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2745 = (1'h0);
  reg [(4'h8):(1'h0)] reg2744 = (1'h0);
  reg [(5'h12):(1'h0)] reg2743 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2742 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2741 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2740 = (1'h0);
  reg [(5'h15):(1'h0)] reg2739 = (1'h0);
  reg [(4'he):(1'h0)] reg2738 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2737 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2736 = (1'h0);
  reg [(4'h9):(1'h0)] reg2735 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2734 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire2733;
  wire [(5'h13):(1'h0)] wire2732;
  wire signed [(5'h16):(1'h0)] wire2731;
  reg signed [(4'hb):(1'h0)] reg2730 = (1'h0);
  reg [(5'h11):(1'h0)] reg2729 = (1'h0);
  reg [(4'hd):(1'h0)] reg2728 = (1'h0);
  wire [(4'hf):(1'h0)] wire2727;
  wire [(4'h9):(1'h0)] wire2726;
  reg signed [(3'h5):(1'h0)] reg2725 = (1'h0);
  reg [(4'hd):(1'h0)] reg2724 = (1'h0);
  reg [(3'h4):(1'h0)] reg2723 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2722 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2721 = (1'h0);
  reg [(2'h2):(1'h0)] reg2720 = (1'h0);
  reg [(5'h18):(1'h0)] reg2719 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2718 = (1'h0);
  reg [(5'h18):(1'h0)] reg2717 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2716 = (1'h0);
  reg [(4'h9):(1'h0)] reg2715 = (1'h0);
  reg [(3'h7):(1'h0)] reg2714 = (1'h0);
  reg [(5'h11):(1'h0)] reg2713 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2712 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2711 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2710 = (1'h0);
  reg [(5'h11):(1'h0)] reg2709 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2708 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2707 = (1'h0);
  reg [(4'hf):(1'h0)] reg2706 = (1'h0);
  reg [(5'h17):(1'h0)] reg2705 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2704 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2703 = (1'h0);
  reg [(3'h6):(1'h0)] reg2702 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2701 = (1'h0);
  assign y = {wire2765,
                 reg2764,
                 reg2763,
                 reg2762,
                 reg2761,
                 reg2760,
                 reg2759,
                 reg2758,
                 reg2757,
                 reg2756,
                 reg2755,
                 reg2754,
                 reg2753,
                 reg2752,
                 reg2751,
                 forvar2750,
                 reg2749,
                 reg2748,
                 reg2747,
                 reg2746,
                 reg2745,
                 reg2744,
                 reg2743,
                 reg2742,
                 forvar2741,
                 forvar2740,
                 reg2739,
                 reg2738,
                 forvar2737,
                 reg2736,
                 reg2735,
                 reg2734,
                 wire2733,
                 wire2732,
                 wire2731,
                 reg2730,
                 reg2729,
                 reg2728,
                 wire2727,
                 wire2726,
                 reg2725,
                 reg2724,
                 reg2723,
                 reg2722,
                 reg2721,
                 reg2720,
                 reg2719,
                 forvar2718,
                 reg2717,
                 reg2716,
                 reg2715,
                 reg2714,
                 reg2713,
                 forvar2712,
                 forvar2711,
                 reg2710,
                 reg2709,
                 reg2708,
                 forvar2707,
                 reg2706,
                 reg2705,
                 reg2704,
                 forvar2703,
                 reg2702,
                 reg2701,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg2701 <= wire2699;
      reg2702 = ((~|("f8gYYTRQ8YJndVzgdF0Hh" < ({reg2701,
          wire2698} ~^ (wire2700 << wire2700)))) >> (|(7'h44)));
      for (forvar2703 = (1'h0); (forvar2703 < (3'h5)); forvar2703 = (forvar2703 + (1'h1)))
        begin
          reg2704 <= ((!$unsigned((~^(^forvar2703)))) * reg2702[(2'h3):(1'h0)]);
          reg2705 <= $signed(((forvar2703[(2'h2):(1'h1)] ?
              "grFmXxF1f4GYVAX8kslZVfiUK" : reg2702) == (+(~^(|(8'ha8))))));
          reg2706 <= ($unsigned(wire2698) ^~ $signed((($unsigned(wire2698) + wire2698[(4'ha):(4'h8)]) >= "tpFmw7fQRe")));
          for (forvar2707 = (1'h0); (forvar2707 < (3'h4)); forvar2707 = (forvar2707 + (1'h1)))
            begin
              reg2708 <= ($signed(("AFU5AL1k3gIuSvQ" - {{wire2700}})) && (~(|($unsigned(reg2702) ?
                  reg2701[(3'h6):(1'h1)] : (wire2700 - reg2706)))));
            end
          reg2709 <= forvar2707;
          reg2710 <= {(-(+"1bttNULRl3fUn8Eq")),
              {$signed((wire2700 <= $signed(reg2705))), reg2702}};
        end
    end
  always
    @(posedge clk) begin
      for (forvar2711 = (1'h0); (forvar2711 < (1'h1)); forvar2711 = (forvar2711 + (1'h1)))
        begin
          for (forvar2712 = (1'h0); (forvar2712 < (2'h3)); forvar2712 = (forvar2712 + (1'h1)))
            begin
              reg2713 <= (|"H");
              reg2714 <= ((^$signed($unsigned((reg2705 + forvar2703)))) ?
                  $unsigned((reg2713 ?
                      (^(~reg2710)) : "ZsL1J7sZfyGIPMCMO7OSxCCqh")) : {$signed({(^(8'h9f)),
                          $unsigned(reg2708)})});
              reg2715 <= "0TSxfDLwzExJItb85nk3";
            end
          reg2716 <= wire2697;
        end
      reg2717 <= (~(reg2702 ? "" : $signed(reg2708)));
      for (forvar2718 = (1'h0); (forvar2718 < (1'h1)); forvar2718 = (forvar2718 + (1'h1)))
        begin
          reg2719 <= (forvar2703 <= (forvar2703[(3'h5):(3'h5)] >> $unsigned(reg2714)));
          reg2720 <= {$signed($signed({"6we0", $signed(reg2705)})),
              "LgUGExFie"};
          reg2721 = $unsigned(wire2699[(1'h0):(1'h0)]);
          reg2722 <= $unsigned($signed(({"5NsQVX9HTUY7izRxP6v"} != (((8'ha1) & reg2713) ?
              (reg2714 ? (7'h46) : reg2717) : (reg2709 & wire2698)))));
        end
      reg2723 = (^(reg2719[(2'h2):(1'h1)] < {($signed(reg2716) ?
              (reg2715 ? forvar2718 : wire2699) : wire2699[(3'h4):(1'h1)]),
          $signed((+wire2699))}));
    end
  always
    @(posedge clk) begin
      reg2724 <= (reg2719[(5'h17):(3'h5)] <<< (($unsigned((^~reg2719)) ?
              {reg2714} : $unsigned($signed(wire2699))) ?
          ((+$unsigned(reg2723)) ^ $signed((~&wire2699))) : (~|(&(7'h4a)))));
      reg2725 <= (^~reg2706);
    end
  assign wire2726 = reg2708;
  assign wire2727 = {(("YkF2bPp3z" >= "L") < $unsigned($signed(reg2709))),
                        ($unsigned(reg2714) ? reg2716 : wire2697)};
  always
    @(posedge clk) begin
      reg2728 <= reg2722;
      reg2729 <= "woJwbkiu";
    end
  always
    @(posedge clk) begin
      reg2730 <= $unsigned(reg2725);
    end
  assign wire2731 = reg2715[(2'h3):(1'h1)];
  assign wire2732 = "EHQkTNF";
  assign wire2733 = (^forvar2711[(3'h7):(3'h7)]);
  always
    @(posedge clk) begin
      reg2734 <= {$signed(($signed((8'hb2)) <<< $signed($unsigned(wire2699)))),
          $signed("")};
      reg2735 = $signed(reg2719[(4'hb):(3'h7)]);
      reg2736 = reg2708;
      for (forvar2737 = (1'h0); (forvar2737 < (3'h5)); forvar2737 = (forvar2737 + (1'h1)))
        begin
          reg2738 = "qg2aSOSSyxpGOL";
          reg2739 <= $unsigned((reg2709 ?
              ($signed(((8'hb0) ?
                  wire2727 : reg2706)) != (8'hb9)) : wire2697[(3'h5):(3'h4)]));
          for (forvar2740 = (1'h0); (forvar2740 < (3'h4)); forvar2740 = (forvar2740 + (1'h1)))
            begin
              for (forvar2741 = (1'h0); (forvar2741 < (2'h3)); forvar2741 = (forvar2741 + (1'h1)))
                begin
                  reg2742 = $signed(("WTonE833tnKvw" ?
                      reg2715[(1'h0):(1'h0)] : (((&reg2730) >> $signed(reg2723)) ?
                          {(^forvar2707)} : {(forvar2741 >>> reg2719),
                              $signed(reg2729)})));
                  reg2743 <= reg2705;
                  reg2744 <= (7'h46);
                  reg2745 <= (~|($signed("Nx") ?
                      $signed(reg2723[(2'h3):(1'h0)]) : forvar2737[(1'h1):(1'h0)]));
                  reg2746 <= ($unsigned($unsigned(wire2699[(1'h0):(1'h0)])) ?
                      $unsigned({$signed($unsigned(reg2716)),
                          (~&(reg2715 >>> reg2714))}) : reg2710);
                end
              reg2747 <= ($unsigned($unsigned({(~^reg2701)})) ?
                  (reg2708 >>> {wire2726,
                      reg2736[(3'h6):(1'h0)]}) : $signed($signed((|$signed(forvar2711)))));
              reg2748 <= (wire2727 ?
                  wire2726[(3'h5):(3'h5)] : reg2704[(4'hc):(4'hb)]);
              reg2749 <= forvar2712;
              for (forvar2750 = (1'h0); (forvar2750 < (2'h3)); forvar2750 = (forvar2750 + (1'h1)))
                begin
                  reg2751 = "sdP";
                  reg2752 <= (&($unsigned((forvar2740[(3'h5):(3'h4)] + (reg2721 & wire2700))) ?
                      {"J4e1lCpJlJ3tOW2XW6UOruTYD",
                          $unsigned($unsigned(reg2713))} : forvar2740));
                  reg2753 = (|"r4GBZR41EDmUpvdcQe2kdb");
                  reg2754 <= (reg2738[(4'h8):(3'h7)] ?
                      $unsigned("ESOZm1kzy8Cc") : reg2723[(1'h1):(1'h1)]);
                end
              reg2755 <= "";
            end
          reg2756 <= "WNgpZ5NiMh";
        end
    end
  always
    @(posedge clk) begin
      reg2757 <= (|reg2738[(3'h5):(1'h1)]);
      reg2758 <= "79fLfO";
      reg2759 <= forvar2703[(1'h0):(1'h0)];
      reg2760 <= {$unsigned((|$unsigned((reg2715 ~^ wire2731)))), reg2729};
      reg2761 <= "DosSNS";
    end
  always
    @(posedge clk) begin
      reg2762 <= $unsigned(($signed(reg2709[(4'hc):(2'h3)]) ?
          (reg2706[(2'h3):(2'h2)] == ("LVOOT0HF" ?
              ((7'h41) && (8'h9c)) : (^reg2705))) : $signed($signed("OHUtGslJ0fhHALWV6J8yKB"))));
      reg2763 <= reg2738[(4'hc):(3'h7)];
      reg2764 <= ({(((reg2714 ? reg2721 : reg2758) ?
                  $unsigned(reg2714) : reg2717[(5'h16):(5'h14)]) == forvar2740[(1'h1):(1'h1)]),
              ("UuKTnzZPC0" ?
                  forvar2718[(3'h7):(2'h3)] : forvar2718[(3'h4):(2'h3)])} ?
          reg2701[(3'h7):(3'h4)] : (((|(reg2757 <<< (8'hbb))) ^ "ohxLlBeC4V") | ((8'ha7) ?
              reg2763[(5'h10):(4'h8)] : reg2749)));
    end
  assign wire2765 = {$signed($signed(reg2754[(4'hd):(4'h9)])), forvar2740};
endmodule