(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param2707 = {(((((7'h43) ? (7'h41) : (8'h9c)) == ((8'ha2) != (8'hbf))) ^ ((~(7'h43)) ? ((8'ha9) ^ (8'hb0)) : (~^(8'hab)))) ? (^~{((8'hb4) ? (8'hac) : (8'hb4))}) : ((8'ha1) ? ({(7'h43), (8'hb9)} < ((8'haf) ^ (8'hb1))) : (((7'h43) ? (7'h40) : (8'hb8)) ? ((8'hbf) & (8'ha8)) : ((8'ha9) ? (7'h41) : (8'h9c)))))} )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h3f8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire3;
  input wire signed [(4'hf):(1'h0)] wire2;
  input wire signed [(4'hd):(1'h0)] wire1;
  input wire [(5'h14):(1'h0)] wire0;
  reg [(5'h10):(1'h0)] reg2706 = (1'h0);
  reg [(2'h2):(1'h0)] reg2705 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2704 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2703 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2702 = (1'h0);
  reg [(5'h14):(1'h0)] reg2701 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2700 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2699 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2698 = (1'h0);
  reg [(3'h4):(1'h0)] reg2697 = (1'h0);
  reg [(3'h4):(1'h0)] reg2696 = (1'h0);
  reg [(5'h10):(1'h0)] reg2695 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2694 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2693 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2692 = (1'h0);
  reg [(5'h11):(1'h0)] reg2691 = (1'h0);
  reg [(5'h15):(1'h0)] reg2690 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2689 = (1'h0);
  reg [(5'h11):(1'h0)] reg2688 = (1'h0);
  reg [(4'hd):(1'h0)] reg2687 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2686 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2685 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2684 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2683 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2682 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2681 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2680 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire2678;
  reg [(3'h6):(1'h0)] reg889 = (1'h0);
  wire signed [(4'he):(1'h0)] wire888;
  wire signed [(4'h8):(1'h0)] wire96;
  wire [(4'ha):(1'h0)] wire54;
  wire signed [(4'h8):(1'h0)] wire53;
  reg signed [(4'he):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg51 = (1'h0);
  reg [(4'h9):(1'h0)] forvar50 = (1'h0);
  reg [(3'h7):(1'h0)] reg49 = (1'h0);
  reg [(5'h15):(1'h0)] reg48 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg47 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar46 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg45 = (1'h0);
  reg [(2'h3):(1'h0)] reg44 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar43 = (1'h0);
  reg [(2'h2):(1'h0)] reg42 = (1'h0);
  reg [(4'h8):(1'h0)] reg41 = (1'h0);
  reg [(5'h14):(1'h0)] reg40 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg39 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg38 = (1'h0);
  reg [(4'hb):(1'h0)] reg37 = (1'h0);
  reg [(2'h3):(1'h0)] reg36 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg35 = (1'h0);
  reg [(4'hb):(1'h0)] reg34 = (1'h0);
  reg [(4'hf):(1'h0)] reg33 = (1'h0);
  reg [(4'hf):(1'h0)] reg32 = (1'h0);
  reg [(4'h8):(1'h0)] forvar31 = (1'h0);
  reg [(5'h12):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg29 = (1'h0);
  reg [(3'h5):(1'h0)] forvar28 = (1'h0);
  reg [(3'h6):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg25 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg24 = (1'h0);
  reg [(5'h12):(1'h0)] reg23 = (1'h0);
  reg [(5'h10):(1'h0)] forvar22 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar20 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire19;
  reg signed [(5'h11):(1'h0)] reg18 = (1'h0);
  reg [(4'h9):(1'h0)] reg17 = (1'h0);
  reg [(4'h8):(1'h0)] reg16 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar15 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg14 = (1'h0);
  reg signed [(4'he):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg9 = (1'h0);
  reg [(4'h8):(1'h0)] forvar8 = (1'h0);
  reg [(4'hc):(1'h0)] reg7 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg5 = (1'h0);
  wire [(4'hd):(1'h0)] wire4;
  wire [(5'h14):(1'h0)] wire98;
  wire [(3'h7):(1'h0)] wire886;
  assign y = {reg2706,
                 reg2705,
                 reg2704,
                 reg2703,
                 reg2702,
                 reg2701,
                 forvar2700,
                 reg2699,
                 reg2698,
                 reg2697,
                 reg2696,
                 reg2695,
                 forvar2694,
                 reg2693,
                 forvar2692,
                 reg2691,
                 reg2690,
                 reg2689,
                 reg2688,
                 reg2687,
                 forvar2686,
                 reg2685,
                 reg2684,
                 reg2683,
                 forvar2682,
                 forvar2681,
                 reg2680,
                 wire2678,
                 reg889,
                 wire888,
                 wire96,
                 wire54,
                 wire53,
                 reg52,
                 reg51,
                 forvar50,
                 reg49,
                 reg48,
                 reg47,
                 forvar46,
                 reg45,
                 reg44,
                 forvar43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 forvar31,
                 reg30,
                 reg29,
                 forvar28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 forvar22,
                 reg21,
                 forvar20,
                 wire19,
                 reg18,
                 reg17,
                 reg16,
                 forvar15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 forvar8,
                 reg7,
                 reg6,
                 reg5,
                 wire4,
                 wire98,
                 wire886,
                 (1'h0)};
  assign wire4 = $signed($signed(({wire2[(2'h3):(1'h1)],
                     {wire3, wire2}} >>> $signed((|wire2)))));
  always
    @(posedge clk) begin
      reg5 = $signed(wire4[(2'h2):(1'h0)]);
      reg6 <= (~&($signed((wire4[(4'hc):(4'h8)] <<< (wire3 ?
          wire0 : wire4))) <<< $signed(wire2[(2'h3):(2'h3)])));
      reg7 = ((8'hab) ?
          (wire4[(3'h6):(1'h0)] ?
              (+$signed(wire2[(2'h3):(1'h1)])) : (|(((8'hb2) ? wire0 : wire0) ?
                  (reg5 ? wire2 : wire2) : (+wire3)))) : wire1[(4'ha):(3'h6)]);
    end
  always
    @(posedge clk) begin
      for (forvar8 = (1'h0); (forvar8 < (3'h4)); forvar8 = (forvar8 + (1'h1)))
        begin
          reg9 = (8'ha0);
        end
      reg10 <= reg7;
      reg11 <= $signed(($unsigned(wire2[(2'h3):(1'h1)]) != reg5[(5'h10):(4'he)]));
      reg12 = reg5;
    end
  always
    @(posedge clk) begin
      reg13 <= ($unsigned((&$signed($signed(reg10)))) ?
          $unsigned($signed(reg12[(4'h9):(3'h7)])) : {$signed(((forvar8 ?
                      reg6 : reg11) ?
                  (reg5 ? reg5 : forvar8) : reg7[(1'h1):(1'h0)]))});
      reg14 = ($signed({({reg6} ? (reg11 - forvar8) : (wire1 | reg12)),
          ((wire2 & (8'hbe)) ^~ $signed(reg13))}) << $signed($signed(reg12[(2'h3):(1'h0)])));
      for (forvar15 = (1'h0); (forvar15 < (3'h4)); forvar15 = (forvar15 + (1'h1)))
        begin
          reg16 <= wire2[(2'h2):(1'h1)];
          reg17 <= $unsigned({reg7, $signed(reg13[(3'h7):(3'h6)])});
          reg18 <= (!$unsigned(reg7));
        end
    end
  assign wire19 = ((+reg10) || $signed(reg13[(3'h7):(1'h1)]));
  always
    @(posedge clk) begin
      for (forvar20 = (1'h0); (forvar20 < (3'h4)); forvar20 = (forvar20 + (1'h1)))
        begin
          reg21 = (reg10[(3'h6):(3'h6)] ?
              {$signed(reg7), ($unsigned($signed(wire0)) & wire0)} : reg12);
          for (forvar22 = (1'h0); (forvar22 < (3'h4)); forvar22 = (forvar22 + (1'h1)))
            begin
              reg23 = (wire19 ?
                  $unsigned((-((8'haa) << forvar15))) : reg11[(4'ha):(2'h3)]);
              reg24 = (&{(~^((reg5 ? reg7 : wire19) || reg5))});
              reg25 <= {(forvar22 ? $unsigned(wire19) : {(~^wire0)})};
              reg26 = $signed({((8'hab) <= (reg9 ? (~&reg18) : reg6)),
                  reg11[(1'h1):(1'h0)]});
            end
        end
      reg27 <= reg21[(4'h8):(3'h4)];
      for (forvar28 = (1'h0); (forvar28 < (1'h1)); forvar28 = (forvar28 + (1'h1)))
        begin
          reg29 <= reg5[(4'hd):(4'hc)];
        end
      reg30 = (!(({$unsigned(reg12)} ?
              (reg25[(3'h6):(3'h4)] <<< wire0[(5'h12):(4'hf)]) : reg16[(3'h4):(3'h4)]) ?
          forvar20[(4'h8):(4'h8)] : $signed((~|reg16))));
      for (forvar31 = (1'h0); (forvar31 < (2'h2)); forvar31 = (forvar31 + (1'h1)))
        begin
          reg32 <= ((~|{$signed((&(8'ha8)))}) ?
              {$signed(reg21),
                  ($signed((reg18 & forvar8)) ?
                      ((+(8'ha0)) ?
                          (reg11 >>> reg30) : $unsigned(reg17)) : (~^$unsigned(forvar20)))} : forvar22);
          if ($unsigned(forvar31))
            begin
              reg33 <= $unsigned(($signed(((^~reg21) ?
                      (+(8'ha9)) : ((8'ha6) ? (8'ha4) : reg16))) ?
                  reg18[(4'h9):(2'h2)] : reg23));
              reg34 = (|((wire19[(3'h4):(2'h2)] ? (8'hb3) : (^~reg13)) ?
                  (8'hbd) : (~&(+$signed(reg5)))));
              reg35 <= (8'h9c);
              reg36 <= {reg32[(4'hd):(4'hc)]};
              reg37 = (((wire0 ? reg14 : reg27[(3'h6):(2'h2)]) ?
                  $unsigned((~&(~reg35))) : (~{wire4[(3'h4):(1'h0)]})) < $unsigned(((+forvar22[(3'h6):(1'h1)]) ?
                  reg24[(2'h2):(2'h2)] : (~&(reg34 > reg11)))));
            end
          else
            begin
              reg33 <= $signed({reg35});
              reg34 <= wire19;
              reg35 <= $unsigned($signed((^~reg14)));
            end
          reg38 <= (($unsigned($signed(reg23[(3'h6):(3'h4)])) >= ({((8'hbf) == (8'hbe))} ?
                  $signed($signed((8'hae))) : (8'hae))) ?
              $unsigned((reg33[(4'ha):(2'h2)] ~^ {{wire3,
                      wire4}})) : reg17[(3'h4):(3'h4)]);
          reg39 <= $unsigned($unsigned($signed(reg10[(3'h5):(2'h2)])));
        end
    end
  always
    @(posedge clk) begin
      reg40 <= $unsigned(((8'hba) != $unsigned(reg34[(4'h8):(2'h3)])));
    end
  always
    @(posedge clk) begin
      reg41 <= {$unsigned($signed(reg14[(3'h7):(1'h1)]))};
      reg42 = $signed($signed(((^~$signed(forvar31)) | $unsigned((reg26 >>> reg40)))));
    end
  always
    @(posedge clk) begin
      for (forvar43 = (1'h0); (forvar43 < (1'h0)); forvar43 = (forvar43 + (1'h1)))
        begin
          reg44 <= reg9[(5'h10):(2'h3)];
          reg45 <= $signed((({$unsigned(reg41)} != reg27) < (($signed(reg30) ?
              reg42[(1'h0):(1'h0)] : (+reg24)) != ((reg40 | reg7) | $unsigned(reg11)))));
          for (forvar46 = (1'h0); (forvar46 < (3'h4)); forvar46 = (forvar46 + (1'h1)))
            begin
              reg47 <= ((8'haa) ?
                  $signed(($signed(reg11) ?
                      ($signed(forvar43) ?
                          reg33 : reg39[(2'h3):(2'h3)]) : ($unsigned(forvar46) <<< reg23))) : forvar22);
              reg48 <= $unsigned(wire0);
            end
          reg49 <= {(^~$signed((~^(^~reg25))))};
        end
      for (forvar50 = (1'h0); (forvar50 < (1'h0)); forvar50 = (forvar50 + (1'h1)))
        begin
          reg51 <= (((|$unsigned((reg26 * reg26))) < reg38[(2'h3):(2'h2)]) ?
              ((wire19[(4'hb):(4'ha)] ?
                  (~^reg27) : $signed(reg30)) < reg10) : (($unsigned({reg12}) ^ forvar28[(3'h4):(1'h1)]) ?
                  $unsigned(reg45[(3'h7):(3'h6)]) : forvar46[(4'hb):(2'h2)]));
          reg52 <= forvar15;
        end
    end
  assign wire53 = $unsigned((!$signed(($unsigned(reg6) ?
                      $signed(forvar8) : $unsigned(reg24)))));
  assign wire54 = (~$signed(reg12[(2'h2):(1'h0)]));
  module55 modinst97 (wire96, clk, reg14, reg49, reg10, reg9, forvar22);
  assign wire98 = {reg11, {forvar22}};
  module99 modinst887 (.clk(clk), .wire103(forvar31), .wire100(reg51), .y(wire886), .wire101(wire2), .wire102(reg47), .wire104(reg14));
  assign wire888 = $signed(((({(8'ha9), reg13} ?
                           $signed(wire96) : ((8'hb4) ?
                               (8'h9e) : reg48)) != {reg44[(1'h0):(1'h0)],
                           $signed(wire96)}) ?
                       $unsigned((~^reg26)) : forvar22[(5'h10):(2'h2)]));
  always
    @(posedge clk) begin
      reg889 <= reg40[(4'hd):(3'h7)];
    end
  module890 modinst2679 (.wire891(forvar43), .wire893(reg36), .wire892(reg9), .y(wire2678), .wire894(wire98), .clk(clk));
  always
    @(posedge clk) begin
      reg2680 = (8'hb1);
      for (forvar2681 = (1'h0); (forvar2681 < (3'h4)); forvar2681 = (forvar2681 + (1'h1)))
        begin
          for (forvar2682 = (1'h0); (forvar2682 < (1'h1)); forvar2682 = (forvar2682 + (1'h1)))
            begin
              reg2683 <= reg47[(1'h0):(1'h0)];
            end
          reg2684 <= (8'ha3);
          reg2685 <= (((&$signed((wire98 > reg34))) == ($unsigned($unsigned(reg40)) + wire19[(3'h4):(2'h2)])) ?
              $signed(((|reg52[(4'hc):(2'h3)]) || $unsigned((reg25 ?
                  reg41 : reg45)))) : $unsigned(($unsigned((reg49 == forvar28)) ?
                  (~$unsigned(reg24)) : $signed((reg42 ? reg39 : wire0)))));
          for (forvar2686 = (1'h0); (forvar2686 < (2'h2)); forvar2686 = (forvar2686 + (1'h1)))
            begin
              reg2687 <= wire886;
              reg2688 <= (($unsigned(((reg17 ? (7'h40) : reg12) ?
                          (reg36 * reg13) : wire2678)) ?
                      $signed({((8'hb4) <<< forvar8)}) : ($signed($unsigned(reg27)) != (8'ha7))) ?
                  $signed($unsigned((|$signed((8'ha6))))) : $signed((~$signed(wire888))));
              reg2689 <= wire886[(3'h6):(3'h4)];
              reg2690 = reg6[(3'h4):(3'h4)];
            end
          reg2691 <= ({(|(reg18 ? (forvar22 ^ reg29) : $unsigned(forvar31))),
                  $signed((wire54[(3'h4):(2'h2)] ?
                      $unsigned(reg37) : forvar2681[(2'h2):(1'h1)]))} ?
              (~^reg14[(4'he):(4'hd)]) : reg7[(3'h5):(3'h4)]);
        end
      for (forvar2692 = (1'h0); (forvar2692 < (2'h2)); forvar2692 = (forvar2692 + (1'h1)))
        begin
          reg2693 = $unsigned((8'hb6));
          for (forvar2694 = (1'h0); (forvar2694 < (3'h4)); forvar2694 = (forvar2694 + (1'h1)))
            begin
              reg2695 = forvar2682[(4'hc):(3'h5)];
              reg2696 <= {wire2[(4'hb):(1'h1)]};
              reg2697 <= (8'h9c);
              reg2698 <= ((+reg2690[(4'hf):(4'hb)]) | reg13);
            end
          reg2699 <= $unsigned(($signed(($signed(reg26) | (reg30 && wire888))) ?
              $unsigned(($signed(reg52) < reg2691)) : $signed(reg2689)));
          for (forvar2700 = (1'h0); (forvar2700 < (2'h3)); forvar2700 = (forvar2700 + (1'h1)))
            begin
              reg2701 <= reg889[(3'h4):(2'h2)];
              reg2702 <= $unsigned($signed({$signed({wire98, (8'hbd)}),
                  reg32[(4'h9):(3'h5)]}));
              reg2703 = ((~|$signed(forvar2692)) ^ $signed((((reg27 << forvar2692) > reg2680) * {(~^(8'h9f)),
                  (8'hb0)})));
              reg2704 <= ((-$signed({(wire0 ? reg2701 : reg13),
                  $signed(reg2688)})) <<< (((^forvar15[(2'h2):(1'h1)]) < reg2698) ?
                  $signed(forvar2686) : reg52[(4'hb):(4'ha)]));
            end
        end
      reg2705 <= $signed(forvar2694);
      reg2706 = ((^($signed(reg40[(4'hf):(4'ha)]) ?
          $unsigned(reg27) : $unsigned((reg11 >> forvar2694)))) <<< $unsigned((|reg11[(5'h13):(2'h2)])));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module890
#( parameter param2676 = {({((8'ha1) ? ((8'had) != (7'h41)) : ((8'hb1) | (8'haf)))} && ((((7'h40) ? (8'hb4) : (8'hb3)) >>> {(8'hb3)}) > (((8'hbf) ? (8'h9c) : (8'hbd)) ^~ ((8'hab) ? (8'h9c) : (7'h43))))), (~^((((8'hbc) - (8'ha1)) ? ((8'hb3) ? (8'hbe) : (7'h44)) : {(8'hb3)}) ? ({(8'hb7), (7'h43)} <= {(8'had)}) : ((+(8'hb8)) ? {(8'hba)} : ((8'ha9) >>> (8'ha1)))))}
, parameter param2677 = (((param2676 ? ((~|param2676) <<< (|param2676)) : {param2676}) ? (|param2676) : (-(^param2676))) ? ((^{param2676}) != (((param2676 ? param2676 : param2676) >>> (param2676 ? param2676 : param2676)) && param2676)) : param2676) )
(y, clk, wire891, wire892, wire893, wire894);
  output wire [(32'h243):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire891;
  input wire signed [(5'h15):(1'h0)] wire892;
  input wire [(2'h3):(1'h0)] wire893;
  input wire signed [(5'h14):(1'h0)] wire894;
  reg [(5'h10):(1'h0)] reg2675 = (1'h0);
  wire [(4'ha):(1'h0)] wire2674;
  wire [(2'h3):(1'h0)] wire2673;
  reg signed [(5'h10):(1'h0)] reg2672 = (1'h0);
  reg [(5'h14):(1'h0)] reg2671 = (1'h0);
  reg [(5'h12):(1'h0)] reg2670 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2669 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2668 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2667 = (1'h0);
  reg [(5'h10):(1'h0)] forvar895 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg896 = (1'h0);
  reg [(5'h12):(1'h0)] reg897 = (1'h0);
  reg signed [(4'he):(1'h0)] reg898 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg899 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar900 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg901 = (1'h0);
  reg [(4'hf):(1'h0)] reg902 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg903 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar904 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg905 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1112;
  wire [(4'hc):(1'h0)] wire1114;
  reg signed [(4'hc):(1'h0)] reg1115 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1116 = (1'h0);
  reg [(3'h5):(1'h0)] reg1117 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1118 = (1'h0);
  wire [(5'h12):(1'h0)] wire1119;
  wire signed [(4'he):(1'h0)] wire1120;
  wire [(2'h2):(1'h0)] wire1121;
  wire [(4'ha):(1'h0)] wire1122;
  wire [(5'h10):(1'h0)] wire1123;
  reg signed [(2'h2):(1'h0)] reg1124 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1125 = (1'h0);
  reg [(5'h11):(1'h0)] reg1126 = (1'h0);
  reg [(4'hc):(1'h0)] reg1127 = (1'h0);
  reg [(5'h14):(1'h0)] reg1128 = (1'h0);
  reg [(5'h12):(1'h0)] reg1129 = (1'h0);
  wire [(5'h15):(1'h0)] wire1130;
  reg [(5'h13):(1'h0)] reg1131 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1132 = (1'h0);
  wire [(5'h14):(1'h0)] wire2665;
  assign y = {reg2675,
                 wire2674,
                 wire2673,
                 reg2672,
                 reg2671,
                 reg2670,
                 reg2669,
                 reg2668,
                 reg2667,
                 forvar895,
                 reg896,
                 reg897,
                 reg898,
                 reg899,
                 forvar900,
                 reg901,
                 reg902,
                 reg903,
                 forvar904,
                 reg905,
                 wire1112,
                 wire1114,
                 reg1115,
                 reg1116,
                 reg1117,
                 reg1118,
                 wire1119,
                 wire1120,
                 wire1121,
                 wire1122,
                 wire1123,
                 reg1124,
                 forvar1125,
                 reg1126,
                 reg1127,
                 reg1128,
                 reg1129,
                 wire1130,
                 reg1131,
                 reg1132,
                 wire2665,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar895 = (1'h0); (forvar895 < (3'h4)); forvar895 = (forvar895 + (1'h1)))
        begin
          reg896 = ({(~^$signed({wire891, (8'ha8)}))} ?
              wire894 : {($unsigned(wire891) ?
                      ($signed((8'hb6)) ?
                          (wire892 || wire893) : $signed(wire893)) : $unsigned(wire894[(1'h0):(1'h0)]))});
          reg897 <= ($signed({$signed((7'h42))}) < $signed((((reg896 ^ wire893) ~^ $signed(forvar895)) ?
              reg896[(5'h12):(5'h11)] : $unsigned(forvar895[(3'h7):(3'h6)]))));
        end
      reg898 <= reg896;
      reg899 <= ($unsigned($unsigned(wire892)) << reg897);
      for (forvar900 = (1'h0); (forvar900 < (1'h1)); forvar900 = (forvar900 + (1'h1)))
        begin
          reg901 <= $signed((~&$signed(reg898)));
          reg902 <= (&$signed(reg901[(2'h2):(1'h1)]));
          reg903 <= reg898[(4'he):(1'h0)];
        end
      for (forvar904 = (1'h0); (forvar904 < (1'h1)); forvar904 = (forvar904 + (1'h1)))
        begin
          reg905 <= (^~{(({(8'hb2)} + (&reg902)) ?
                  reg901 : wire894[(2'h2):(2'h2)]),
              (+forvar895)});
        end
    end
  module906 modinst1113 (.clk(clk), .wire909(forvar904), .y(wire1112), .wire910(reg896), .wire908(reg899), .wire907(reg902));
  assign wire1114 = $signed($signed($unsigned(((reg901 < reg899) >> forvar904[(1'h0):(1'h0)]))));
  always
    @(posedge clk) begin
      reg1115 <= (8'hbe);
      reg1116 <= $unsigned($signed((^~((wire892 != forvar895) ?
          (8'hbc) : $signed(reg903)))));
      reg1117 <= wire1114;
    end
  always
    @(posedge clk) begin
      reg1118 = reg1117;
    end
  assign wire1119 = $unsigned({($signed((wire892 && reg896)) >= forvar895),
                        reg898[(1'h1):(1'h1)]});
  assign wire1120 = ($unsigned(((+forvar895) ?
                        (~$unsigned(reg899)) : forvar895)) >> $unsigned((~|$signed($signed(reg1116)))));
  assign wire1121 = ((7'h40) ?
                        $unsigned(reg903[(3'h5):(2'h3)]) : wire892[(1'h1):(1'h1)]);
  assign wire1122 = forvar900[(1'h0):(1'h0)];
  assign wire1123 = ($signed((reg897 != ((^~reg1116) ?
                            wire1122[(1'h1):(1'h1)] : (~^reg905)))) ?
                        {{((wire1114 ? wire1114 : reg1118) ?
                                    (~(8'ha5)) : (reg1117 ?
                                        reg898 : wire891))}} : reg1115[(4'hc):(4'h9)]);
  always
    @(posedge clk) begin
      reg1124 = (~|(~&$unsigned($signed((forvar904 ? wire893 : reg896)))));
      for (forvar1125 = (1'h0); (forvar1125 < (2'h3)); forvar1125 = (forvar1125 + (1'h1)))
        begin
          reg1126 = (&(|$unsigned((~|{(8'had), wire1119}))));
          reg1127 = $signed($signed((!$unsigned($signed(reg905)))));
          reg1128 <= (+reg902[(4'h9):(3'h7)]);
          reg1129 <= $signed($signed(reg896[(4'hb):(3'h4)]));
        end
    end
  assign wire1130 = (($signed(wire1119[(4'hf):(4'hc)]) ?
                        ((|(reg1124 ? (8'hb7) : reg901)) ?
                            reg1117[(1'h0):(1'h0)] : reg898) : ($unsigned($unsigned(forvar895)) <= $signed(forvar904[(1'h1):(1'h1)]))) ~^ $signed($signed(reg1118[(3'h7):(3'h7)])));
  always
    @(posedge clk) begin
      reg1131 <= reg898;
      reg1132 <= {(^$signed((~&{reg899, (8'hbe)})))};
    end
  module1133 modinst2666 (wire2665, clk, wire1120, reg1129, reg1131, forvar1125, wire894);
  always
    @(posedge clk) begin
      reg2667 <= $unsigned($unsigned((wire1122 ?
          $unsigned({reg896}) : {$unsigned(wire1122), $signed(forvar895)})));
      if (wire1130[(3'h6):(3'h4)])
        begin
          reg2668 = ((($unsigned((|wire1119)) ?
                      (~^$signed(wire892)) : (-$unsigned(forvar895))) ?
                  (reg1116 >>> ($unsigned(reg1124) == $unsigned((8'hb5)))) : forvar900[(3'h5):(3'h4)]) ?
              $signed((($signed(wire2665) ?
                  (wire1123 ?
                      reg1126 : reg902) : $unsigned(wire1119)) - {(reg1126 == reg903),
                  reg896[(4'ha):(2'h3)]})) : ($signed(({reg1131} ?
                  $signed(wire891) : ((8'hb2) + wire893))) ~^ $unsigned((reg1129[(4'h9):(1'h0)] ?
                  (~|wire1123) : $unsigned(wire1120)))));
        end
      else
        begin
          reg2668 <= ((~&wire894[(1'h1):(1'h1)]) != wire891[(1'h1):(1'h0)]);
          reg2669 <= (8'haf);
          reg2670 = reg1132;
          reg2671 <= (7'h44);
          reg2672 <= (|$signed($unsigned((8'h9f))));
        end
    end
  assign wire2673 = wire1112[(1'h1):(1'h1)];
  assign wire2674 = wire1112[(3'h4):(1'h1)];
  always
    @(posedge clk) begin
      reg2675 = ($signed((($unsigned((8'hac)) != $signed(reg2667)) - ((forvar904 ?
              reg1126 : (7'h42)) + wire1123))) ?
          (($unsigned($signed(reg2672)) << (8'hb3)) ?
              $unsigned($signed(((8'ha3) > reg1116))) : wire1130[(2'h2):(1'h1)]) : ($signed(wire1122) && ((^(wire1112 ?
                  reg1118 : reg899)) ?
              $unsigned($unsigned(wire2673)) : $signed((8'h9f)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module99
#( parameter param884 = ((^((~|(^(8'hb6))) | (((8'hbb) ? (8'hbb) : (8'hb6)) ? ((8'ha4) ? (7'h42) : (8'hbe)) : ((7'h41) > (7'h42))))) ? (({(+(8'h9c))} ? (~^(^(8'hb6))) : (^(8'h9e))) ? ((|(^~(8'ha4))) ^ {(~^(8'hba))}) : (({(8'ha8)} ? (!(8'hb6)) : ((7'h43) ? (8'ha1) : (8'ha1))) & (~^((8'ha4) ^ (7'h41))))) : ((~((~(8'ha7)) ? ((8'ha6) ? (8'hb3) : (8'ha5)) : {(8'ha5), (8'ha8)})) || (((8'ha8) ? (~(8'hb3)) : (~^(8'hb4))) ? (^((7'h42) <= (8'hbc))) : ((~(8'h9d)) >= ((8'haf) ^ (8'hb7))))))
, parameter param885 = {(^~{((~^param884) ? param884 : (+param884))})} )
(y, clk, wire100, wire101, wire102, wire103, wire104);
  output wire [(32'h18a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire100;
  input wire [(4'hf):(1'h0)] wire101;
  input wire signed [(5'h15):(1'h0)] wire102;
  input wire signed [(4'h8):(1'h0)] wire103;
  input wire signed [(4'hc):(1'h0)] wire104;
  reg [(4'hc):(1'h0)] reg883 = (1'h0);
  reg signed [(4'he):(1'h0)] reg882 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg881 = (1'h0);
  reg [(4'hb):(1'h0)] reg880 = (1'h0);
  reg [(4'he):(1'h0)] forvar879 = (1'h0);
  reg [(4'hf):(1'h0)] reg878 = (1'h0);
  reg signed [(4'he):(1'h0)] reg877 = (1'h0);
  wire [(4'hd):(1'h0)] wire875;
  wire [(5'h15):(1'h0)] wire180;
  reg [(5'h14):(1'h0)] reg179 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg178 = (1'h0);
  reg [(4'hc):(1'h0)] reg177 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg176 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg175 = (1'h0);
  reg [(4'hf):(1'h0)] reg174 = (1'h0);
  reg [(5'h10):(1'h0)] forvar173 = (1'h0);
  wire [(4'h8):(1'h0)] wire172;
  wire [(4'h9):(1'h0)] wire105;
  wire [(5'h13):(1'h0)] wire106;
  wire signed [(4'hd):(1'h0)] wire107;
  reg [(5'h10):(1'h0)] reg108 = (1'h0);
  reg signed [(4'he):(1'h0)] reg109 = (1'h0);
  reg [(5'h12):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg111 = (1'h0);
  reg [(5'h10):(1'h0)] reg112 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg113 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg114 = (1'h0);
  wire [(5'h14):(1'h0)] wire170;
  assign y = {reg883,
                 reg882,
                 reg881,
                 reg880,
                 forvar879,
                 reg878,
                 reg877,
                 wire875,
                 wire180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 forvar173,
                 wire172,
                 wire105,
                 wire106,
                 wire107,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 reg112,
                 reg113,
                 reg114,
                 wire170,
                 (1'h0)};
  assign wire105 = wire104;
  assign wire106 = ($unsigned((|$signed(((8'ha1) >> wire101)))) ?
                       {$unsigned((-(wire104 < (8'hbf))))} : (~^$signed((8'ha5))));
  assign wire107 = (^wire101);
  always
    @(posedge clk) begin
      reg108 <= $unsigned($signed(wire102));
      reg109 <= {wire102};
    end
  always
    @(posedge clk) begin
      reg110 <= (+($unsigned($unsigned((reg108 + wire105))) >> (&$signed($signed((8'hb8))))));
      reg111 <= wire104[(4'hc):(4'hb)];
      reg112 <= $signed((($signed(wire106) ?
          {(reg111 ?
                  reg109 : wire103)} : {$signed(wire103)}) <<< (^~(~(&reg111)))));
      reg113 = wire104[(3'h4):(1'h0)];
      reg114 = {$signed(($unsigned({wire100}) ?
              reg110[(3'h4):(2'h2)] : $signed($unsigned(wire101))))};
    end
  module115 modinst171 (wire170, clk, reg114, reg110, wire100, reg111, reg109);
  assign wire172 = ($signed($signed(wire105[(1'h0):(1'h0)])) ^ $signed(($unsigned(reg108) ?
                       wire105 : reg108)));
  always
    @(posedge clk) begin
      for (forvar173 = (1'h0); (forvar173 < (3'h4)); forvar173 = (forvar173 + (1'h1)))
        begin
          reg174 = wire103[(4'h8):(1'h0)];
          reg175 <= (8'ha3);
          reg176 = $unsigned((^(reg108 != $unsigned(reg108[(3'h4):(3'h4)]))));
        end
    end
  always
    @(posedge clk) begin
      reg177 = (|(reg110[(2'h2):(1'h0)] ?
          (($unsigned((8'hbf)) & $unsigned(wire102)) == {wire102[(2'h2):(1'h1)]}) : ((~(wire104 ?
              reg110 : wire100)) * reg112[(3'h5):(2'h3)])));
      reg178 <= $unsigned((({$unsigned(reg112)} ?
          ((~&forvar173) ?
              reg108 : (wire100 ?
                  reg112 : reg176)) : $signed(wire102[(2'h2):(2'h2)])) << $signed($signed((forvar173 && reg175)))));
      reg179 <= wire172;
    end
  assign wire180 = $unsigned($unsigned($signed(reg178)));
  module181 modinst876 (.wire185(wire102), .clk(clk), .wire183(wire172), .wire184(reg112), .wire182(reg174), .y(wire875));
  always
    @(posedge clk) begin
      reg877 = $unsigned((reg110 ? wire100 : $unsigned(reg114[(3'h6):(3'h4)])));
      reg878 = (!wire180[(4'he):(4'hb)]);
      for (forvar879 = (1'h0); (forvar879 < (1'h0)); forvar879 = (forvar879 + (1'h1)))
        begin
          reg880 <= reg113[(3'h7):(3'h4)];
          reg881 = (+(^~(forvar879[(4'hb):(3'h7)] ?
              $unsigned($unsigned(wire102)) : (!wire172))));
          reg882 <= (~|reg108[(4'hb):(2'h2)]);
          reg883 <= ({((wire103 != (!wire875)) ?
                  reg179[(4'he):(1'h0)] : $signed(wire875)),
              reg178[(4'he):(2'h3)]} << $unsigned((wire106[(4'he):(4'ha)] ?
              wire170[(4'h9):(3'h4)] : (forvar173 ?
                  $unsigned(wire180) : (reg113 ? (8'haa) : wire101)))));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module55
#( parameter param94 = (7'h42)
, parameter param95 = ((param94 ? (param94 < param94) : (^~(^(^param94)))) == (~^((param94 >>> (!param94)) ? param94 : (~&(param94 >= param94))))) )
(y, clk, wire60, wire59, wire58, wire57, wire56);
  output wire [(32'h1a7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire60;
  input wire [(3'h7):(1'h0)] wire59;
  input wire signed [(5'h13):(1'h0)] wire58;
  input wire signed [(5'h12):(1'h0)] wire57;
  input wire signed [(5'h10):(1'h0)] wire56;
  wire [(2'h2):(1'h0)] wire93;
  reg [(4'h9):(1'h0)] reg92 = (1'h0);
  reg [(4'ha):(1'h0)] reg91 = (1'h0);
  reg [(5'h15):(1'h0)] reg90 = (1'h0);
  reg [(5'h15):(1'h0)] reg89 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar88 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg87 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg86 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg85 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg84 = (1'h0);
  reg [(5'h11):(1'h0)] reg83 = (1'h0);
  reg [(5'h12):(1'h0)] reg82 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar81 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg79 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar78 = (1'h0);
  reg [(3'h6):(1'h0)] reg77 = (1'h0);
  reg [(4'hd):(1'h0)] forvar76 = (1'h0);
  reg [(5'h14):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg74 = (1'h0);
  reg [(5'h14):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg72 = (1'h0);
  reg [(4'h8):(1'h0)] forvar71 = (1'h0);
  reg [(4'he):(1'h0)] reg70 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire69;
  reg [(3'h6):(1'h0)] reg68 = (1'h0);
  wire [(5'h12):(1'h0)] wire67;
  wire [(5'h12):(1'h0)] wire66;
  wire signed [(3'h6):(1'h0)] wire65;
  wire [(4'hf):(1'h0)] wire64;
  reg [(5'h11):(1'h0)] reg63 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg62 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg61 = (1'h0);
  assign y = {wire93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 forvar88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 forvar81,
                 reg80,
                 reg79,
                 forvar78,
                 reg77,
                 forvar76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 forvar71,
                 reg70,
                 wire69,
                 reg68,
                 wire67,
                 wire66,
                 wire65,
                 wire64,
                 reg63,
                 reg62,
                 reg61,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg61 <= (wire57 >> wire60);
      reg62 = wire56;
      reg63 <= $signed({$unsigned((reg61[(2'h2):(1'h1)] ?
              (~&wire59) : wire58[(3'h5):(1'h1)]))});
    end
  assign wire64 = $signed((reg61 >>> wire56[(3'h6):(1'h0)]));
  assign wire65 = (wire59 ?
                      {($unsigned(wire59) ?
                              ({wire57} ^ $unsigned(wire57)) : {$signed(wire56),
                                  $unsigned(wire57)})} : ((reg63[(2'h3):(2'h2)] || wire57) | (^~wire56)));
  assign wire66 = ((!(reg62[(3'h4):(1'h1)] ^~ ($unsigned(wire57) || $unsigned(wire58)))) << $signed(($unsigned(((8'hb8) >> (8'hbb))) < wire57[(4'he):(4'hb)])));
  assign wire67 = wire57;
  always
    @(posedge clk) begin
      reg68 <= (($unsigned(((~&wire58) ?
              $unsigned(wire59) : (reg61 ^ wire60))) ?
          (wire64[(4'ha):(1'h1)] ?
              ((wire65 ? wire57 : wire66) ?
                  wire57[(1'h1):(1'h1)] : (~|wire67)) : ((8'hb8) <<< {wire59})) : ((^{(8'hbe)}) <<< $unsigned((wire60 ~^ wire65)))) * {(~((wire64 >> wire57) ?
              (wire65 <<< reg63) : (reg61 ^ wire60)))});
    end
  assign wire69 = $signed($unsigned((((8'hbc) == $signed(wire57)) >>> $signed($unsigned(wire60)))));
  always
    @(posedge clk) begin
      reg70 <= {wire60[(4'hb):(4'h8)]};
      for (forvar71 = (1'h0); (forvar71 < (3'h4)); forvar71 = (forvar71 + (1'h1)))
        begin
          reg72 = reg61;
          reg73 <= $unsigned((&(wire58[(5'h12):(4'ha)] & ($signed(wire57) ?
              (wire67 ? reg68 : (8'ha8)) : (reg68 ? reg72 : wire59)))));
        end
    end
  always
    @(posedge clk) begin
      reg74 <= $unsigned($signed(((&(reg73 ?
          reg68 : wire69)) != wire64[(2'h3):(2'h3)])));
      reg75 <= (8'hb1);
      for (forvar76 = (1'h0); (forvar76 < (3'h4)); forvar76 = (forvar76 + (1'h1)))
        begin
          reg77 <= reg63;
        end
      for (forvar78 = (1'h0); (forvar78 < (3'h4)); forvar78 = (forvar78 + (1'h1)))
        begin
          reg79 <= $signed((~(&(!wire64[(3'h6):(3'h5)]))));
          reg80 <= (($signed({$signed(reg73), (reg63 ? (8'ha0) : (8'ha4))}) ?
              $signed(wire67[(4'he):(1'h0)]) : (7'h42)) != (8'h9f));
          for (forvar81 = (1'h0); (forvar81 < (3'h4)); forvar81 = (forvar81 + (1'h1)))
            begin
              reg82 = {{(+($signed(reg72) >>> (wire56 * (8'ha4)))),
                      wire59[(3'h4):(1'h0)]}};
              reg83 = {reg80};
              reg84 <= {(reg77 != wire66[(4'hb):(4'h9)])};
              reg85 <= (~|$signed(reg77[(1'h1):(1'h0)]));
              reg86 <= ($unsigned({(8'hb9),
                      {(reg82 ? (8'ha7) : reg68), (-wire60)}}) ?
                  (~{reg75[(1'h1):(1'h0)]}) : {(~$signed($signed(reg68))),
                      (($signed(reg84) ?
                              ((8'haa) ?
                                  (8'hb3) : wire60) : (forvar78 << reg70)) ?
                          reg79 : ((&wire57) ?
                              (wire59 || (8'haf)) : reg84[(3'h4):(1'h0)]))});
            end
          reg87 = ((wire64[(4'hb):(3'h4)] >> (((reg68 ?
                  reg73 : forvar81) << reg62) << $signed($signed((8'h9f))))) ?
              {($signed($unsigned(reg62)) ^ $signed({reg77})),
                  reg61[(2'h3):(1'h1)]} : $signed((&(7'h40))));
          for (forvar88 = (1'h0); (forvar88 < (1'h1)); forvar88 = (forvar88 + (1'h1)))
            begin
              reg89 <= (reg80[(2'h2):(1'h0)] ?
                  (($unsigned((reg74 - forvar78)) - (-(forvar71 | reg77))) | $signed($signed({wire59,
                      wire57}))) : $signed(reg75));
              reg90 = $signed((!$signed((reg73 ?
                  reg89[(3'h4):(1'h0)] : (wire65 && reg87)))));
              reg91 <= (8'ha1);
            end
        end
      reg92 <= $signed(reg85[(2'h2):(1'h1)]);
    end
  assign wire93 = wire56[(4'h8):(4'h8)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module181
#( parameter param873 = ({(!{{(8'ha2), (8'ha3)}})} ? {((((8'hac) != (8'hb4)) >> (-(8'ha0))) <<< (((8'ha8) <= (8'hbd)) ? (-(8'hae)) : ((8'haa) + (8'ha6))))} : (^(|((+(8'haa)) ? (8'ha3) : ((8'h9d) ? (8'hb8) : (8'ha2))))))
, parameter param874 = ((&((param873 < (param873 >> param873)) ? ((|param873) ? (-param873) : (param873 ^~ param873)) : {(-param873)})) || (~|param873)) )
(y, clk, wire182, wire183, wire184, wire185);
  output wire [(32'h7f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire182;
  input wire signed [(4'h8):(1'h0)] wire183;
  input wire signed [(4'h8):(1'h0)] wire184;
  input wire [(5'h15):(1'h0)] wire185;
  wire signed [(4'h8):(1'h0)] wire872;
  wire [(5'h11):(1'h0)] wire186;
  wire signed [(4'hd):(1'h0)] wire187;
  reg [(5'h13):(1'h0)] reg188 = (1'h0);
  reg signed [(4'he):(1'h0)] reg189 = (1'h0);
  wire [(5'h13):(1'h0)] wire190;
  wire signed [(5'h12):(1'h0)] wire191;
  wire [(5'h12):(1'h0)] wire870;
  assign y = {wire872,
                 wire186,
                 wire187,
                 reg188,
                 reg189,
                 wire190,
                 wire191,
                 wire870,
                 (1'h0)};
  assign wire186 = $signed(wire183);
  assign wire187 = wire182;
  always
    @(posedge clk) begin
      reg188 = wire185;
      reg189 <= {wire186};
    end
  assign wire190 = ($signed((8'ha7)) >>> (((|(8'ha1)) <= {(wire184 || wire183)}) ?
                       wire182[(3'h5):(1'h0)] : ($unsigned($unsigned(wire186)) - $signed(((8'ha5) || wire183)))));
  assign wire191 = {(8'ha1), $unsigned($signed((~&wire182)))};
  module192 modinst871 (.wire195(reg188), .clk(clk), .wire196(wire186), .y(wire870), .wire197(wire190), .wire194(wire185), .wire193(wire187));
  assign wire872 = $signed($unsigned({((+wire185) - (8'hbd)),
                       (-(wire182 >> wire186))}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module115
#( parameter param169 = (|{(|(((8'hbe) ? (8'hbb) : (8'haa)) ? ((8'hbe) ? (8'had) : (8'hb5)) : ((8'hbc) ? (8'hba) : (8'hbe)))), (&{(^~(8'haa)), ((8'ha1) ? (8'hb3) : (8'hab))})}) )
(y, clk, wire120, wire119, wire118, wire117, wire116);
  output wire [(32'h23c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire120;
  input wire signed [(5'h12):(1'h0)] wire119;
  input wire signed [(5'h12):(1'h0)] wire118;
  input wire [(5'h15):(1'h0)] wire117;
  input wire [(4'he):(1'h0)] wire116;
  reg signed [(5'h10):(1'h0)] reg168 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg167 = (1'h0);
  reg [(5'h14):(1'h0)] reg166 = (1'h0);
  reg [(5'h14):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg164 = (1'h0);
  reg [(5'h11):(1'h0)] reg157 = (1'h0);
  reg [(3'h7):(1'h0)] reg163 = (1'h0);
  reg [(3'h6):(1'h0)] reg162 = (1'h0);
  reg [(3'h5):(1'h0)] reg161 = (1'h0);
  reg [(4'hf):(1'h0)] reg160 = (1'h0);
  reg signed [(4'he):(1'h0)] reg159 = (1'h0);
  reg [(4'h8):(1'h0)] reg158 = (1'h0);
  reg [(4'h9):(1'h0)] forvar157 = (1'h0);
  reg [(5'h14):(1'h0)] reg156 = (1'h0);
  wire [(3'h5):(1'h0)] wire155;
  reg [(4'hc):(1'h0)] reg154 = (1'h0);
  reg [(5'h11):(1'h0)] reg153 = (1'h0);
  reg [(5'h15):(1'h0)] reg152 = (1'h0);
  reg [(5'h15):(1'h0)] forvar151 = (1'h0);
  wire [(3'h4):(1'h0)] wire150;
  reg [(4'hd):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg148 = (1'h0);
  reg [(2'h3):(1'h0)] reg147 = (1'h0);
  reg [(4'ha):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg145 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg144 = (1'h0);
  reg [(5'h12):(1'h0)] forvar143 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire142;
  wire [(3'h6):(1'h0)] wire141;
  reg [(4'he):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg139 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg138 = (1'h0);
  reg [(3'h5):(1'h0)] reg137 = (1'h0);
  reg [(4'h9):(1'h0)] reg136 = (1'h0);
  reg [(5'h15):(1'h0)] reg135 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire134;
  reg [(5'h12):(1'h0)] reg133 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg132 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg131 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg129 = (1'h0);
  reg [(2'h2):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar127 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg126 = (1'h0);
  reg [(3'h4):(1'h0)] forvar125 = (1'h0);
  reg [(2'h2):(1'h0)] reg124 = (1'h0);
  reg [(5'h10):(1'h0)] reg123 = (1'h0);
  reg [(3'h4):(1'h0)] forvar122 = (1'h0);
  reg [(5'h10):(1'h0)] reg121 = (1'h0);
  assign y = {reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg157,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 forvar157,
                 reg156,
                 wire155,
                 reg154,
                 reg153,
                 reg152,
                 forvar151,
                 wire150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 forvar143,
                 wire142,
                 wire141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 wire134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 forvar127,
                 reg126,
                 forvar125,
                 reg124,
                 reg123,
                 forvar122,
                 reg121,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg121 <= $unsigned($unsigned($signed(wire116[(1'h1):(1'h1)])));
      for (forvar122 = (1'h0); (forvar122 < (3'h4)); forvar122 = (forvar122 + (1'h1)))
        begin
          reg123 <= ($signed({((reg121 ? wire116 : wire118) ?
                  (wire116 | (8'ha1)) : (-(8'haf))),
              ($unsigned((8'hba)) > (|forvar122))}) | reg121[(3'h4):(2'h3)]);
        end
      reg124 = {$unsigned(($unsigned(wire119) ?
              ((wire120 >> reg123) >= $signed(wire118)) : reg123[(2'h3):(2'h3)])),
          $signed($signed(($signed(wire118) ? $unsigned(wire117) : wire118)))};
      for (forvar125 = (1'h0); (forvar125 < (3'h4)); forvar125 = (forvar125 + (1'h1)))
        begin
          reg126 <= $signed(wire119[(2'h3):(1'h1)]);
          for (forvar127 = (1'h0); (forvar127 < (2'h2)); forvar127 = (forvar127 + (1'h1)))
            begin
              reg128 = $unsigned({$unsigned(forvar125[(2'h3):(2'h3)]),
                  $unsigned((forvar122[(2'h2):(1'h0)] ?
                      forvar125[(1'h1):(1'h1)] : $signed((8'ha8))))});
              reg129 <= forvar127;
            end
          if ((($unsigned($signed($signed(reg129))) ?
                  {($unsigned((8'hbf)) & wire119)} : reg128[(1'h0):(1'h0)]) ?
              reg129 : forvar125))
            begin
              reg130 <= $signed(wire119);
              reg131 = ({((wire116[(2'h3):(1'h0)] - reg121) >>> {$signed(wire119),
                          forvar122[(2'h3):(1'h1)]}),
                      (($signed(forvar127) ?
                          $unsigned(reg126) : {reg124,
                              wire117}) >= {$signed(wire117),
                          forvar125[(1'h1):(1'h1)]})} ?
                  $signed($signed((~&{reg124,
                      forvar125}))) : $unsigned({$unsigned(reg129[(4'hd):(3'h4)])}));
              reg132 <= wire117[(4'he):(3'h7)];
            end
          else
            begin
              reg130 <= $unsigned((((!((7'h40) ? reg132 : wire118)) ?
                      ({reg129} ?
                          reg126[(2'h3):(2'h2)] : (reg126 ?
                              wire117 : reg130)) : $unsigned(reg126[(4'hb):(3'h6)])) ?
                  $unsigned(reg132) : (8'hac)));
              reg131 <= ($unsigned(wire120) ^ $unsigned($unsigned($signed($signed(reg126)))));
              reg132 = (~forvar122);
            end
        end
      reg133 <= reg123;
    end
  assign wire134 = wire116[(4'h8):(1'h0)];
  always
    @(posedge clk) begin
      reg135 <= reg123[(2'h3):(2'h2)];
      reg136 <= reg131;
    end
  always
    @(posedge clk) begin
      reg137 <= {$unsigned((&$signed(reg135[(4'hc):(2'h3)]))),
          $signed(wire118[(2'h3):(1'h0)])};
      reg138 <= $signed(((((reg132 ? reg129 : reg123) ?
              (^(8'hb0)) : (-forvar125)) ?
          $signed(((8'ha4) && (7'h41))) : {{wire134},
              (7'h44)}) <= $signed(($signed(reg129) ?
          $unsigned((8'ha2)) : $signed(reg135)))));
      reg139 <= reg136[(4'h8):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg140 = {(reg135 ? $unsigned(wire117[(4'hc):(3'h5)]) : reg123)};
    end
  assign wire141 = wire119[(5'h12):(1'h1)];
  assign wire142 = $signed($signed($signed((!(reg121 ? reg140 : wire117)))));
  always
    @(posedge clk) begin
      for (forvar143 = (1'h0); (forvar143 < (1'h0)); forvar143 = (forvar143 + (1'h1)))
        begin
          reg144 <= (forvar127[(3'h6):(3'h6)] ?
              forvar125[(1'h1):(1'h0)] : $unsigned((-$signed((reg133 >> forvar143)))));
          reg145 = $signed($signed((^($unsigned((7'h43)) ?
              ((8'haf) > wire142) : reg137))));
          reg146 <= ($signed($signed(reg133)) ?
              $unsigned((((8'h9d) || $signed(reg133)) ?
                  $unsigned($signed((8'hb6))) : $signed((reg130 - reg137)))) : $unsigned((($unsigned((8'hba)) < $unsigned((8'hb5))) == (!reg133))));
          reg147 <= reg135[(3'h5):(2'h3)];
          reg148 <= forvar122[(3'h4):(2'h3)];
        end
      reg149 <= $signed($signed($unsigned({{reg139},
          (reg148 ? (8'hac) : reg144)})));
    end
  assign wire150 = ($signed(({(&reg137),
                       reg149[(3'h4):(1'h0)]} && (~wire119))) >= (-$signed(({reg148} <<< (reg129 > (8'hb0))))));
  always
    @(posedge clk) begin
      for (forvar151 = (1'h0); (forvar151 < (2'h3)); forvar151 = (forvar151 + (1'h1)))
        begin
          reg152 <= ((+wire118[(4'hb):(4'hb)]) ?
              (forvar125[(2'h2):(1'h0)] != wire120[(2'h3):(2'h3)]) : (~^(&$signed(reg131[(4'hc):(4'h9)]))));
          reg153 <= (~$unsigned((reg146 ?
              $signed($unsigned(reg138)) : $unsigned($signed(reg128)))));
          reg154 = $signed($unsigned(($unsigned((^wire117)) ?
              (((8'had) ?
                  reg128 : forvar125) ^~ $unsigned(reg123)) : (reg131[(5'h10):(4'hc)] << (~|reg152)))));
        end
    end
  assign wire155 = wire120[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      reg156 <= reg131[(5'h11):(4'ha)];
      if (({(!{$signed(reg121)}), $unsigned($unsigned(reg124))} ?
          wire116 : reg139))
        begin
          for (forvar157 = (1'h0); (forvar157 < (2'h3)); forvar157 = (forvar157 + (1'h1)))
            begin
              reg158 = (|$unsigned(reg146[(2'h2):(1'h0)]));
              reg159 = $signed($signed(((~|reg145[(2'h2):(2'h2)]) ?
                  (reg137[(2'h3):(1'h1)] | $signed(wire117)) : ($unsigned(reg132) ?
                      $unsigned((8'hae)) : wire116[(1'h1):(1'h0)]))));
              reg160 = ($signed({forvar127[(2'h3):(1'h0)]}) != (reg140 ?
                  (~|(~^(8'hac))) : (~&(reg138 ?
                      wire116[(4'hc):(4'ha)] : (reg146 ? reg136 : reg147)))));
              reg161 <= reg124;
            end
          reg162 <= (^~reg123);
          reg163 <= {reg138[(2'h3):(2'h2)], (~&reg138)};
        end
      else
        begin
          reg157 = forvar127[(5'h11):(2'h2)];
          reg158 <= forvar157;
        end
      reg164 <= wire119;
      reg165 = $unsigned(((({wire117} ^ (reg156 ?
              reg152 : (7'h40))) > (reg158[(4'h8):(1'h0)] >= (reg136 ?
              reg136 : reg136))) ?
          $unsigned((wire134 ?
              $unsigned(reg153) : $signed(wire155))) : (forvar122[(1'h0):(1'h0)] ?
              reg162[(1'h0):(1'h0)] : ((reg121 ?
                  reg153 : (8'hb2)) > (forvar157 ? reg123 : reg121)))));
      reg166 = $signed(reg128[(1'h1):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg167 <= reg138[(2'h2):(1'h1)];
      reg168 <= reg123;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module192
#( parameter param868 = {(8'ha3), ((^~{(8'hbf), ((8'ha6) && (8'hbc))}) ? (^(~^(&(8'ha0)))) : ((8'ha8) ^ (((8'hb4) - (8'haa)) ? {(7'h44), (7'h40)} : ((8'h9c) <<< (8'hba)))))}
, parameter param869 = (+((^~((~&param868) ? (param868 ? param868 : param868) : (param868 | param868))) & (&{param868, (~&param868)}))) )
(y, clk, wire193, wire194, wire195, wire196, wire197);
  output wire [(32'h24f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire193;
  input wire signed [(5'h15):(1'h0)] wire194;
  input wire [(5'h13):(1'h0)] wire195;
  input wire signed [(5'h11):(1'h0)] wire196;
  input wire signed [(5'h13):(1'h0)] wire197;
  wire signed [(3'h5):(1'h0)] wire866;
  reg [(4'hf):(1'h0)] reg745 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg744 = (1'h0);
  reg [(2'h3):(1'h0)] reg743 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg742 = (1'h0);
  reg [(4'h9):(1'h0)] reg741 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar740 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg739 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg738 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg737 = (1'h0);
  reg [(5'h10):(1'h0)] reg736 = (1'h0);
  reg [(5'h10):(1'h0)] forvar735 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg734 = (1'h0);
  reg [(3'h7):(1'h0)] forvar733 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg732 = (1'h0);
  reg [(5'h12):(1'h0)] reg731 = (1'h0);
  reg [(4'hd):(1'h0)] reg730 = (1'h0);
  wire signed [(4'he):(1'h0)] wire729;
  wire [(5'h12):(1'h0)] wire728;
  reg signed [(3'h5):(1'h0)] reg727 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg726 = (1'h0);
  reg [(4'h8):(1'h0)] reg725 = (1'h0);
  wire [(5'h14):(1'h0)] wire724;
  reg [(4'ha):(1'h0)] reg723 = (1'h0);
  reg [(5'h15):(1'h0)] reg722 = (1'h0);
  wire signed [(4'he):(1'h0)] wire720;
  wire [(3'h6):(1'h0)] wire198;
  reg [(5'h10):(1'h0)] reg199 = (1'h0);
  reg [(5'h12):(1'h0)] reg200 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg201 = (1'h0);
  wire [(5'h10):(1'h0)] wire499;
  reg [(3'h4):(1'h0)] reg501 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire502;
  reg signed [(5'h10):(1'h0)] reg503 = (1'h0);
  reg [(4'hc):(1'h0)] forvar504 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg505 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg506 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg507 = (1'h0);
  reg [(3'h5):(1'h0)] forvar508 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg509 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar511 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg512 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg513 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg514 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg515 = (1'h0);
  wire [(4'ha):(1'h0)] wire611;
  assign y = {wire866,
                 reg745,
                 reg744,
                 reg743,
                 reg742,
                 reg741,
                 forvar740,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 forvar735,
                 reg734,
                 forvar733,
                 reg732,
                 reg731,
                 reg730,
                 wire729,
                 wire728,
                 reg727,
                 reg726,
                 reg725,
                 wire724,
                 reg723,
                 reg722,
                 wire720,
                 wire198,
                 reg199,
                 reg200,
                 reg201,
                 wire499,
                 reg501,
                 wire502,
                 reg503,
                 forvar504,
                 reg505,
                 reg506,
                 reg507,
                 forvar508,
                 reg509,
                 reg510,
                 forvar511,
                 reg512,
                 reg513,
                 reg514,
                 reg515,
                 wire611,
                 (1'h0)};
  assign wire198 = ((!{(!$signed(wire195)),
                       wire195[(2'h2):(1'h0)]}) & ((wire194[(5'h11):(4'ha)] ?
                           (wire195[(3'h6):(3'h5)] ?
                               (^~wire196) : (wire194 ?
                                   wire194 : wire193)) : wire193[(4'ha):(3'h7)]) ?
                       $signed($signed((wire197 ?
                           wire197 : wire196))) : wire193));
  always
    @(posedge clk) begin
      reg199 <= wire197[(3'h7):(3'h6)];
      reg200 = wire196;
      reg201 <= $signed($unsigned((~&({(7'h43)} ?
          $signed((8'hab)) : (wire193 * wire198)))));
    end
  module202 modinst500 (wire499, clk, reg200, wire193, wire195, wire194);
  always
    @(posedge clk) begin
      reg501 <= (($signed(($signed((7'h43)) ?
              (wire194 ~^ wire197) : (wire193 ? wire193 : wire499))) ?
          wire197 : {$signed(wire194[(5'h11):(3'h5)])}) < {(^~(^~wire197))});
    end
  assign wire502 = reg201[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg503 <= (~^wire502);
      for (forvar504 = (1'h0); (forvar504 < (3'h4)); forvar504 = (forvar504 + (1'h1)))
        begin
          reg505 = $unsigned(($unsigned((&(reg501 << wire196))) ?
              wire193 : wire502[(5'h14):(4'hf)]));
          reg506 <= reg501;
          reg507 <= ((reg201[(2'h3):(1'h1)] ?
                  $unsigned(((wire194 && reg501) ?
                      (wire195 || reg201) : $unsigned(wire499))) : (~(8'hba))) ?
              (~|reg201[(2'h3):(2'h2)]) : ((~wire194) + $signed(wire502)));
        end
      for (forvar508 = (1'h0); (forvar508 < (2'h3)); forvar508 = (forvar508 + (1'h1)))
        begin
          reg509 <= wire198[(2'h2):(2'h2)];
          reg510 <= $signed({($unsigned({(7'h41),
                  reg200}) << ((~wire196) ~^ {reg501})),
              wire193[(4'ha):(1'h1)]});
          for (forvar511 = (1'h0); (forvar511 < (1'h1)); forvar511 = (forvar511 + (1'h1)))
            begin
              reg512 <= reg506;
              reg513 <= $unsigned(forvar511);
            end
          reg514 = reg201;
        end
      reg515 <= $unsigned(wire193);
    end
  module516 modinst612 (wire611, clk, reg503, reg514, reg509, wire499, wire193);
  module613 modinst721 (.wire617(reg200), .wire616(wire499), .y(wire720), .wire615(forvar511), .clk(clk), .wire614(reg509));
  always
    @(posedge clk) begin
      reg722 <= $unsigned(reg510[(4'hc):(4'hc)]);
      reg723 <= reg509;
    end
  assign wire724 = (|$signed((~|$unsigned((wire193 ? wire195 : reg512)))));
  always
    @(posedge clk) begin
      reg725 = wire611[(3'h5):(3'h5)];
      reg726 = (8'h9f);
      reg727 <= (reg200 ? reg726[(2'h3):(1'h1)] : forvar511[(3'h4):(1'h0)]);
    end
  assign wire728 = reg514;
  assign wire729 = $unsigned(reg507[(3'h7):(2'h3)]);
  always
    @(posedge clk) begin
      reg730 = (wire197[(1'h1):(1'h1)] ?
          ($signed({((8'ha5) & reg510)}) ?
              (reg501 << ($signed(reg200) <<< forvar508)) : reg505) : ({(~^forvar504),
              $unsigned($signed(reg510))} * (($unsigned((8'ha9)) ?
                  wire196 : (8'haf)) ?
              (forvar508 != $signed(reg201)) : ($signed(wire502) ?
                  $signed((8'hbf)) : reg515[(1'h1):(1'h1)]))));
      reg731 <= $signed($signed(($signed(reg727[(1'h0):(1'h0)]) == $signed($signed(reg513)))));
      reg732 <= $unsigned($signed((-({reg506, reg512} ?
          $signed(reg200) : (reg730 ? wire611 : wire502)))));
      for (forvar733 = (1'h0); (forvar733 < (2'h3)); forvar733 = (forvar733 + (1'h1)))
        begin
          reg734 = $unsigned($unsigned($signed(wire499)));
          for (forvar735 = (1'h0); (forvar735 < (2'h3)); forvar735 = (forvar735 + (1'h1)))
            begin
              reg736 <= (8'ha0);
              reg737 <= $signed({(8'h9f), (^~reg200)});
              reg738 <= reg514[(1'h1):(1'h0)];
              reg739 = (($unsigned($signed(forvar733[(2'h2):(2'h2)])) << {(((8'had) != wire724) ?
                      $signed((8'hbb)) : (-reg736)),
                  reg722[(1'h1):(1'h1)]}) | $signed($unsigned((reg514[(1'h1):(1'h0)] - (reg515 << reg503)))));
            end
        end
      for (forvar740 = (1'h0); (forvar740 < (1'h1)); forvar740 = (forvar740 + (1'h1)))
        begin
          reg741 <= ($unsigned(wire724) <<< ((-$signed((-wire729))) > reg515));
          reg742 <= reg722;
          reg743 <= ((forvar511 ?
                  (($unsigned(reg515) >= (reg730 <<< wire194)) > {forvar740[(4'h9):(4'h9)]}) : wire724) ?
              $signed((~^$signed(reg739[(2'h2):(1'h1)]))) : $signed(wire502[(5'h10):(4'h9)]));
          reg744 <= $unsigned((wire196[(4'ha):(2'h2)] ?
              reg201[(2'h3):(1'h1)] : $signed($signed(wire728[(4'hf):(1'h1)]))));
          reg745 <= ((-$unsigned(($signed(reg738) ?
              $signed(reg199) : (reg201 ?
                  reg201 : (8'h9c))))) - $unsigned(wire499[(4'h9):(4'h8)]));
        end
    end
  module746 modinst867 (.wire748(wire193), .wire750(reg731), .wire747(reg503), .clk(clk), .wire749(reg722), .y(wire866));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module746
#( parameter param865 = (^~{({(|(8'ha8)), ((7'h44) ? (8'hbd) : (7'h42))} < {{(8'hb2)}, ((8'hbc) ? (8'haa) : (8'ha1))}), {{((8'h9c) ? (8'ha2) : (8'h9c)), ((8'ha4) <= (8'hb8))}, ((^(8'haf)) ? (^(8'ha6)) : (8'haf))}}) )
(y, clk, wire747, wire748, wire749, wire750);
  output wire [(32'h2e6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire747;
  input wire [(4'hd):(1'h0)] wire748;
  input wire signed [(5'h15):(1'h0)] wire749;
  input wire signed [(5'h11):(1'h0)] wire750;
  reg [(4'he):(1'h0)] reg864 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg863 = (1'h0);
  reg [(3'h6):(1'h0)] reg862 = (1'h0);
  reg [(4'ha):(1'h0)] reg861 = (1'h0);
  reg signed [(4'he):(1'h0)] reg860 = (1'h0);
  reg [(3'h4):(1'h0)] forvar859 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg858 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg857 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg856 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg855 = (1'h0);
  reg [(3'h4):(1'h0)] reg854 = (1'h0);
  reg [(4'h9):(1'h0)] reg853 = (1'h0);
  reg [(5'h15):(1'h0)] forvar852 = (1'h0);
  reg [(4'h9):(1'h0)] reg851 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire850;
  reg signed [(5'h15):(1'h0)] reg849 = (1'h0);
  reg [(5'h13):(1'h0)] reg848 = (1'h0);
  reg [(5'h15):(1'h0)] reg847 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg846 = (1'h0);
  reg [(4'hd):(1'h0)] reg845 = (1'h0);
  reg [(5'h12):(1'h0)] forvar844 = (1'h0);
  reg [(4'hc):(1'h0)] reg843 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg842 = (1'h0);
  reg [(2'h3):(1'h0)] reg751 = (1'h0);
  reg [(3'h7):(1'h0)] reg752 = (1'h0);
  wire [(4'hb):(1'h0)] wire753;
  wire [(4'ha):(1'h0)] wire754;
  wire [(4'hb):(1'h0)] wire755;
  wire [(4'hd):(1'h0)] wire756;
  reg signed [(5'h14):(1'h0)] reg757 = (1'h0);
  reg [(5'h14):(1'h0)] reg758 = (1'h0);
  reg [(4'h9):(1'h0)] reg759 = (1'h0);
  reg [(3'h7):(1'h0)] reg760 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg761 = (1'h0);
  reg [(4'hf):(1'h0)] reg762 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg763 = (1'h0);
  reg [(5'h14):(1'h0)] reg764 = (1'h0);
  reg [(5'h11):(1'h0)] reg765 = (1'h0);
  reg [(3'h7):(1'h0)] reg766 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg767 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg768 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg769 = (1'h0);
  reg signed [(4'he):(1'h0)] reg770 = (1'h0);
  reg [(3'h4):(1'h0)] forvar771 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar772 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg773 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg774 = (1'h0);
  reg [(5'h10):(1'h0)] reg775 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg776 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg777 = (1'h0);
  reg [(3'h6):(1'h0)] reg778 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg779 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg780 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg781 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar782 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg783 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg784 = (1'h0);
  reg signed [(4'he):(1'h0)] reg785 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg786 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar779 = (1'h0);
  reg [(2'h3):(1'h0)] reg782 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg787 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire840;
  assign y = {reg864,
                 reg863,
                 reg862,
                 reg861,
                 reg860,
                 forvar859,
                 reg858,
                 reg857,
                 reg856,
                 reg855,
                 reg854,
                 reg853,
                 forvar852,
                 reg851,
                 wire850,
                 reg849,
                 reg848,
                 reg847,
                 reg846,
                 reg845,
                 forvar844,
                 reg843,
                 reg842,
                 reg751,
                 reg752,
                 wire753,
                 wire754,
                 wire755,
                 wire756,
                 reg757,
                 reg758,
                 reg759,
                 reg760,
                 reg761,
                 reg762,
                 reg763,
                 reg764,
                 reg765,
                 reg766,
                 reg767,
                 reg768,
                 reg769,
                 reg770,
                 forvar771,
                 forvar772,
                 reg773,
                 reg774,
                 reg775,
                 reg776,
                 reg777,
                 reg778,
                 reg779,
                 reg780,
                 reg781,
                 forvar782,
                 reg783,
                 reg784,
                 reg785,
                 reg786,
                 forvar779,
                 reg782,
                 reg787,
                 wire840,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg751 <= $signed($unsigned($signed(wire748)));
      reg752 <= wire748[(3'h5):(2'h3)];
    end
  assign wire753 = (~|((($signed(wire749) ?
                           $unsigned((7'h41)) : $signed((8'had))) + (~^(reg751 ~^ wire749))) ?
                       $signed({(wire750 >> wire747),
                           wire750[(5'h11):(2'h3)]}) : wire747[(3'h5):(2'h2)]));
  assign wire754 = $signed((~&wire749));
  assign wire755 = reg751;
  assign wire756 = $signed(wire754);
  always
    @(posedge clk) begin
      reg757 <= {((8'hbb) ?
              $signed(reg751[(1'h1):(1'h0)]) : $signed(wire755[(3'h4):(3'h4)])),
          $unsigned({(~^$signed(wire754)),
              $unsigned((wire755 ? wire754 : wire749))})};
      reg758 <= wire756[(2'h3):(1'h1)];
      reg759 = (!wire748);
      reg760 <= wire749;
      reg761 = $signed((~((&{wire755, (7'h44)}) ?
          ((reg751 ^ wire754) ?
              $unsigned(wire756) : {wire747}) : reg751[(1'h1):(1'h1)])));
    end
  always
    @(posedge clk) begin
      reg762 <= ($signed($unsigned(wire750[(3'h4):(3'h4)])) + {{$signed($signed(reg751)),
              $unsigned(wire756[(4'hb):(4'h9)])}});
      reg763 <= (~reg761);
      reg764 <= (8'ha4);
      reg765 <= {(^~$unsigned(reg752))};
      reg766 <= reg758;
    end
  always
    @(posedge clk) begin
      reg767 <= reg759[(4'h8):(1'h1)];
      reg768 = $unsigned((reg762[(4'h8):(1'h1)] && reg763[(3'h4):(2'h2)]));
    end
  always
    @(posedge clk) begin
      reg769 <= $signed({$unsigned(((&(8'hb3)) ?
              reg764[(5'h10):(4'hf)] : (~&wire753))),
          reg758[(5'h10):(3'h6)]});
    end
  always
    @(posedge clk) begin
      reg770 <= $signed(((reg764[(5'h10):(4'hd)] ?
          (8'ha1) : $unsigned(reg762[(4'ha):(2'h2)])) ^~ reg762));
      for (forvar771 = (1'h0); (forvar771 < (1'h0)); forvar771 = (forvar771 + (1'h1)))
        begin
          for (forvar772 = (1'h0); (forvar772 < (3'h4)); forvar772 = (forvar772 + (1'h1)))
            begin
              reg773 = (7'h42);
              reg774 <= wire747;
              reg775 <= reg751[(2'h2):(1'h0)];
              reg776 <= (~|$unsigned(wire750));
              reg777 <= reg773;
            end
        end
      reg778 = reg757;
      if ((((((!reg758) ? (reg760 << reg774) : {reg776, (8'hb7)}) ?
          reg751[(2'h2):(1'h1)] : ($signed(reg773) ?
              (reg751 | reg759) : $signed(forvar771))) < $signed($unsigned($signed(reg775)))) >>> ($unsigned((^(~|(7'h40)))) ^ ({wire756} ?
          (^~reg778) : ($signed(reg769) ? {reg776} : reg774[(2'h3):(1'h1)])))))
        begin
          reg779 <= reg761;
          reg780 <= ($signed(wire755) ?
              {$unsigned($unsigned((reg765 - reg760)))} : $signed(reg776[(4'hc):(4'hb)]));
          reg781 <= $unsigned(reg777[(2'h3):(2'h3)]);
          for (forvar782 = (1'h0); (forvar782 < (3'h4)); forvar782 = (forvar782 + (1'h1)))
            begin
              reg783 <= $unsigned(reg751[(2'h3):(1'h0)]);
              reg784 <= $unsigned(reg762[(1'h0):(1'h0)]);
              reg785 = ($unsigned(reg779) >> reg773);
              reg786 <= $signed({{reg775[(4'hd):(4'h9)],
                      $signed((reg763 ? forvar782 : reg785))},
                  (forvar771 && wire754)});
            end
        end
      else
        begin
          for (forvar779 = (1'h0); (forvar779 < (2'h3)); forvar779 = (forvar779 + (1'h1)))
            begin
              reg780 <= (($unsigned((((8'hba) ?
                  (8'h9e) : reg765) ^~ (reg759 != (8'hb1)))) ^~ (reg773[(4'hc):(4'hb)] ?
                  $unsigned($unsigned(reg759)) : ($signed(wire747) ?
                      ((8'ha1) >>> reg758) : $signed(reg784)))) < $signed({$signed($signed(wire749)),
                  reg783}));
            end
          reg781 <= wire755[(4'h8):(3'h7)];
          reg782 = {(8'h9f),
              (reg761[(3'h7):(1'h0)] ? (8'h9d) : forvar771[(2'h3):(1'h0)])};
          reg783 <= {((~^$signed($signed(reg780))) >= ((reg751 ?
                      reg751[(1'h0):(1'h0)] : reg778) ?
                  reg779[(3'h7):(1'h0)] : ((reg786 ?
                      (8'hbd) : forvar772) >>> forvar779[(1'h0):(1'h0)])))};
          reg784 <= reg774[(2'h3):(1'h0)];
        end
      reg787 = (&((&($unsigned((8'hb8)) >>> reg757)) < $signed($signed($signed(reg778)))));
    end
  module788 modinst841 (wire840, clk, reg769, reg787, forvar782, reg764, reg770);
  always
    @(posedge clk) begin
      reg842 = (forvar779 >= ($unsigned(($unsigned(reg760) >= $signed((8'h9c)))) ?
          $unsigned((&$signed((8'h9e)))) : ($signed(((8'haf) ?
                  wire755 : forvar779)) ?
              (reg787 ?
                  $signed(reg769) : {reg786,
                      reg770}) : $signed($signed((8'hb1))))));
      reg843 <= (((^wire748) << (^~(^$unsigned(reg759)))) && (&(reg781[(2'h2):(2'h2)] ?
          (^~reg757[(3'h5):(2'h3)]) : ($signed(wire750) && $unsigned(reg786)))));
      for (forvar844 = (1'h0); (forvar844 < (1'h1)); forvar844 = (forvar844 + (1'h1)))
        begin
          reg845 <= (reg769 & reg751[(1'h0):(1'h0)]);
          reg846 = wire840[(1'h1):(1'h1)];
          reg847 <= ({($signed($unsigned(reg761)) ? (-(-(8'hbe))) : (8'h9c)),
                  reg763} ?
              reg775 : ($signed($signed({forvar772,
                  (8'ha2)})) || (~|forvar782[(1'h0):(1'h0)])));
          reg848 <= ({$unsigned((^wire750[(2'h2):(1'h1)]))} ?
              ({reg782[(1'h0):(1'h0)]} ?
                  reg757[(1'h1):(1'h0)] : reg776) : wire748);
          reg849 = $signed((($signed((~&reg780)) ?
              (8'hb2) : reg768[(1'h0):(1'h0)]) != forvar779[(1'h1):(1'h1)]));
        end
    end
  assign wire850 = $unsigned((reg775 ?
                       {reg781, $unsigned(wire756)} : (((reg782 ?
                                   reg765 : reg763) ?
                               $signed(reg775) : (^~reg787)) ?
                           ((8'hb4) != reg847) : (+$unsigned(reg778)))));
  always
    @(posedge clk) begin
      reg851 = (((^~reg845) <<< reg760) == reg757[(4'h8):(3'h4)]);
      for (forvar852 = (1'h0); (forvar852 < (1'h0)); forvar852 = (forvar852 + (1'h1)))
        begin
          reg853 <= (reg776[(2'h2):(1'h0)] + {reg758,
              (reg775 ? reg782[(1'h1):(1'h0)] : $unsigned($signed((8'hb9))))});
          reg854 <= (~^(7'h41));
          reg855 <= {(8'hbb)};
          reg856 <= {reg781};
          reg857 <= reg854;
        end
      reg858 <= ((($unsigned((-(7'h43))) ?
              $signed((reg773 ^ (8'hac))) : (8'h9c)) * reg857[(2'h3):(1'h1)]) ?
          (|((8'ha6) > (~^$unsigned((8'had))))) : (~(~|(~^wire756[(4'hb):(4'ha)]))));
      for (forvar859 = (1'h0); (forvar859 < (1'h1)); forvar859 = (forvar859 + (1'h1)))
        begin
          reg860 = $unsigned($signed(((&((8'hbd) ? reg773 : reg856)) ?
              $unsigned({reg752}) : {reg773})));
        end
    end
  always
    @(posedge clk) begin
      reg861 <= $signed(($signed(((wire748 ? reg760 : reg760) ?
          reg780 : $signed((8'ha8)))) ~^ reg787[(1'h0):(1'h0)]));
      reg862 <= reg785;
      reg863 <= {(+forvar779), wire850};
      reg864 <= ($signed(($signed(reg847[(5'h12):(1'h1)]) ?
          reg779[(1'h0):(1'h0)] : $unsigned(reg782))) && (+$signed(({(7'h44)} ?
          (reg787 || reg758) : reg860))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module613
#( parameter param718 = ((((+((8'hba) ^ (8'hb9))) + (((8'hab) ? (7'h44) : (7'h40)) & {(8'h9e), (8'ha3)})) ? (^~((~(8'ha0)) ? ((8'ha7) || (8'ha5)) : (~&(8'hae)))) : ((!(8'hae)) != (^~(~&(8'ha6))))) <<< ((|({(8'ha4), (8'hbe)} ? (~(7'h40)) : (8'haa))) >>> ((~|((8'ha3) > (8'ha6))) ? ((8'hbd) ? (+(8'hb2)) : ((8'ha6) ? (8'h9d) : (8'hb0))) : (!{(8'hbe)}))))
, parameter param719 = ((param718 ^~ (((param718 <= param718) ^~ (param718 ? (8'hbe) : param718)) | param718)) ^~ ((^(~((7'h44) ? param718 : param718))) ? (param718 ? (param718 | (~|param718)) : ((param718 ? param718 : (7'h44)) ? (^~param718) : (param718 * param718))) : param718)) )
(y, clk, wire614, wire615, wire616, wire617);
  output wire [(32'hed):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire614;
  input wire [(3'h4):(1'h0)] wire615;
  input wire signed [(3'h7):(1'h0)] wire616;
  input wire signed [(5'h12):(1'h0)] wire617;
  reg [(5'h15):(1'h0)] reg717 = (1'h0);
  reg [(3'h6):(1'h0)] reg716 = (1'h0);
  reg [(4'he):(1'h0)] reg715 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg714 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg713 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg712 = (1'h0);
  wire [(2'h2):(1'h0)] wire711;
  reg [(5'h15):(1'h0)] reg710 = (1'h0);
  wire [(5'h13):(1'h0)] wire709;
  reg [(4'he):(1'h0)] reg618 = (1'h0);
  reg [(2'h3):(1'h0)] reg619 = (1'h0);
  reg [(2'h3):(1'h0)] reg620 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire621;
  wire signed [(5'h13):(1'h0)] wire622;
  reg signed [(5'h13):(1'h0)] reg623 = (1'h0);
  reg [(2'h2):(1'h0)] reg624 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg625 = (1'h0);
  reg [(2'h2):(1'h0)] reg626 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg627 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg628 = (1'h0);
  wire [(2'h3):(1'h0)] wire707;
  assign y = {reg717,
                 reg716,
                 reg715,
                 reg714,
                 reg713,
                 reg712,
                 wire711,
                 reg710,
                 wire709,
                 reg618,
                 reg619,
                 reg620,
                 wire621,
                 wire622,
                 reg623,
                 reg624,
                 reg625,
                 reg626,
                 reg627,
                 reg628,
                 wire707,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg618 <= wire614[(4'ha):(3'h6)];
    end
  always
    @(posedge clk) begin
      reg619 <= ((wire615 ?
          reg618[(2'h2):(2'h2)] : ((((8'hb4) >> wire617) == (wire614 ?
              wire617 : wire616)) != $signed((8'hb4)))) <= (~&(~(-wire616[(3'h6):(1'h0)]))));
      reg620 <= {reg618};
    end
  assign wire621 = (^~($signed((reg620 ?
                       wire614 : $unsigned(wire615))) && reg618));
  assign wire622 = wire616[(3'h7):(3'h4)];
  always
    @(posedge clk) begin
      reg623 = (reg618[(3'h6):(1'h1)] >>> (wire621[(3'h7):(3'h5)] + $signed(wire621[(4'hb):(4'hb)])));
      reg624 = {(~&reg623),
          (~&$signed((reg623[(4'hf):(3'h4)] > ((8'hac) ? (8'hbb) : reg619))))};
      reg625 <= {wire621[(3'h4):(1'h0)],
          ($unsigned((~|$signed(wire616))) >> (!$unsigned(wire614[(4'h9):(3'h5)])))};
      reg626 = (~^wire617);
      reg627 <= $unsigned(wire614[(3'h7):(3'h5)]);
    end
  always
    @(posedge clk) begin
      reg628 <= wire617;
    end
  module629 modinst708 (.wire630(reg619), .wire632(reg628), .y(wire707), .wire634(wire617), .clk(clk), .wire631(reg623), .wire633(wire622));
  assign wire709 = reg619[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg710 <= reg624;
    end
  assign wire711 = (-wire616[(3'h6):(3'h5)]);
  always
    @(posedge clk) begin
      reg712 <= $unsigned(wire621[(3'h6):(3'h6)]);
      reg713 <= ((~|$signed($signed((^~reg624)))) ? (8'ha5) : wire621);
      reg714 <= $signed(((({wire621, reg618} >>> ((8'hae) * (8'haf))) ?
          $signed($unsigned(wire711)) : reg624[(2'h2):(1'h0)]) > {reg628,
          $signed($signed((8'h9c)))}));
      reg715 <= $signed(wire621);
      reg716 = (^~(^~$unsigned((+(reg714 <<< reg625)))));
    end
  always
    @(posedge clk) begin
      reg717 <= reg625;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module516
#( parameter param609 = (-((~|((8'hb2) != (~&(8'hba)))) >= (~(((8'haa) ? (8'h9d) : (8'ha6)) ? ((8'hb6) + (8'h9f)) : (7'h43)))))
, parameter param610 = param609 )
(y, clk, wire517, wire518, wire519, wire520, wire521);
  output wire [(32'h8d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire517;
  input wire [(4'hb):(1'h0)] wire518;
  input wire [(5'h12):(1'h0)] wire519;
  input wire [(5'h10):(1'h0)] wire520;
  input wire [(4'hb):(1'h0)] wire521;
  wire signed [(2'h3):(1'h0)] wire608;
  reg signed [(2'h3):(1'h0)] reg607 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar606 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg605 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg604 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar603 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg602 = (1'h0);
  reg [(4'h9):(1'h0)] forvar601 = (1'h0);
  wire [(3'h6):(1'h0)] wire522;
  wire [(2'h2):(1'h0)] wire523;
  wire [(5'h13):(1'h0)] wire524;
  wire [(4'hd):(1'h0)] wire525;
  wire signed [(3'h6):(1'h0)] wire526;
  wire [(4'he):(1'h0)] wire599;
  assign y = {wire608,
                 reg607,
                 forvar606,
                 reg605,
                 reg604,
                 forvar603,
                 reg602,
                 forvar601,
                 wire522,
                 wire523,
                 wire524,
                 wire525,
                 wire526,
                 wire599,
                 (1'h0)};
  assign wire522 = $signed({wire519[(3'h5):(1'h0)],
                       {wire519, (+$signed(wire519))}});
  assign wire523 = (~^($unsigned($signed(wire518[(2'h3):(2'h3)])) ?
                       ({{wire522},
                           (-wire521)} ~^ $signed({wire518})) : wire522[(3'h4):(1'h1)]));
  assign wire524 = {((8'hbe) ?
                           wire518[(3'h6):(2'h2)] : ($unsigned({wire517,
                                   wire520}) ?
                               ((wire520 ? wire522 : wire517) ?
                                   (!wire517) : $signed(wire518)) : {wire518,
                                   wire522}))};
  assign wire525 = (+({wire520[(4'hf):(4'he)]} ^~ ((wire523[(1'h0):(1'h0)] ?
                       $signed(wire520) : (!wire517)) | (~|wire517))));
  assign wire526 = wire520;
  module527 modinst600 (.wire528(wire520), .wire529(wire519), .clk(clk), .wire532(wire517), .wire530(wire524), .y(wire599), .wire531(wire518));
  always
    @(posedge clk) begin
      for (forvar601 = (1'h0); (forvar601 < (2'h2)); forvar601 = (forvar601 + (1'h1)))
        begin
          reg602 <= $unsigned(wire520);
          for (forvar603 = (1'h0); (forvar603 < (1'h0)); forvar603 = (forvar603 + (1'h1)))
            begin
              reg604 <= wire521;
              reg605 <= (((wire523[(2'h2):(2'h2)] ?
                  ($unsigned(forvar603) & $unsigned(wire522)) : $signed($unsigned(forvar601))) - ($signed(wire525) ?
                  wire519 : ((+wire526) < (&wire526)))) | $unsigned(wire520));
            end
        end
      for (forvar606 = (1'h0); (forvar606 < (1'h1)); forvar606 = (forvar606 + (1'h1)))
        begin
          reg607 <= ((forvar606[(1'h1):(1'h0)] >>> (wire523[(2'h2):(1'h1)] ?
              {(wire525 * forvar601)} : wire522)) ^~ (wire517[(1'h0):(1'h0)] ?
              {$unsigned((~&wire524))} : ({{wire525}, wire523[(1'h1):(1'h0)]} ?
                  ((~|wire523) ?
                      wire517 : $unsigned(forvar603)) : {(wire519 && wire525)})));
        end
    end
  assign wire608 = ((($unsigned((reg605 ? forvar601 : (8'ha3))) ?
                           $unsigned(wire523) : (~&wire520)) ?
                       wire517 : reg602) <<< $signed($unsigned((-((8'hb1) ?
                       wire523 : forvar601)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module202
#( parameter param497 = ((8'hbd) ^~ (({((7'h44) <<< (8'hb0)), ((8'ha7) << (8'h9e))} ? ({(8'haf)} >> (^(8'hae))) : {(8'ha9), ((7'h43) ? (8'hb3) : (8'ha5))}) ? (-(((8'haf) ? (8'ha1) : (8'hb6)) ? (!(8'hbb)) : ((8'h9f) * (7'h44)))) : ((8'hbd) ? (((8'hbf) ? (8'hb6) : (8'hb5)) ? ((8'haf) ? (8'hbd) : (8'ha8)) : ((8'ha6) ? (8'ha6) : (8'ha5))) : (((8'hb9) ? (8'haf) : (8'hb2)) * (^(8'ha9))))))
, parameter param498 = {param497} )
(y, clk, wire203, wire204, wire205, wire206);
  output wire [(32'h248):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire203;
  input wire [(4'hc):(1'h0)] wire204;
  input wire [(5'h13):(1'h0)] wire205;
  input wire [(5'h15):(1'h0)] wire206;
  wire signed [(4'hb):(1'h0)] wire496;
  wire [(4'he):(1'h0)] wire495;
  wire [(5'h10):(1'h0)] wire494;
  wire [(4'h8):(1'h0)] wire493;
  reg [(4'hc):(1'h0)] reg492 = (1'h0);
  reg [(3'h4):(1'h0)] reg491 = (1'h0);
  wire [(3'h6):(1'h0)] wire490;
  wire [(2'h3):(1'h0)] wire489;
  wire signed [(2'h3):(1'h0)] wire488;
  reg signed [(4'hf):(1'h0)] forvar207 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg208 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar209 = (1'h0);
  reg [(4'hb):(1'h0)] reg210 = (1'h0);
  reg [(4'h8):(1'h0)] reg211 = (1'h0);
  reg [(5'h10):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg213 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg214 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg215 = (1'h0);
  wire [(4'h8):(1'h0)] wire216;
  reg signed [(5'h10):(1'h0)] reg217 = (1'h0);
  reg [(4'he):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg219 = (1'h0);
  reg [(4'he):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar221 = (1'h0);
  reg [(4'h9):(1'h0)] reg222 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg223 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar224 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg225 = (1'h0);
  reg [(2'h2):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg228 = (1'h0);
  reg [(4'he):(1'h0)] reg229 = (1'h0);
  reg [(5'h15):(1'h0)] forvar230 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg231 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire232;
  wire [(5'h12):(1'h0)] wire337;
  wire [(5'h15):(1'h0)] wire339;
  reg [(4'ha):(1'h0)] reg340 = (1'h0);
  reg [(4'he):(1'h0)] reg341 = (1'h0);
  reg [(4'hc):(1'h0)] reg342 = (1'h0);
  reg [(4'hc):(1'h0)] reg343 = (1'h0);
  reg [(5'h13):(1'h0)] reg344 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg345 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg346 = (1'h0);
  wire [(5'h10):(1'h0)] wire399;
  wire signed [(5'h13):(1'h0)] wire486;
  assign y = {wire496,
                 wire495,
                 wire494,
                 wire493,
                 reg492,
                 reg491,
                 wire490,
                 wire489,
                 wire488,
                 forvar207,
                 reg208,
                 forvar209,
                 reg210,
                 reg211,
                 reg212,
                 reg213,
                 reg214,
                 reg215,
                 wire216,
                 reg217,
                 reg218,
                 reg219,
                 reg220,
                 forvar221,
                 reg222,
                 reg223,
                 forvar224,
                 reg225,
                 reg226,
                 reg227,
                 reg228,
                 reg229,
                 forvar230,
                 reg231,
                 wire232,
                 wire337,
                 wire339,
                 reg340,
                 reg341,
                 reg342,
                 reg343,
                 reg344,
                 reg345,
                 reg346,
                 wire399,
                 wire486,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar207 = (1'h0); (forvar207 < (2'h2)); forvar207 = (forvar207 + (1'h1)))
        begin
          reg208 = wire206;
          for (forvar209 = (1'h0); (forvar209 < (1'h1)); forvar209 = (forvar209 + (1'h1)))
            begin
              reg210 <= (~^($signed(wire203) ^~ $unsigned((^~reg208))));
              reg211 <= forvar209;
              reg212 <= (~&$signed($signed((!$unsigned(wire203)))));
              reg213 <= $unsigned($unsigned($signed(($unsigned(reg210) ?
                  (~&wire203) : $unsigned(reg208)))));
            end
        end
      reg214 <= $signed($signed($signed((^(~&forvar209)))));
      reg215 <= $signed(((|$unsigned(reg208)) ?
          ($signed({(8'ha1), wire204}) != (!(reg210 ?
              (8'hb7) : reg210))) : (wire205 ?
              wire205 : ((forvar207 ? reg212 : forvar207) ^ {(8'hbc),
                  wire203}))));
    end
  assign wire216 = wire206;
  always
    @(posedge clk) begin
      reg217 <= $signed((((~(reg211 == wire205)) ?
              wire216 : wire203[(4'hd):(3'h4)]) ?
          (+$signed((forvar207 && wire203))) : $unsigned(({reg212} ?
              $unsigned((8'h9f)) : (forvar207 ? wire206 : forvar207)))));
      reg218 <= (~&((|{wire216[(3'h5):(3'h4)], wire216}) ?
          $unsigned(wire206) : wire216));
      reg219 <= (!(~$signed((~(-reg208)))));
    end
  always
    @(posedge clk) begin
      reg220 <= {wire205[(3'h7):(3'h5)],
          ({reg208[(4'h8):(2'h2)],
              $unsigned(((7'h43) ? reg212 : reg210))} > wire204)};
      for (forvar221 = (1'h0); (forvar221 < (2'h3)); forvar221 = (forvar221 + (1'h1)))
        begin
          reg222 <= wire216[(1'h1):(1'h0)];
          reg223 <= (7'h41);
        end
      for (forvar224 = (1'h0); (forvar224 < (2'h3)); forvar224 = (forvar224 + (1'h1)))
        begin
          reg225 = (((^$signed(reg219[(4'hb):(4'ha)])) ?
              $signed(({reg217} ?
                  wire206[(2'h3):(1'h0)] : $unsigned(reg217))) : (-(!(forvar224 ?
                  reg219 : reg215)))) >> {({$signed(reg219),
                  (reg208 ? wire205 : reg210)} ~^ $unsigned($signed(wire204))),
              ($unsigned($unsigned(forvar207)) < (8'had))});
          reg226 <= $unsigned(forvar207[(4'ha):(3'h4)]);
          reg227 <= {($signed(reg208) << reg222),
              ((wire206 ?
                  $unsigned((reg214 ?
                      forvar207 : wire203)) : (+wire216[(1'h0):(1'h0)])) <= reg222[(3'h7):(3'h4)])};
          reg228 = $unsigned(reg222);
        end
      reg229 <= reg226[(1'h0):(1'h0)];
      for (forvar230 = (1'h0); (forvar230 < (1'h0)); forvar230 = (forvar230 + (1'h1)))
        begin
          reg231 = (^~$unsigned(reg213));
        end
    end
  assign wire232 = reg231[(3'h7):(3'h7)];
  module233 modinst338 (wire337, clk, reg229, reg212, wire204, reg215);
  assign wire339 = reg211[(3'h6):(3'h4)];
  always
    @(posedge clk) begin
      reg340 <= reg223;
      reg341 <= (^$unsigned(reg227[(4'h8):(3'h7)]));
    end
  always
    @(posedge clk) begin
      reg342 <= reg218[(4'hd):(4'h9)];
      reg343 = (($unsigned($unsigned((wire204 ? (8'hb5) : (7'h42)))) ?
              reg340[(2'h3):(2'h2)] : (({(7'h44)} * $signed(reg215)) ^ forvar221)) ?
          ({$unsigned((reg212 - (8'hb5))),
              {((8'ha2) <<< (8'hbe)), (-(8'hbd))}} >= ({(wire337 <= reg222),
              wire339[(4'ha):(2'h3)]} <= (wire232[(2'h2):(2'h2)] ?
              (wire206 | wire337) : (wire232 ~^ reg218)))) : forvar221[(4'hd):(3'h4)]);
      reg344 = $signed(((reg227 || $signed($unsigned(forvar224))) ?
          $signed($signed(reg211[(2'h3):(2'h2)])) : wire339));
      reg345 <= ($signed(($signed((^~reg222)) ?
          $signed($signed(reg220)) : (8'hb8))) ^~ $signed($unsigned((reg226 ?
          (^reg228) : reg223[(3'h6):(3'h5)]))));
      reg346 <= $unsigned(({reg212[(3'h4):(2'h3)], wire216} ?
          (reg345[(3'h6):(1'h0)] ?
              forvar209 : reg208) : (^$unsigned((reg222 < forvar221)))));
    end
  module347 modinst400 (.clk(clk), .wire351(reg214), .wire350(wire205), .wire349(reg212), .y(wire399), .wire348(reg227));
  module401 modinst487 (.wire404(reg208), .wire406(wire204), .clk(clk), .wire403(reg211), .y(wire486), .wire405(reg341), .wire402(reg210));
  assign wire488 = wire203;
  assign wire489 = ((reg218 ?
                       $signed((|(reg344 != wire203))) : {(((8'h9d) ?
                                   reg344 : reg217) ?
                               (forvar221 * wire206) : (+reg217))}) ~^ ($unsigned(((8'ha2) > $unsigned((8'hb6)))) ?
                       ({$unsigned(wire339), reg231} ?
                           $unsigned({reg223}) : reg226) : {((reg345 > wire337) ?
                               ((8'hac) | wire399) : (reg343 ?
                                   wire399 : reg220)),
                           {$signed(wire216), (reg220 <= wire486)}}));
  assign wire490 = $signed(forvar230);
  always
    @(posedge clk) begin
      reg491 <= (forvar221 << reg229);
      reg492 <= forvar207;
    end
  assign wire493 = ((reg223 ? reg222[(1'h1):(1'h0)] : reg227) * reg226);
  assign wire494 = (7'h44);
  assign wire495 = (8'hb1);
  assign wire496 = reg344;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module401
#( parameter param484 = ({((((8'had) * (8'hbb)) ? (+(7'h41)) : ((8'h9e) ? (8'haf) : (8'h9c))) ? {((8'hae) ? (8'ha3) : (8'hba)), (^~(8'hbb))} : ((8'hbb) ^~ ((8'haf) <= (8'hbb)))), {{((8'hae) + (8'hab))}}} ? (((8'hb2) ~^ (((8'hac) ? (8'ha6) : (8'ha7)) ? ((8'h9d) ? (8'hae) : (8'hb5)) : ((8'had) ? (8'h9e) : (8'hbe)))) * {(((8'h9c) && (8'hb3)) >> ((8'ha4) > (8'hbd)))}) : {(^((~|(8'hac)) >= {(7'h40)})), ((((8'ha3) >= (8'ha5)) ? ((8'ha4) != (8'hbf)) : ((8'had) < (8'hb2))) >= (((8'ha3) ? (8'h9d) : (8'ha3)) && ((8'ha5) | (8'ha8))))})
, parameter param485 = param484 )
(y, clk, wire406, wire405, wire404, wire403, wire402);
  output wire [(32'h395):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire406;
  input wire [(4'he):(1'h0)] wire405;
  input wire [(5'h11):(1'h0)] wire404;
  input wire [(3'h5):(1'h0)] wire403;
  input wire [(4'hb):(1'h0)] wire402;
  wire signed [(4'h9):(1'h0)] wire483;
  reg [(4'hd):(1'h0)] reg482 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg481 = (1'h0);
  reg [(3'h6):(1'h0)] forvar480 = (1'h0);
  reg [(5'h12):(1'h0)] reg479 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg478 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg477 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg476 = (1'h0);
  reg [(4'ha):(1'h0)] reg475 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg474 = (1'h0);
  reg signed [(4'he):(1'h0)] reg473 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg472 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg471 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar470 = (1'h0);
  reg [(3'h4):(1'h0)] reg469 = (1'h0);
  reg [(3'h4):(1'h0)] reg468 = (1'h0);
  reg [(5'h10):(1'h0)] reg467 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg466 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg465 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg464 = (1'h0);
  reg [(2'h3):(1'h0)] reg463 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar462 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg461 = (1'h0);
  reg signed [(4'he):(1'h0)] reg460 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg459 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg458 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg457 = (1'h0);
  wire [(3'h6):(1'h0)] wire456;
  reg signed [(5'h13):(1'h0)] reg455 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg452 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg451 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg450 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg449 = (1'h0);
  reg [(5'h13):(1'h0)] reg448 = (1'h0);
  reg [(5'h14):(1'h0)] reg447 = (1'h0);
  reg [(5'h13):(1'h0)] forvar446 = (1'h0);
  reg [(5'h14):(1'h0)] reg445 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg444 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar443 = (1'h0);
  reg [(2'h3):(1'h0)] reg442 = (1'h0);
  reg [(5'h13):(1'h0)] reg441 = (1'h0);
  reg [(4'hc):(1'h0)] reg440 = (1'h0);
  reg [(3'h6):(1'h0)] forvar439 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg438 = (1'h0);
  reg [(5'h10):(1'h0)] forvar437 = (1'h0);
  reg [(3'h7):(1'h0)] reg436 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg435 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg434 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg433 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg432 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg431 = (1'h0);
  reg [(5'h11):(1'h0)] forvar430 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg429 = (1'h0);
  reg [(4'hb):(1'h0)] reg428 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire427;
  wire signed [(4'hf):(1'h0)] wire426;
  wire signed [(3'h6):(1'h0)] wire425;
  wire [(2'h3):(1'h0)] wire424;
  reg [(4'hd):(1'h0)] reg423 = (1'h0);
  reg [(2'h3):(1'h0)] reg422 = (1'h0);
  reg [(4'hd):(1'h0)] reg421 = (1'h0);
  wire signed [(4'he):(1'h0)] wire420;
  reg signed [(3'h6):(1'h0)] reg419 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar418 = (1'h0);
  reg [(4'he):(1'h0)] reg417 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg416 = (1'h0);
  reg [(3'h4):(1'h0)] reg415 = (1'h0);
  reg [(5'h15):(1'h0)] reg414 = (1'h0);
  reg [(5'h10):(1'h0)] forvar413 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg412 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg411 = (1'h0);
  reg [(4'he):(1'h0)] forvar410 = (1'h0);
  reg [(4'hc):(1'h0)] reg409 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg408 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg407 = (1'h0);
  assign y = {wire483,
                 reg482,
                 reg481,
                 forvar480,
                 reg479,
                 reg478,
                 reg477,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 forvar470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 forvar462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 wire456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 reg447,
                 forvar446,
                 reg445,
                 reg444,
                 forvar443,
                 reg442,
                 reg441,
                 reg440,
                 forvar439,
                 reg438,
                 forvar437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 forvar430,
                 reg429,
                 reg428,
                 wire427,
                 wire426,
                 wire425,
                 wire424,
                 reg423,
                 reg422,
                 reg421,
                 wire420,
                 reg419,
                 forvar418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 forvar413,
                 reg412,
                 reg411,
                 forvar410,
                 reg409,
                 reg408,
                 reg407,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg407 = $unsigned($signed((~{$unsigned((8'hac))})));
      reg408 <= $unsigned(reg407[(1'h0):(1'h0)]);
      reg409 = ((reg407 ?
              (wire406[(1'h0):(1'h0)] | (~&$signed(wire406))) : ($signed((wire402 ^~ (8'haf))) <<< $signed($signed(wire405)))) ?
          (reg407 <<< $signed($signed(wire402))) : wire406);
    end
  always
    @(posedge clk) begin
      for (forvar410 = (1'h0); (forvar410 < (1'h0)); forvar410 = (forvar410 + (1'h1)))
        begin
          reg411 = (wire405 | {wire402});
        end
      reg412 = wire404[(4'h9):(1'h1)];
      for (forvar413 = (1'h0); (forvar413 < (2'h3)); forvar413 = (forvar413 + (1'h1)))
        begin
          reg414 = $unsigned((~|$unsigned({forvar413[(4'h9):(3'h7)],
              $unsigned(reg407)})));
          reg415 <= (+(~|$unsigned((!$unsigned((8'ha9))))));
        end
    end
  always
    @(posedge clk) begin
      reg416 <= $unsigned(wire404[(3'h7):(1'h0)]);
      reg417 <= (8'hac);
      for (forvar418 = (1'h0); (forvar418 < (1'h0)); forvar418 = (forvar418 + (1'h1)))
        begin
          reg419 <= reg407[(3'h5):(3'h4)];
        end
    end
  assign wire420 = (($unsigned($signed($unsigned(reg416))) * (|wire406)) ?
                       reg409[(1'h1):(1'h1)] : reg419);
  always
    @(posedge clk) begin
      reg421 <= $signed({reg414[(4'h9):(1'h0)],
          $unsigned($unsigned((|wire406)))});
      reg422 = {{$unsigned(reg409)}};
      reg423 <= (|wire406);
    end
  assign wire424 = $unsigned($unsigned((wire403 ~^ reg415)));
  assign wire425 = (^(($unsigned($unsigned((8'hb7))) <<< (8'hb5)) >= $signed((wire403 ^~ (reg423 ?
                       wire406 : wire405)))));
  assign wire426 = {(&$unsigned(((wire405 & (8'hac)) ?
                           (reg416 < reg414) : {reg412, (8'hb5)})))};
  assign wire427 = (~|(forvar418 && $unsigned(reg412)));
  always
    @(posedge clk) begin
      reg428 <= reg408;
      reg429 <= $signed((|wire404[(3'h5):(2'h2)]));
    end
  always
    @(posedge clk) begin
      for (forvar430 = (1'h0); (forvar430 < (2'h3)); forvar430 = (forvar430 + (1'h1)))
        begin
          reg431 <= ((^((8'h9d) <= ((^~reg428) ?
                  $signed((8'hbe)) : forvar430[(1'h0):(1'h0)]))) ?
              (forvar418 ?
                  $signed((~$unsigned(forvar430))) : (^wire426)) : (wire403[(3'h4):(1'h0)] >= reg422));
          reg432 <= (8'hbf);
          reg433 <= ({(forvar418[(4'h8):(3'h4)] + {reg419}),
              (|($unsigned(wire425) ?
                  reg409[(4'hc):(4'h9)] : reg412[(5'h10):(3'h5)]))} * $signed((+$unsigned(reg414))));
          reg434 <= (8'hba);
        end
      reg435 <= ((((~wire406) ? (^reg432[(1'h1):(1'h0)]) : (8'h9e)) ?
          {(&$unsigned((8'hbb)))} : reg407) > wire426);
      reg436 <= (reg416 | {$unsigned(wire425[(2'h3):(1'h1)])});
    end
  always
    @(posedge clk) begin
      for (forvar437 = (1'h0); (forvar437 < (1'h0)); forvar437 = (forvar437 + (1'h1)))
        begin
          reg438 = (+reg409[(2'h2):(1'h1)]);
          for (forvar439 = (1'h0); (forvar439 < (1'h1)); forvar439 = (forvar439 + (1'h1)))
            begin
              reg440 <= (|reg408);
            end
          reg441 <= ({$signed(reg435)} - reg436);
        end
      reg442 <= ($signed($unsigned({wire425})) ?
          wire425[(1'h1):(1'h1)] : (-$signed(((^reg422) ^ (reg440 ?
              wire425 : forvar437)))));
      for (forvar443 = (1'h0); (forvar443 < (2'h2)); forvar443 = (forvar443 + (1'h1)))
        begin
          reg444 = reg411;
          reg445 <= (~&$unsigned($signed(reg442[(2'h3):(1'h1)])));
          for (forvar446 = (1'h0); (forvar446 < (1'h1)); forvar446 = (forvar446 + (1'h1)))
            begin
              reg447 = (forvar446 ?
                  (^~$unsigned(((reg429 >> reg442) != (8'hb4)))) : (|($signed(reg416[(2'h3):(2'h2)]) == $signed($signed((8'had))))));
              reg448 = $signed($signed(wire427[(4'he):(4'hb)]));
              reg449 <= $unsigned(reg447);
            end
          reg450 <= (8'ha0);
          reg451 <= ($signed(((^~(reg417 - reg445)) ?
                  ($signed(reg429) ?
                      $unsigned(reg412) : reg442[(2'h3):(1'h1)]) : $signed({reg433}))) ?
              $signed((8'ha3)) : ($unsigned(((~&forvar430) == wire403)) ?
                  ($signed((forvar446 || wire425)) ^ wire405) : {(((8'hb1) * reg447) - reg435)}));
        end
      reg452 <= {forvar446};
      reg453 = forvar418[(2'h2):(1'h1)];
    end
  always
    @(posedge clk) begin
      reg454 = (forvar437 <= forvar443);
      reg455 <= $unsigned((reg441 + ({{(7'h44)}} ?
          (+((8'hb4) ? reg435 : reg436)) : ((forvar413 ? forvar443 : reg417) ?
              reg451[(1'h1):(1'h0)] : (wire424 * wire420)))));
    end
  assign wire456 = $unsigned((~&(-(~^(|(8'ha9))))));
  always
    @(posedge clk) begin
      reg457 <= $unsigned($unsigned(reg441[(2'h3):(2'h3)]));
      reg458 <= ($unsigned((+(((8'hb3) ? reg411 : reg421) ?
          (reg452 ?
              (8'hb1) : reg433) : (&forvar443)))) ^ (({{reg438}} <<< (reg407 & $signed(wire426))) ?
          (((forvar418 ? forvar437 : reg435) ^~ (|wire456)) ?
              $signed($unsigned(reg450)) : (^reg433)) : $unsigned(wire425)));
    end
  always
    @(posedge clk) begin
      reg459 <= (((reg415[(3'h4):(3'h4)] ?
              {$signed(forvar413), $unsigned(reg449)} : reg432) ?
          (({reg448} < (forvar418 < reg429)) ?
              reg428[(2'h2):(1'h1)] : $signed(reg458[(4'h9):(1'h0)])) : (reg415[(3'h4):(1'h1)] ?
              {wire427, $signed(wire404)} : forvar413)) || reg417);
      reg460 <= $unsigned((~&forvar437));
      reg461 = ((8'hb7) ? $unsigned(reg451) : $unsigned(forvar446));
    end
  always
    @(posedge clk) begin
      for (forvar462 = (1'h0); (forvar462 < (1'h1)); forvar462 = (forvar462 + (1'h1)))
        begin
          reg463 <= $signed((!$unsigned((^$signed(reg448)))));
          reg464 = (~|reg445);
          reg465 <= reg411;
        end
      reg466 <= reg423[(2'h3):(2'h2)];
      reg467 <= $signed($unsigned(((^$unsigned(reg434)) ?
          (^~reg421) : $unsigned(forvar430))));
      if ($unsigned((~{$signed((^(8'ha6))), reg459[(1'h0):(1'h0)]})))
        begin
          reg468 <= (forvar413[(1'h0):(1'h0)] | $unsigned($unsigned(reg464[(3'h7):(3'h5)])));
          reg469 <= $signed($signed((-(+(reg451 * reg466)))));
          for (forvar470 = (1'h0); (forvar470 < (1'h1)); forvar470 = (forvar470 + (1'h1)))
            begin
              reg471 <= (~^wire456[(2'h3):(2'h2)]);
              reg472 <= (reg454 <= $signed((({(8'h9c),
                  reg419} <<< reg468[(1'h0):(1'h0)]) << reg415)));
              reg473 = $unsigned((+($signed((^~reg409)) ?
                  (&(~^(8'h9f))) : $unsigned((!reg461)))));
            end
          reg474 = (&({($signed(reg458) & {reg450})} ?
              ((~^$signed(forvar418)) ?
                  $unsigned($unsigned(reg442)) : $unsigned((|reg448))) : reg467));
        end
      else
        begin
          reg468 <= $unsigned((forvar437[(4'h9):(4'h9)] ?
              $unsigned(({reg416, wire420} ?
                  $signed(reg412) : (reg468 || wire405))) : (|($unsigned(reg440) == (forvar470 ?
                  reg464 : reg451)))));
          reg469 <= (8'ha4);
          for (forvar470 = (1'h0); (forvar470 < (3'h4)); forvar470 = (forvar470 + (1'h1)))
            begin
              reg471 = (wire403[(3'h4):(1'h1)] && reg469);
            end
          reg472 <= $signed((8'hb9));
        end
      reg475 = ({$unsigned($unsigned(reg411[(4'he):(3'h6)]))} ?
          (~($unsigned({reg450}) > reg471[(4'hf):(4'h9)])) : ($signed($signed(((8'haf) ?
              reg474 : reg440))) != forvar443[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg476 <= $unsigned((reg433 ?
          $unsigned($signed((reg459 ?
              wire425 : wire420))) : $signed($unsigned((reg423 == reg457)))));
      reg477 <= $unsigned({(^~(&$unsigned(reg476))),
          $signed(reg432[(1'h0):(1'h0)])});
      reg478 <= ((~|(|reg432[(1'h1):(1'h1)])) <<< (($unsigned((forvar446 ?
              (8'hb9) : reg411)) ?
          ((reg436 ? reg467 : reg433) ?
              $signed(reg411) : (-reg416)) : (reg449 >> (reg415 << (8'hb3)))) + (reg468[(2'h3):(2'h2)] ?
          ((reg463 ? reg474 : reg458) ^ $signed(reg474)) : wire403)));
      reg479 = reg460;
    end
  always
    @(posedge clk) begin
      for (forvar480 = (1'h0); (forvar480 < (1'h0)); forvar480 = (forvar480 + (1'h1)))
        begin
          reg481 <= {(^({(reg412 ? reg450 : forvar430), (forvar446 != reg433)} ?
                  (reg475[(1'h0):(1'h0)] ?
                      (reg469 ?
                          reg469 : forvar462) : (reg407 >>> forvar413)) : wire405[(4'hc):(3'h6)]))};
          reg482 <= {reg475,
              $unsigned(((^~(^~reg457)) * wire425[(3'h6):(1'h0)]))};
        end
    end
  assign wire483 = reg442[(1'h0):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module347
#(parameter param398 = (!(8'hba)))
(y, clk, wire351, wire350, wire349, wire348);
  output wire [(32'h222):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire351;
  input wire signed [(4'he):(1'h0)] wire350;
  input wire [(4'he):(1'h0)] wire349;
  input wire [(5'h15):(1'h0)] wire348;
  wire [(5'h15):(1'h0)] wire397;
  reg signed [(4'he):(1'h0)] reg396 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg395 = (1'h0);
  reg [(3'h6):(1'h0)] reg394 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg393 = (1'h0);
  reg [(5'h13):(1'h0)] forvar392 = (1'h0);
  reg [(2'h2):(1'h0)] reg391 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg390 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire389;
  reg signed [(3'h5):(1'h0)] reg388 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg387 = (1'h0);
  wire [(4'he):(1'h0)] wire386;
  wire [(5'h11):(1'h0)] wire385;
  reg signed [(4'hd):(1'h0)] reg384 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg383 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg382 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg381 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar380 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar379 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg378 = (1'h0);
  wire [(4'hd):(1'h0)] wire377;
  reg signed [(4'hc):(1'h0)] reg376 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg375 = (1'h0);
  reg [(2'h2):(1'h0)] reg374 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg373 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg372 = (1'h0);
  reg [(4'he):(1'h0)] reg371 = (1'h0);
  reg [(5'h15):(1'h0)] reg370 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg369 = (1'h0);
  reg signed [(4'he):(1'h0)] reg368 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar367 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar366 = (1'h0);
  reg [(4'hd):(1'h0)] reg365 = (1'h0);
  reg [(4'hb):(1'h0)] reg364 = (1'h0);
  reg [(2'h2):(1'h0)] reg363 = (1'h0);
  reg [(5'h11):(1'h0)] reg362 = (1'h0);
  reg [(5'h12):(1'h0)] forvar361 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg360 = (1'h0);
  reg [(3'h5):(1'h0)] reg359 = (1'h0);
  reg [(4'hf):(1'h0)] reg358 = (1'h0);
  reg [(4'hb):(1'h0)] reg357 = (1'h0);
  reg [(3'h4):(1'h0)] forvar356 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar355 = (1'h0);
  reg signed [(4'he):(1'h0)] reg354 = (1'h0);
  reg signed [(4'he):(1'h0)] reg353 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar352 = (1'h0);
  assign y = {wire397,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 forvar392,
                 reg391,
                 reg390,
                 wire389,
                 reg388,
                 reg387,
                 wire386,
                 wire385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 forvar380,
                 forvar379,
                 reg378,
                 wire377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 forvar367,
                 forvar366,
                 reg365,
                 reg364,
                 reg363,
                 reg362,
                 forvar361,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 forvar356,
                 forvar355,
                 reg354,
                 reg353,
                 forvar352,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar352 = (1'h0); (forvar352 < (1'h1)); forvar352 = (forvar352 + (1'h1)))
        begin
          reg353 <= wire351;
          reg354 = (!(8'ha6));
        end
      for (forvar355 = (1'h0); (forvar355 < (3'h4)); forvar355 = (forvar355 + (1'h1)))
        begin
          for (forvar356 = (1'h0); (forvar356 < (2'h3)); forvar356 = (forvar356 + (1'h1)))
            begin
              reg357 <= ((forvar355 ?
                      ($unsigned($unsigned(wire348)) ?
                          $signed(forvar352) : $signed(reg353)) : (^$signed({wire348,
                          forvar356}))) ?
                  (reg353 ?
                      forvar352 : wire351[(3'h5):(2'h2)]) : $unsigned({(~|(~^reg354))}));
            end
          reg358 <= {$signed($signed((^$unsigned(wire349))))};
          reg359 <= {reg354[(3'h4):(3'h4)],
              $unsigned({$unsigned($unsigned(wire348)),
                  $signed(((7'h40) ^ wire349))})};
          reg360 <= reg358;
          for (forvar361 = (1'h0); (forvar361 < (1'h0)); forvar361 = (forvar361 + (1'h1)))
            begin
              reg362 <= (wire351 ^ ((-{reg360}) - (~wire348)));
              reg363 = wire351;
              reg364 <= wire348;
              reg365 <= {((^~((8'ha6) ?
                          (reg363 ? reg363 : (7'h44)) : (~|reg360))) ?
                      $signed($unsigned(wire348[(5'h13):(2'h3)])) : $unsigned(((forvar355 << reg358) < ((8'hbb) ?
                          forvar361 : forvar352))))};
            end
        end
      for (forvar366 = (1'h0); (forvar366 < (1'h1)); forvar366 = (forvar366 + (1'h1)))
        begin
          for (forvar367 = (1'h0); (forvar367 < (2'h3)); forvar367 = (forvar367 + (1'h1)))
            begin
              reg368 = ((^$unsigned(reg358[(3'h4):(2'h2)])) ^~ forvar361[(4'hf):(3'h7)]);
              reg369 = $unsigned((^reg358[(2'h3):(1'h1)]));
              reg370 <= $signed($signed($signed($unsigned((^forvar367)))));
              reg371 = $unsigned(forvar355);
              reg372 = (|{wire351[(2'h3):(2'h2)], reg363});
            end
          reg373 <= (~&$unsigned({((reg368 ? reg354 : forvar356) ?
                  reg365 : {reg368})}));
          reg374 <= $unsigned(((^forvar355) ?
              {($unsigned(reg358) ?
                      (+wire350) : (~|reg358))} : $unsigned((-(wire350 >> forvar355)))));
          reg375 <= $signed($signed({{{reg370, (8'hba)}},
              $signed($signed((8'hbf)))}));
        end
      reg376 = ($signed(reg358[(4'hd):(3'h4)]) ?
          ({(8'had)} ^ $signed(reg371[(3'h7):(2'h3)])) : reg364);
    end
  assign wire377 = reg376[(4'hc):(1'h0)];
  always
    @(posedge clk) begin
      reg378 <= $unsigned(({(+(~&forvar356))} > $unsigned($unsigned($unsigned(reg364)))));
      for (forvar379 = (1'h0); (forvar379 < (1'h1)); forvar379 = (forvar379 + (1'h1)))
        begin
          for (forvar380 = (1'h0); (forvar380 < (3'h4)); forvar380 = (forvar380 + (1'h1)))
            begin
              reg381 <= reg359[(2'h2):(1'h0)];
              reg382 <= (($signed(($unsigned(forvar355) == $signed(reg364))) + $unsigned(forvar355[(4'h8):(1'h1)])) ^ (~^reg354));
            end
          reg383 <= (&({forvar367[(4'ha):(3'h5)]} ?
              $signed($signed((reg372 * reg363))) : ($unsigned((reg369 ?
                  reg369 : reg368)) >>> {wire351[(2'h3):(2'h3)],
                  $signed(wire349)})));
          reg384 = $unsigned(((+(~reg365[(2'h3):(1'h1)])) * forvar380));
        end
    end
  assign wire385 = reg364;
  assign wire386 = reg363[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg387 <= (!(^$signed((~(reg378 * (8'had))))));
      reg388 <= reg363;
    end
  assign wire389 = wire349;
  always
    @(posedge clk) begin
      reg390 = ((wire348 ?
          (wire389[(1'h1):(1'h1)] >>> $signed((&reg353))) : (|$signed(reg359[(1'h1):(1'h0)]))) >>> ((^$signed($unsigned(forvar355))) ^~ $unsigned((^(reg382 ?
          wire350 : forvar355)))));
      reg391 = wire350;
      for (forvar392 = (1'h0); (forvar392 < (2'h3)); forvar392 = (forvar392 + (1'h1)))
        begin
          reg393 <= ($unsigned((~(forvar361[(3'h4):(2'h2)] ?
                  reg363 : reg381))) ?
              $unsigned($unsigned(($signed(reg354) >= (-wire386)))) : wire351[(2'h3):(2'h3)]);
        end
      reg394 <= $unsigned(forvar356[(2'h3):(1'h1)]);
      reg395 <= {$unsigned(reg391)};
    end
  always
    @(posedge clk) begin
      reg396 <= (reg393[(1'h0):(1'h0)] ?
          forvar392 : $signed(($unsigned($unsigned(forvar379)) ?
              $unsigned(((8'hae) ?
                  (8'hb2) : (7'h40))) : ((reg360 ^ reg353) != $signed((8'h9e))))));
    end
  assign wire397 = (reg396 ?
                       reg363 : $signed($unsigned(($unsigned(reg360) ?
                           (reg393 > reg383) : (~&reg387)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module233
#( parameter param336 = {{({(-(8'hbd)), ((8'hb3) ? (7'h42) : (8'hb3))} ? ({(8'hba)} ? (-(8'ha8)) : ((8'hb5) ^ (8'ha3))) : (((8'hb4) ^~ (8'hbf)) * ((8'ha3) == (8'hae))))}} )
(y, clk, wire237, wire236, wire235, wire234);
  output wire [(32'h473):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire237;
  input wire signed [(5'h10):(1'h0)] wire236;
  input wire [(4'hc):(1'h0)] wire235;
  input wire [(3'h4):(1'h0)] wire234;
  reg [(4'ha):(1'h0)] reg335 = (1'h0);
  wire [(5'h12):(1'h0)] wire334;
  wire [(4'ha):(1'h0)] wire333;
  wire [(5'h14):(1'h0)] wire332;
  wire [(4'hc):(1'h0)] wire331;
  wire [(5'h14):(1'h0)] wire330;
  wire [(3'h6):(1'h0)] wire329;
  wire signed [(3'h7):(1'h0)] wire328;
  reg signed [(5'h13):(1'h0)] reg327 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire326;
  reg [(5'h12):(1'h0)] reg325 = (1'h0);
  reg signed [(4'he):(1'h0)] reg324 = (1'h0);
  reg [(2'h2):(1'h0)] reg323 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar322 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg321 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar320 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg319 = (1'h0);
  reg [(5'h10):(1'h0)] reg318 = (1'h0);
  reg [(5'h13):(1'h0)] reg317 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg316 = (1'h0);
  reg [(4'he):(1'h0)] forvar315 = (1'h0);
  reg [(4'h8):(1'h0)] reg314 = (1'h0);
  reg [(5'h11):(1'h0)] reg313 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg312 = (1'h0);
  reg [(3'h5):(1'h0)] reg311 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar310 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg307 = (1'h0);
  reg [(3'h6):(1'h0)] forvar306 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar305 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg304 = (1'h0);
  reg [(2'h2):(1'h0)] reg303 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar302 = (1'h0);
  reg [(5'h11):(1'h0)] reg301 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg300 = (1'h0);
  wire [(5'h12):(1'h0)] wire299;
  reg signed [(4'hf):(1'h0)] reg298 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg297 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg296 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg295 = (1'h0);
  reg [(5'h13):(1'h0)] reg294 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg293 = (1'h0);
  reg [(3'h6):(1'h0)] reg292 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar291 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg290 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg289 = (1'h0);
  reg signed [(4'he):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg287 = (1'h0);
  reg [(3'h4):(1'h0)] reg286 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg285 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg284 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar283 = (1'h0);
  reg [(4'hf):(1'h0)] reg282 = (1'h0);
  reg [(3'h5):(1'h0)] reg281 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire280;
  reg signed [(5'h14):(1'h0)] reg279 = (1'h0);
  reg [(3'h5):(1'h0)] reg278 = (1'h0);
  reg [(3'h7):(1'h0)] reg277 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg276 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg275 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg274 = (1'h0);
  reg [(4'hf):(1'h0)] forvar273 = (1'h0);
  reg [(4'h8):(1'h0)] reg272 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg271 = (1'h0);
  reg [(5'h12):(1'h0)] forvar270 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg269 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg268 = (1'h0);
  reg [(4'h8):(1'h0)] forvar267 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg266 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar265 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg264 = (1'h0);
  reg [(3'h5):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg262 = (1'h0);
  reg [(2'h3):(1'h0)] reg261 = (1'h0);
  reg [(5'h10):(1'h0)] reg260 = (1'h0);
  reg [(3'h6):(1'h0)] reg259 = (1'h0);
  reg [(4'hc):(1'h0)] reg258 = (1'h0);
  reg [(5'h14):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg256 = (1'h0);
  reg [(3'h5):(1'h0)] reg255 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar254 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg253 = (1'h0);
  reg [(4'hb):(1'h0)] reg252 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar251 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg250 = (1'h0);
  reg [(4'hf):(1'h0)] reg249 = (1'h0);
  reg [(4'hc):(1'h0)] reg248 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg247 = (1'h0);
  reg [(4'hb):(1'h0)] reg246 = (1'h0);
  reg [(5'h12):(1'h0)] forvar245 = (1'h0);
  reg [(2'h2):(1'h0)] reg244 = (1'h0);
  wire [(4'h9):(1'h0)] wire243;
  reg [(4'hb):(1'h0)] reg242 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg241 = (1'h0);
  reg [(4'hc):(1'h0)] reg240 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire239;
  wire signed [(5'h14):(1'h0)] wire238;
  assign y = {reg335,
                 wire334,
                 wire333,
                 wire332,
                 wire331,
                 wire330,
                 wire329,
                 wire328,
                 reg327,
                 wire326,
                 reg325,
                 reg324,
                 reg323,
                 forvar322,
                 reg321,
                 forvar320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 forvar315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 forvar310,
                 reg309,
                 reg308,
                 reg307,
                 forvar306,
                 forvar305,
                 reg304,
                 reg303,
                 forvar302,
                 reg301,
                 reg300,
                 wire299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 forvar291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 forvar283,
                 reg282,
                 reg281,
                 wire280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 forvar273,
                 reg272,
                 reg271,
                 forvar270,
                 reg269,
                 reg268,
                 forvar267,
                 reg266,
                 forvar265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 forvar254,
                 reg253,
                 reg252,
                 forvar251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 forvar245,
                 reg244,
                 wire243,
                 reg242,
                 reg241,
                 reg240,
                 wire239,
                 wire238,
                 (1'h0)};
  assign wire238 = $signed(wire237[(4'hc):(4'hc)]);
  assign wire239 = ($signed($signed(wire236[(3'h6):(2'h2)])) ?
                       (+wire234[(2'h2):(2'h2)]) : $signed(((+(wire236 ?
                           wire236 : wire235)) <= $unsigned((+wire234)))));
  always
    @(posedge clk) begin
      reg240 <= $unsigned((((8'hbd) << $unsigned((wire239 ?
              (8'ha8) : wire235))) ?
          $signed($signed(wire238[(2'h3):(1'h1)])) : wire239));
      reg241 = (-(+((+wire237) ?
          wire235 : ((reg240 ? wire239 : wire237) ?
              (~&reg240) : $unsigned(wire237)))));
      reg242 <= (((~|({wire239, wire238} & $signed(reg241))) ?
          $signed((~^(reg240 >>> (8'hbc)))) : wire238[(5'h12):(3'h6)]) >> wire237);
    end
  assign wire243 = ($signed(reg241[(3'h5):(3'h5)]) ?
                       wire238 : $unsigned({wire236[(3'h7):(2'h2)]}));
  always
    @(posedge clk) begin
      reg244 <= ({wire236, {{$signed(reg240)}, $signed($signed(wire234))}} ?
          (|wire239[(2'h2):(1'h1)]) : {{$signed((wire235 ? wire237 : reg241)),
                  reg242[(1'h0):(1'h0)]}});
      for (forvar245 = (1'h0); (forvar245 < (1'h0)); forvar245 = (forvar245 + (1'h1)))
        begin
          reg246 <= {$unsigned((^~($signed((8'hbe)) << {wire236})))};
          reg247 <= wire234;
          reg248 <= $unsigned(wire235);
          reg249 <= (|reg244);
        end
      reg250 <= ((8'h9e) << reg240);
    end
  always
    @(posedge clk) begin
      for (forvar251 = (1'h0); (forvar251 < (1'h0)); forvar251 = (forvar251 + (1'h1)))
        begin
          reg252 <= reg250;
          reg253 = reg249[(3'h7):(2'h2)];
          for (forvar254 = (1'h0); (forvar254 < (3'h4)); forvar254 = (forvar254 + (1'h1)))
            begin
              reg255 <= (((wire235[(3'h7):(2'h2)] ?
                          forvar254 : $signed($unsigned(reg248))) ?
                      (($unsigned(reg246) ?
                          (wire235 <= wire237) : forvar251) + {(reg250 ^~ wire237),
                          {wire235, reg240}}) : (!{wire235[(4'h9):(1'h0)],
                          (8'hb2)})) ?
                  (~^wire237[(2'h3):(1'h1)]) : $signed($unsigned(reg246)));
              reg256 = $unsigned($signed({$signed((8'hbd))}));
              reg257 <= wire238[(4'hd):(3'h6)];
              reg258 <= $signed((($unsigned((reg252 ? wire237 : reg252)) ?
                  {((8'hab) * reg255)} : $unsigned((reg244 ~^ reg242))) || reg252));
              reg259 <= {(8'h9e), $signed($signed(reg255))};
            end
          reg260 = reg259;
        end
      reg261 <= (!$signed(((^~$unsigned((8'hbd))) ^ {(reg259 ?
              wire238 : (7'h44))})));
      reg262 <= (^~reg244[(1'h0):(1'h0)]);
      reg263 <= (reg249 ?
          ({reg259[(3'h5):(2'h2)], (~(reg246 ? reg261 : reg256))} ?
              (wire234[(2'h3):(2'h2)] ?
                  $signed($unsigned(reg246)) : {(reg255 ~^ reg240),
                      (wire237 > forvar245)}) : $signed((~|wire236[(4'hc):(2'h2)]))) : reg249);
      reg264 <= $signed(reg247);
    end
  always
    @(posedge clk) begin
      for (forvar265 = (1'h0); (forvar265 < (2'h3)); forvar265 = (forvar265 + (1'h1)))
        begin
          reg266 = wire236;
          for (forvar267 = (1'h0); (forvar267 < (2'h3)); forvar267 = (forvar267 + (1'h1)))
            begin
              reg268 = reg240;
            end
          reg269 <= ($unsigned((^(~&$signed(reg263)))) <<< (forvar245 ^~ (+($unsigned(wire238) << reg268))));
          for (forvar270 = (1'h0); (forvar270 < (3'h4)); forvar270 = (forvar270 + (1'h1)))
            begin
              reg271 <= (&$unsigned({(reg259 ^~ (reg255 ?
                      reg269 : forvar265))}));
              reg272 <= (($signed(reg247[(4'h9):(3'h6)]) || $signed(forvar270)) ?
                  $signed(reg246) : reg257[(4'he):(2'h2)]);
            end
          for (forvar273 = (1'h0); (forvar273 < (2'h3)); forvar273 = (forvar273 + (1'h1)))
            begin
              reg274 <= (-forvar273);
              reg275 <= forvar270;
              reg276 <= {($unsigned((+$signed(reg269))) ?
                      $signed(((&reg258) || (&reg263))) : forvar245)};
              reg277 <= $signed($unsigned((reg255[(2'h3):(1'h1)] | $unsigned($signed((8'hb0))))));
              reg278 = {reg269[(4'hc):(2'h2)],
                  ((reg255[(1'h1):(1'h1)] == (reg248[(2'h2):(2'h2)] || reg260)) * (~$signed(forvar273)))};
            end
        end
      reg279 <= ({$signed(reg260[(4'ha):(3'h5)]),
              (wire237[(4'h9):(3'h7)] != reg249)} ?
          $signed(reg253[(1'h0):(1'h0)]) : wire234);
    end
  assign wire280 = reg248;
  always
    @(posedge clk) begin
      reg281 <= forvar254[(3'h7):(2'h3)];
      reg282 <= $signed({(^(~|$unsigned(wire280))),
          (&(-wire235[(3'h6):(1'h1)]))});
      for (forvar283 = (1'h0); (forvar283 < (2'h2)); forvar283 = (forvar283 + (1'h1)))
        begin
          reg284 <= $unsigned($signed(((forvar273 ?
                  forvar251 : $unsigned(reg266)) ?
              wire235[(1'h1):(1'h0)] : (((8'hb3) ? reg281 : wire235) ?
                  reg244[(1'h1):(1'h0)] : forvar283))));
          reg285 <= ((($unsigned((reg274 || wire236)) ?
              ($unsigned(wire243) ?
                  {wire280} : wire238) : (+$unsigned(reg271))) < reg247[(2'h3):(2'h2)]) || reg240);
          if (wire236[(3'h6):(3'h5)])
            begin
              reg286 <= (reg246 ?
                  $signed({(^~(reg249 ? (7'h41) : forvar270)),
                      reg274}) : $unsigned(wire236[(4'hb):(3'h5)]));
              reg287 <= $unsigned(reg285[(3'h7):(2'h2)]);
              reg288 <= reg250;
              reg289 <= (~^(~^$unsigned($signed(reg286[(2'h3):(2'h3)]))));
              reg290 <= (8'ha1);
            end
          else
            begin
              reg286 = ($signed(reg257) ?
                  ((reg253 ~^ $unsigned((reg246 ? reg242 : forvar265))) ?
                      $signed({reg244,
                          $signed(reg262)}) : (!{forvar245})) : ((8'hb9) ?
                      $unsigned($unsigned(reg257)) : ($signed({(8'hb6),
                              (7'h44)}) ?
                          reg263 : ($unsigned(reg248) ?
                              (&reg263) : {wire236, (8'hb2)}))));
              reg287 = reg261;
              reg288 = ({(8'h9e)} ?
                  $signed({$unsigned($signed(forvar251))}) : $signed({{reg252[(1'h0):(1'h0)]},
                      ($unsigned((8'hba)) ? (^reg286) : reg261)}));
            end
          for (forvar291 = (1'h0); (forvar291 < (2'h2)); forvar291 = (forvar291 + (1'h1)))
            begin
              reg292 = (reg258 << reg269);
              reg293 <= (8'hae);
              reg294 <= ($unsigned((~((wire243 & reg240) ?
                  (8'hbd) : $signed((8'ha8))))) + $unsigned((~&(|(^reg241)))));
              reg295 = reg240[(4'hb):(4'hb)];
              reg296 <= {($unsigned(($unsigned(reg246) <<< reg269)) * wire239[(4'hf):(4'hd)]),
                  (((&(reg266 ~^ reg289)) ?
                          forvar245 : $unsigned(reg284[(2'h2):(1'h1)])) ?
                      $unsigned($unsigned(forvar273[(4'hd):(1'h0)])) : {(!wire280[(1'h1):(1'h1)])})};
            end
        end
      reg297 <= (^($unsigned($unsigned((reg294 ? (8'haf) : wire234))) ?
          reg277[(1'h0):(1'h0)] : wire235));
    end
  always
    @(posedge clk) begin
      reg298 = (^$signed((reg292[(3'h5):(3'h5)] ?
          (reg281[(3'h4):(2'h2)] >= reg276[(3'h7):(3'h7)]) : ((reg255 ?
                  reg290 : reg285) ?
              (reg272 ? wire234 : reg274) : reg277[(1'h0):(1'h0)]))));
    end
  assign wire299 = (reg281 ?
                       (reg284[(3'h6):(2'h3)] - (((~&wire280) ?
                           $signed(wire236) : reg286) ^~ ($signed(reg240) ?
                           (~^reg248) : (!reg279)))) : ($unsigned((~{reg286,
                           wire234})) >= $unsigned($unsigned((+(8'ha9))))));
  always
    @(posedge clk) begin
      reg300 <= $signed(({reg279[(5'h13):(1'h0)], (|(reg285 << reg244))} ?
          {((reg296 * reg260) == (^~wire299))} : (^~$signed((|reg249)))));
      reg301 <= (forvar251[(4'hd):(4'hc)] ?
          {$signed((8'haf))} : (~$signed(reg297)));
    end
  always
    @(posedge clk) begin
      for (forvar302 = (1'h0); (forvar302 < (1'h0)); forvar302 = (forvar302 + (1'h1)))
        begin
          reg303 <= $unsigned($unsigned($unsigned(reg295)));
          reg304 <= reg287[(1'h0):(1'h0)];
        end
      for (forvar305 = (1'h0); (forvar305 < (1'h0)); forvar305 = (forvar305 + (1'h1)))
        begin
          for (forvar306 = (1'h0); (forvar306 < (2'h3)); forvar306 = (forvar306 + (1'h1)))
            begin
              reg307 <= reg279[(4'hf):(1'h1)];
              reg308 = $signed((($unsigned(reg266) << $unsigned(reg248[(4'h9):(1'h0)])) ?
                  $unsigned(reg264[(3'h4):(3'h4)]) : (^(8'haf))));
              reg309 = $signed((({(&reg242), (forvar273 <= reg296)} ?
                      (reg272 ?
                          $signed(reg287) : (reg244 & (8'h9e))) : ((8'ha0) ?
                          reg287[(3'h7):(3'h7)] : (|reg252))) ?
                  (^~(reg301 << reg253[(3'h4):(1'h0)])) : (reg281 && $unsigned((wire234 ?
                      wire236 : reg269)))));
            end
          for (forvar310 = (1'h0); (forvar310 < (1'h0)); forvar310 = (forvar310 + (1'h1)))
            begin
              reg311 <= (wire239 - wire238);
              reg312 <= wire239;
              reg313 <= (!((((~|(8'hb3)) ? reg297 : (|reg289)) ?
                  $signed(wire280) : $signed((reg297 ?
                      reg312 : reg241))) >= $signed($unsigned($unsigned((8'hb5))))));
            end
          reg314 <= reg259[(3'h4):(3'h4)];
          for (forvar315 = (1'h0); (forvar315 < (1'h0)); forvar315 = (forvar315 + (1'h1)))
            begin
              reg316 <= reg241[(4'h9):(3'h5)];
              reg317 <= $signed($signed(reg253[(2'h2):(1'h0)]));
            end
          reg318 <= ($signed($signed(reg264)) + ((~^$unsigned($signed(forvar310))) ^~ reg244[(1'h1):(1'h1)]));
        end
      reg319 <= $unsigned((reg271[(3'h6):(3'h4)] ? wire235 : reg258));
      for (forvar320 = (1'h0); (forvar320 < (2'h2)); forvar320 = (forvar320 + (1'h1)))
        begin
          reg321 <= reg298;
          for (forvar322 = (1'h0); (forvar322 < (3'h4)); forvar322 = (forvar322 + (1'h1)))
            begin
              reg323 <= {(((~(forvar305 ? (8'ha2) : (8'haf))) ?
                      {(forvar245 ? reg242 : forvar283),
                          {forvar315}} : {(reg249 ?
                              reg309 : reg253)}) + (reg271 >>> $unsigned(((8'h9d) == reg321)))),
                  ((-(~^$unsigned(reg252))) <= ((+$signed(reg293)) ?
                      reg311 : ((8'haa) | forvar245)))};
              reg324 <= ((!reg311[(2'h2):(1'h0)]) == (^$unsigned($signed(reg298))));
            end
          reg325 = {(reg264[(2'h3):(2'h3)] ?
                  ((!(reg271 ~^ reg314)) ?
                      (~|(~reg287)) : (-(reg241 <<< forvar254))) : ($signed((~^reg289)) ?
                      reg314[(3'h5):(1'h0)] : {$unsigned(reg272)})),
              (8'hb0)};
        end
    end
  assign wire326 = reg292[(2'h3):(1'h0)];
  always
    @(posedge clk) begin
      reg327 <= (|($signed($unsigned($unsigned(reg295))) ?
          $unsigned($unsigned(reg258[(4'h8):(2'h3)])) : reg272));
    end
  assign wire328 = $unsigned(((~&$unsigned((reg260 <= (8'hac)))) ?
                       $unsigned($signed({reg276,
                           reg325})) : (((wire326 < reg285) ?
                               $signed(reg290) : (forvar270 ^ reg325)) ?
                           ((wire234 ?
                               forvar306 : reg284) <<< (~|reg261)) : {$signed(reg260)})));
  assign wire329 = $unsigned(($signed(((~^reg247) ?
                       $unsigned(forvar302) : $signed(reg274))) >>> $unsigned((reg284[(3'h5):(3'h5)] > forvar291))));
  assign wire330 = reg272;
  assign wire331 = (reg313 ?
                       (&(~|wire243[(4'h8):(4'h8)])) : $signed(($unsigned(forvar305[(1'h1):(1'h1)]) * $unsigned($unsigned(reg255)))));
  assign wire332 = {(|$unsigned($unsigned((~(8'hbf)))))};
  assign wire333 = (+reg313);
  assign wire334 = $unsigned(reg327[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg335 <= $signed($signed($signed($signed($signed(forvar291)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module527  (y, clk, wire532, wire531, wire530, wire529, wire528);
  output wire [(32'h2d0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire532;
  input wire [(4'h9):(1'h0)] wire531;
  input wire signed [(5'h13):(1'h0)] wire530;
  input wire [(5'h12):(1'h0)] wire529;
  input wire [(5'h10):(1'h0)] wire528;
  wire [(2'h3):(1'h0)] wire598;
  reg [(3'h7):(1'h0)] reg597 = (1'h0);
  reg [(3'h5):(1'h0)] reg596 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg595 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg594 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire593;
  reg [(4'he):(1'h0)] reg592 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg591 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg590 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg589 = (1'h0);
  reg [(4'hd):(1'h0)] reg588 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar587 = (1'h0);
  reg [(4'hb):(1'h0)] reg586 = (1'h0);
  reg [(3'h6):(1'h0)] reg585 = (1'h0);
  reg [(4'h9):(1'h0)] reg584 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar583 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg582 = (1'h0);
  wire [(4'hb):(1'h0)] wire581;
  wire [(3'h5):(1'h0)] wire580;
  wire [(2'h2):(1'h0)] wire579;
  reg signed [(3'h7):(1'h0)] reg578 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg577 = (1'h0);
  reg [(4'he):(1'h0)] reg576 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg575 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg574 = (1'h0);
  reg [(5'h15):(1'h0)] forvar573 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar572 = (1'h0);
  reg [(4'hb):(1'h0)] reg571 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg570 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire569;
  reg signed [(5'h10):(1'h0)] reg568 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg567 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg566 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg565 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg564 = (1'h0);
  reg [(3'h4):(1'h0)] forvar563 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg562 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg561 = (1'h0);
  reg [(5'h10):(1'h0)] reg560 = (1'h0);
  reg [(4'hd):(1'h0)] reg559 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar558 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg557 = (1'h0);
  reg [(2'h3):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg555 = (1'h0);
  wire [(4'hf):(1'h0)] wire554;
  reg [(5'h15):(1'h0)] reg553 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg552 = (1'h0);
  reg [(5'h14):(1'h0)] reg551 = (1'h0);
  reg [(3'h4):(1'h0)] reg550 = (1'h0);
  reg [(5'h15):(1'h0)] reg549 = (1'h0);
  reg [(4'ha):(1'h0)] reg548 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg547 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar546 = (1'h0);
  reg [(4'hb):(1'h0)] reg545 = (1'h0);
  reg [(2'h3):(1'h0)] reg544 = (1'h0);
  wire [(4'hb):(1'h0)] wire543;
  wire signed [(5'h13):(1'h0)] wire542;
  wire [(4'h8):(1'h0)] wire541;
  wire [(4'h9):(1'h0)] wire540;
  wire signed [(5'h10):(1'h0)] wire539;
  wire [(5'h11):(1'h0)] wire538;
  reg signed [(5'h12):(1'h0)] reg537 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg536 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg535 = (1'h0);
  reg [(5'h12):(1'h0)] reg534 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg533 = (1'h0);
  assign y = {wire598,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 wire593,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 forvar587,
                 reg586,
                 reg585,
                 reg584,
                 forvar583,
                 reg582,
                 wire581,
                 wire580,
                 wire579,
                 reg578,
                 reg577,
                 reg576,
                 reg575,
                 reg574,
                 forvar573,
                 forvar572,
                 reg571,
                 reg570,
                 wire569,
                 reg568,
                 reg567,
                 reg566,
                 reg565,
                 reg564,
                 forvar563,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 forvar558,
                 reg557,
                 reg556,
                 reg555,
                 wire554,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 forvar546,
                 reg545,
                 reg544,
                 wire543,
                 wire542,
                 wire541,
                 wire540,
                 wire539,
                 wire538,
                 reg537,
                 reg536,
                 reg535,
                 reg534,
                 reg533,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg533 <= (($unsigned($signed(wire531)) | wire531[(3'h7):(3'h7)]) <<< (+(~|($signed(wire529) ?
          (wire530 ? wire532 : wire532) : wire528[(4'he):(3'h7)]))));
      reg534 <= wire528;
      reg535 = (wire530 << ($unsigned(reg533) - (wire529[(4'hb):(4'h8)] ?
          {(reg534 ? wire530 : wire530)} : reg533[(1'h0):(1'h0)])));
      reg536 <= ($signed({$signed(((8'ha2) ? wire530 : wire531))}) ?
          reg535[(1'h0):(1'h0)] : $signed((((wire532 ? wire531 : wire528) ?
                  reg535[(2'h3):(2'h2)] : $signed(reg534)) ?
              wire528 : $unsigned(wire531[(1'h0):(1'h0)]))));
      reg537 = {$signed(wire530), reg535[(1'h0):(1'h0)]};
    end
  assign wire538 = $signed(reg533);
  assign wire539 = reg535[(3'h6):(2'h2)];
  assign wire540 = (^~({reg537[(4'hc):(4'ha)]} != (+$unsigned((wire528 - wire531)))));
  assign wire541 = $unsigned(reg535);
  assign wire542 = wire532;
  assign wire543 = wire529;
  always
    @(posedge clk) begin
      reg544 <= wire531[(3'h5):(2'h2)];
      reg545 <= ((|(|wire541)) + ((((wire530 ?
              wire543 : reg537) - wire530) >> ((&wire532) ^~ (|wire532))) ?
          (((&wire539) ?
              {wire531,
                  (8'ha3)} : {(8'hbd)}) > $unsigned($unsigned(reg537))) : ($signed($unsigned((8'haa))) * (-reg533[(1'h0):(1'h0)]))));
      for (forvar546 = (1'h0); (forvar546 < (2'h3)); forvar546 = (forvar546 + (1'h1)))
        begin
          reg547 = wire538[(4'h9):(2'h2)];
          reg548 = (reg547[(4'hc):(1'h0)] ?
              (reg533 ?
                  reg533[(1'h0):(1'h0)] : {reg533,
                      $unsigned($signed((8'ha6)))}) : (+$unsigned($unsigned($signed((8'hbf))))));
        end
      reg549 <= (^$unsigned((reg536 & ((wire528 | wire541) ^~ (8'hac)))));
      reg550 <= wire542[(1'h1):(1'h1)];
    end
  always
    @(posedge clk) begin
      reg551 <= wire529[(4'h8):(3'h4)];
      reg552 <= (|{reg549, (|(^~(wire531 <= wire528)))});
    end
  always
    @(posedge clk) begin
      reg553 <= $unsigned((reg547[(4'hf):(3'h5)] >= (~&(wire531[(2'h2):(1'h0)] ?
          wire541[(1'h1):(1'h1)] : $unsigned(reg536)))));
    end
  assign wire554 = $signed($unsigned($signed($signed((reg537 ?
                       wire538 : wire532)))));
  always
    @(posedge clk) begin
      reg555 <= ((~&reg550[(1'h0):(1'h0)]) != $signed((^$signed((reg553 || wire540)))));
      reg556 = wire539;
      reg557 = $unsigned(reg534);
      for (forvar558 = (1'h0); (forvar558 < (2'h2)); forvar558 = (forvar558 + (1'h1)))
        begin
          reg559 <= (^wire530);
          reg560 = reg549;
          reg561 <= reg534[(3'h7):(1'h0)];
          reg562 <= reg537[(4'hc):(2'h3)];
          for (forvar563 = (1'h0); (forvar563 < (1'h0)); forvar563 = (forvar563 + (1'h1)))
            begin
              reg564 <= wire543;
              reg565 <= (~{(reg561[(3'h6):(3'h4)] ?
                      (7'h43) : ((-(8'hb4)) <<< ((8'h9c) || (8'hb9)))),
                  (^~forvar546)});
              reg566 <= $unsigned(reg537);
              reg567 <= $unsigned(wire531[(2'h3):(2'h3)]);
              reg568 <= reg556[(1'h0):(1'h0)];
            end
        end
    end
  assign wire569 = $unsigned($signed(reg533));
  always
    @(posedge clk) begin
      reg570 = (wire569[(3'h6):(1'h1)] ?
          wire541 : ((($signed((8'hb0)) ? (+wire531) : (wire538 < wire539)) ?
              $signed(wire532[(3'h7):(1'h0)]) : (reg533 ?
                  (wire531 ? reg557 : reg544) : ((8'ha3) ?
                      (8'hb0) : reg548))) ~^ $unsigned((wire531[(1'h0):(1'h0)] ?
              (reg533 ? (8'ha9) : forvar546) : wire540))));
      reg571 <= $unsigned((reg562 || (!reg556)));
      for (forvar572 = (1'h0); (forvar572 < (3'h4)); forvar572 = (forvar572 + (1'h1)))
        begin
          for (forvar573 = (1'h0); (forvar573 < (3'h4)); forvar573 = (forvar573 + (1'h1)))
            begin
              reg574 <= $signed(($signed(({reg544} ?
                      (reg549 ? (8'hbb) : forvar563) : (reg544 | (8'h9d)))) ?
                  {((wire529 || wire539) || $unsigned(forvar573)),
                      forvar558[(3'h4):(2'h3)]} : reg557[(1'h1):(1'h0)]));
              reg575 <= $unsigned(wire539);
              reg576 <= $unsigned($signed((8'ha1)));
              reg577 = (!reg548[(2'h2):(1'h0)]);
            end
        end
      reg578 <= (reg551[(4'hd):(1'h0)] ?
          (wire542[(1'h0):(1'h0)] ?
              {reg544,
                  reg544} : $unsigned(forvar563[(1'h1):(1'h0)])) : {($unsigned($signed(forvar558)) ?
                  $signed($unsigned(forvar546)) : $unsigned(reg577))});
    end
  assign wire579 = (8'hae);
  assign wire580 = $unsigned({(($signed(reg560) ?
                           (wire554 ?
                               (8'hba) : wire530) : $signed(wire530)) >> $unsigned((&reg552)))});
  assign wire581 = reg534;
  always
    @(posedge clk) begin
      reg582 <= (({{$unsigned((8'hab))}} ?
          reg537[(5'h11):(3'h7)] : (~&reg567)) != reg535);
      for (forvar583 = (1'h0); (forvar583 < (1'h1)); forvar583 = (forvar583 + (1'h1)))
        begin
          reg584 <= ($unsigned((~&reg570)) & reg550[(1'h1):(1'h1)]);
          reg585 = (~^$signed($unsigned({$signed(wire543),
              $unsigned(wire542)})));
          reg586 <= $unsigned($unsigned({forvar546[(2'h3):(2'h2)]}));
          for (forvar587 = (1'h0); (forvar587 < (2'h2)); forvar587 = (forvar587 + (1'h1)))
            begin
              reg588 = ($signed(((~&(wire532 ~^ wire540)) ?
                  (forvar563 >>> reg535[(3'h5):(2'h3)]) : (reg562 ^~ (forvar546 ?
                      reg545 : reg537)))) < (reg551 << forvar583));
              reg589 <= ((~&$signed((~|(+forvar573)))) >> $unsigned(reg557[(1'h1):(1'h0)]));
              reg590 = reg565;
            end
          reg591 <= forvar587[(2'h2):(2'h2)];
        end
      reg592 = (~|$unsigned($unsigned(wire581)));
    end
  assign wire593 = reg551[(4'hf):(4'hf)];
  always
    @(posedge clk) begin
      reg594 <= $signed(reg537);
      reg595 = $unsigned(reg550[(2'h2):(2'h2)]);
      reg596 = ($unsigned(reg560[(5'h10):(4'hc)]) ?
          {(~^$unsigned($signed(reg585))),
              {((^~reg535) ?
                      {(8'h9f)} : (wire542 | reg550))}} : $unsigned((~{(8'ha5)})));
    end
  always
    @(posedge clk) begin
      reg597 <= $unsigned((8'h9e));
    end
  assign wire598 = {(($unsigned(wire531) ~^ ($signed((8'ha1)) ?
                               (reg575 == wire579) : (!reg559))) ?
                           $unsigned({{(7'h41),
                                   wire528}}) : ((~|$unsigned(forvar563)) ?
                               $signed({forvar546}) : $unsigned((reg535 || (8'hb6)))))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module629
#( parameter param706 = (((({(8'ha7), (7'h44)} ? ((7'h40) | (8'hbf)) : (+(8'h9c))) - (((8'hb0) <= (8'hab)) ? {(8'hb8), (8'hbb)} : {(8'hbc), (8'haa)})) & ((((8'hba) ? (8'hb0) : (8'ha1)) ? (|(8'ha7)) : ((8'hb9) ? (8'hbe) : (8'ha4))) << (~&{(8'ha4), (8'hb9)}))) == ((({(8'ha7)} ? ((8'hb8) ? (8'haa) : (8'hab)) : (-(8'hb3))) <= ({(8'hb1), (8'hb9)} ? {(7'h42), (8'hbd)} : ((8'ha3) >> (8'haf)))) ? (8'ha7) : (8'hb9))) )
(y, clk, wire634, wire633, wire632, wire631, wire630);
  output wire [(32'h312):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire634;
  input wire [(2'h3):(1'h0)] wire633;
  input wire [(4'hf):(1'h0)] wire632;
  input wire [(4'hb):(1'h0)] wire631;
  input wire signed [(2'h3):(1'h0)] wire630;
  wire [(3'h5):(1'h0)] wire705;
  reg signed [(5'h13):(1'h0)] reg704 = (1'h0);
  reg [(4'hb):(1'h0)] forvar703 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg702 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire701;
  wire [(5'h12):(1'h0)] wire700;
  wire signed [(2'h3):(1'h0)] wire699;
  wire [(5'h10):(1'h0)] wire698;
  reg [(4'hd):(1'h0)] reg697 = (1'h0);
  reg [(3'h4):(1'h0)] reg696 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg695 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg694 = (1'h0);
  reg [(4'ha):(1'h0)] reg693 = (1'h0);
  reg [(4'h8):(1'h0)] reg692 = (1'h0);
  reg [(5'h11):(1'h0)] reg691 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg690 = (1'h0);
  reg [(5'h11):(1'h0)] reg689 = (1'h0);
  reg signed [(4'he):(1'h0)] reg688 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg687 = (1'h0);
  reg [(5'h11):(1'h0)] reg686 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg685 = (1'h0);
  reg [(3'h5):(1'h0)] reg684 = (1'h0);
  wire [(5'h13):(1'h0)] wire683;
  wire [(5'h14):(1'h0)] wire682;
  reg [(4'h8):(1'h0)] reg681 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg680 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg679 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg678 = (1'h0);
  reg [(3'h6):(1'h0)] reg677 = (1'h0);
  reg [(5'h11):(1'h0)] reg676 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar675 = (1'h0);
  wire [(3'h6):(1'h0)] wire674;
  reg [(3'h7):(1'h0)] reg673 = (1'h0);
  reg [(3'h7):(1'h0)] reg672 = (1'h0);
  reg [(4'hb):(1'h0)] reg671 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg670 = (1'h0);
  reg [(4'h8):(1'h0)] reg669 = (1'h0);
  reg [(5'h10):(1'h0)] reg668 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg667 = (1'h0);
  reg [(2'h3):(1'h0)] reg666 = (1'h0);
  reg [(4'ha):(1'h0)] forvar665 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar664 = (1'h0);
  reg signed [(4'he):(1'h0)] reg663 = (1'h0);
  reg [(3'h4):(1'h0)] reg662 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire661;
  reg signed [(4'hf):(1'h0)] reg660 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg659 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg658 = (1'h0);
  reg [(2'h3):(1'h0)] reg657 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire656;
  reg [(3'h7):(1'h0)] reg655 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg654 = (1'h0);
  reg [(2'h2):(1'h0)] forvar653 = (1'h0);
  reg [(4'h9):(1'h0)] reg652 = (1'h0);
  reg [(3'h6):(1'h0)] reg651 = (1'h0);
  reg [(2'h3):(1'h0)] reg650 = (1'h0);
  reg [(4'hd):(1'h0)] reg649 = (1'h0);
  reg [(3'h5):(1'h0)] reg648 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire647;
  reg [(3'h7):(1'h0)] reg646 = (1'h0);
  reg [(5'h14):(1'h0)] reg645 = (1'h0);
  reg [(2'h2):(1'h0)] reg643 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg640 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar639 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg644 = (1'h0);
  reg [(5'h13):(1'h0)] forvar643 = (1'h0);
  reg [(5'h12):(1'h0)] reg642 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg641 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar640 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg639 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg638 = (1'h0);
  reg [(3'h7):(1'h0)] reg637 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg636 = (1'h0);
  wire [(5'h14):(1'h0)] wire635;
  assign y = {wire705,
                 reg704,
                 forvar703,
                 reg702,
                 wire701,
                 wire700,
                 wire699,
                 wire698,
                 reg697,
                 reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 reg691,
                 reg690,
                 reg689,
                 reg688,
                 reg687,
                 reg686,
                 reg685,
                 reg684,
                 wire683,
                 wire682,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 reg676,
                 forvar675,
                 wire674,
                 reg673,
                 reg672,
                 reg671,
                 reg670,
                 reg669,
                 reg668,
                 reg667,
                 reg666,
                 forvar665,
                 forvar664,
                 reg663,
                 reg662,
                 wire661,
                 reg660,
                 reg659,
                 reg658,
                 reg657,
                 wire656,
                 reg655,
                 reg654,
                 forvar653,
                 reg652,
                 reg651,
                 reg650,
                 reg649,
                 reg648,
                 wire647,
                 reg646,
                 reg645,
                 reg643,
                 reg640,
                 forvar639,
                 reg644,
                 forvar643,
                 reg642,
                 reg641,
                 forvar640,
                 reg639,
                 reg638,
                 reg637,
                 reg636,
                 wire635,
                 (1'h0)};
  assign wire635 = wire631[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg636 <= (!(~|($signed((!wire635)) ? wire635 : $unsigned({(8'hb9)}))));
      reg637 = (wire635[(5'h14):(2'h2)] ?
          $unsigned($signed(((~wire630) * {(8'h9c),
              wire634}))) : $unsigned((reg636[(4'ha):(4'h9)] >> $signed((wire635 ?
              wire633 : wire635)))));
      reg638 = (~&wire631[(3'h6):(2'h3)]);
    end
  always
    @(posedge clk) begin
      if ($signed(wire633))
        begin
          reg639 <= $unsigned(reg636);
          for (forvar640 = (1'h0); (forvar640 < (3'h4)); forvar640 = (forvar640 + (1'h1)))
            begin
              reg641 <= (|(^reg638));
              reg642 = (~$signed((($unsigned(wire634) ?
                  forvar640 : wire630) >>> (((8'ha0) ? reg639 : wire632) ?
                  (forvar640 << reg641) : reg641))));
            end
          for (forvar643 = (1'h0); (forvar643 < (1'h1)); forvar643 = (forvar643 + (1'h1)))
            begin
              reg644 <= (~&(forvar643[(4'h9):(4'h9)] ?
                  reg641 : $signed($signed((reg641 ? (7'h41) : forvar640)))));
            end
        end
      else
        begin
          for (forvar639 = (1'h0); (forvar639 < (2'h2)); forvar639 = (forvar639 + (1'h1)))
            begin
              reg640 <= (|$signed((&$unsigned(wire630[(2'h2):(2'h2)]))));
              reg641 <= reg638;
              reg642 <= ((~&(wire635 != (8'hb2))) >>> (8'haa));
              reg643 <= (-{(-(^(wire633 + (8'ha7))))});
            end
        end
      reg645 = ((!(($signed(reg639) <<< forvar639) ?
              $signed($signed(reg639)) : reg640)) ?
          ((|((~&wire634) >> (reg642 + wire630))) > ((~^$unsigned((8'hb5))) ~^ (+wire632))) : (wire634[(1'h1):(1'h0)] + $signed($signed((forvar640 ?
              wire635 : wire630)))));
      reg646 <= forvar639;
    end
  assign wire647 = (!$signed((($unsigned(forvar643) ?
                           reg642[(4'he):(1'h0)] : reg644[(1'h0):(1'h0)]) ?
                       forvar643 : (&{reg641}))));
  always
    @(posedge clk) begin
      reg648 <= reg636[(4'h9):(3'h5)];
      reg649 <= (((~{(forvar639 >>> wire634),
          (~^reg641)}) || $signed($unsigned($signed(reg644)))) >>> $unsigned(wire632[(4'hb):(3'h6)]));
      reg650 <= (!($signed(((forvar640 ? reg644 : wire631) ?
              ((8'had) ? reg646 : reg640) : (reg646 >>> reg640))) ?
          $unsigned((reg638 ^ reg645)) : $signed((~&$unsigned(reg637)))));
    end
  always
    @(posedge clk) begin
      reg651 <= ((|({(8'hb9)} ?
          {wire632[(2'h2):(2'h2)],
              wire631} : wire630[(2'h3):(1'h0)])) || (&(-forvar640[(2'h3):(1'h0)])));
      reg652 <= $signed($signed($unsigned((wire635[(4'hf):(4'hb)] >> $signed((8'ha1))))));
      for (forvar653 = (1'h0); (forvar653 < (3'h4)); forvar653 = (forvar653 + (1'h1)))
        begin
          reg654 = (!reg649);
          reg655 <= $signed($unsigned(reg648[(1'h0):(1'h0)]));
        end
    end
  assign wire656 = {(-reg638[(1'h1):(1'h1)])};
  always
    @(posedge clk) begin
      reg657 <= wire635;
      reg658 <= $unsigned((($signed(reg655) ?
              ($signed((8'h9f)) ^ (8'h9d)) : $unsigned(wire634)) ?
          {(reg655[(1'h0):(1'h0)] ?
                  reg642[(5'h12):(4'he)] : reg639[(1'h1):(1'h0)]),
              forvar643} : $signed((reg642[(2'h3):(2'h3)] <= (reg649 & reg644)))));
      reg659 <= $signed((~|(~|$unsigned(forvar643[(1'h0):(1'h0)]))));
    end
  always
    @(posedge clk) begin
      reg660 <= (reg658[(1'h1):(1'h0)] ? reg646[(3'h4):(2'h2)] : wire630);
    end
  assign wire661 = reg657[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg662 = $unsigned(({((~|forvar639) ? (reg636 ~^ reg649) : {reg636}),
          reg657} | {reg650, reg648[(2'h3):(1'h1)]}));
      reg663 = $signed($unsigned(((reg654 != $unsigned(reg643)) ~^ (reg652 >= (reg637 <<< (8'h9d))))));
      for (forvar664 = (1'h0); (forvar664 < (2'h2)); forvar664 = (forvar664 + (1'h1)))
        begin
          for (forvar665 = (1'h0); (forvar665 < (3'h4)); forvar665 = (forvar665 + (1'h1)))
            begin
              reg666 <= {$signed(((^~reg648) ?
                      (~&(8'hb1)) : ((~(8'h9d)) >>> $unsigned(forvar665))))};
              reg667 <= $signed((!($signed($unsigned((8'ha6))) & (^~(~&(8'hab))))));
              reg668 <= (^(reg651[(1'h1):(1'h1)] ?
                  (|$unsigned({reg655})) : wire656[(2'h3):(1'h1)]));
              reg669 <= $unsigned($unsigned($signed(($unsigned(reg652) ~^ (reg648 >= reg663)))));
              reg670 <= ($unsigned($unsigned(wire631)) && reg650[(2'h3):(2'h2)]);
            end
          reg671 <= $unsigned($signed($signed($unsigned((~^wire647)))));
        end
      reg672 <= reg660[(1'h0):(1'h0)];
      reg673 <= wire632;
    end
  assign wire674 = wire632;
  always
    @(posedge clk) begin
      for (forvar675 = (1'h0); (forvar675 < (2'h2)); forvar675 = (forvar675 + (1'h1)))
        begin
          if ((wire656[(1'h1):(1'h0)] ?
              $unsigned(reg672[(3'h7):(2'h3)]) : reg663))
            begin
              reg676 <= {wire633[(1'h1):(1'h0)]};
              reg677 <= (8'haa);
            end
          else
            begin
              reg676 <= (+(^~reg667[(3'h7):(3'h7)]));
            end
          if ((($signed(((~&(7'h41)) ?
              (^reg677) : (~|(8'hab)))) & $signed($unsigned($unsigned(reg637)))) + (~$unsigned($signed(forvar640)))))
            begin
              reg678 <= {reg667[(4'hb):(3'h4)],
                  $signed(((|(wire632 ? forvar665 : reg668)) ?
                      (reg654 == ((8'hb2) - reg636)) : reg646[(3'h5):(3'h5)]))};
              reg679 <= forvar664;
            end
          else
            begin
              reg678 <= ($signed((wire632 ?
                      {(wire661 ? wire632 : wire635)} : reg671)) ?
                  reg640 : ((wire633[(1'h0):(1'h0)] << $unsigned((reg679 ?
                      reg642 : reg673))) | $signed(reg659)));
              reg679 = $unsigned(((~|$unsigned((^~forvar675))) ?
                  $unsigned(wire674) : (reg640 ?
                      reg663 : $signed((wire634 >= (8'ha7))))));
            end
          reg680 <= (^reg666[(2'h3):(1'h0)]);
          reg681 = {((~forvar653) ? reg650[(2'h2):(1'h1)] : $unsigned(reg636)),
              (wire661[(4'hf):(2'h2)] ?
                  (|((reg666 ^ reg641) ?
                      (reg669 ?
                          forvar643 : reg655) : $unsigned(wire630))) : reg678)};
        end
    end
  assign wire682 = (forvar664 ?
                       {reg636[(3'h5):(2'h2)],
                           $unsigned(reg638[(1'h1):(1'h0)])} : reg678);
  assign wire683 = $unsigned({reg673});
  always
    @(posedge clk) begin
      reg684 = (wire631 ?
          $signed(((((8'hb6) ? reg667 : reg639) ?
              reg667 : reg636) <= ($unsigned(reg680) ?
              (reg636 - forvar639) : $unsigned(reg648)))) : (!reg666));
      reg685 = (7'h44);
      reg686 <= (-(reg636[(4'hb):(3'h7)] ?
          reg655[(3'h4):(2'h2)] : ($signed((~|wire634)) || (~^$unsigned(reg652)))));
      reg687 = ({$unsigned($unsigned($signed(reg663)))} ?
          $signed(((-(reg685 + wire633)) ?
              $signed(reg658) : reg648[(2'h3):(2'h2)])) : (~(((wire635 <<< forvar640) - (wire635 ?
              forvar639 : reg667)) - $unsigned((reg645 <<< reg636)))));
    end
  always
    @(posedge clk) begin
      if (reg659[(2'h3):(2'h2)])
        begin
          reg688 <= reg669[(3'h4):(2'h3)];
        end
      else
        begin
          reg688 = $signed(reg667[(2'h3):(1'h0)]);
          reg689 <= {$unsigned(reg659[(3'h6):(2'h2)]),
              ((($signed(reg688) <<< (reg670 <= wire661)) ?
                      {wire631[(4'h8):(1'h0)], reg673} : (|((8'ha2) ?
                          reg676 : reg641))) ?
                  {(~|(^(8'ha4))),
                      wire683[(4'hf):(2'h3)]} : $signed(($unsigned(forvar653) ~^ $unsigned(reg638))))};
          if (({$signed({wire634[(3'h6):(3'h4)]})} >= (~&(reg659 && (!(|reg666))))))
            begin
              reg690 <= $unsigned((+(~&{$signed(reg678), reg655})));
              reg691 <= reg649[(2'h2):(1'h0)];
              reg692 <= (forvar675 >> (~((~(reg648 >>> reg684)) ?
                  reg663[(2'h3):(2'h3)] : reg652)));
              reg693 <= $signed(reg639[(4'he):(4'h9)]);
              reg694 <= $unsigned(($unsigned(reg650[(2'h3):(1'h0)]) >> (reg657[(1'h1):(1'h0)] >> wire634[(2'h2):(1'h1)])));
            end
          else
            begin
              reg690 <= ($signed($unsigned($unsigned($signed(reg652)))) & reg660[(2'h3):(2'h3)]);
              reg691 <= (($signed((!(&reg638))) + reg651[(1'h1):(1'h0)]) ?
                  $unsigned(($signed($unsigned(reg680)) ?
                      {(reg636 && reg686)} : ((reg657 ^~ (8'ha6)) ?
                          $unsigned((8'hb0)) : wire647[(4'hf):(4'hf)]))) : $signed(({(-reg640),
                          $unsigned(wire634)} ?
                      (+$signed(forvar665)) : reg640[(4'ha):(4'h8)])));
              reg692 <= {($signed($unsigned(reg648)) ~^ $signed($signed(reg679[(4'h9):(2'h3)])))};
              reg693 <= forvar675;
            end
          reg695 = {reg672[(2'h2):(1'h1)]};
        end
      reg696 = $unsigned(($unsigned((&$unsigned(reg695))) ?
          $signed(reg691[(4'he):(4'hc)]) : reg691));
      reg697 <= reg694[(3'h4):(1'h0)];
    end
  assign wire698 = (((reg693[(1'h1):(1'h0)] ?
                               {$signed(reg687)} : ((reg681 ^ reg637) ?
                                   reg637 : forvar665[(3'h6):(1'h1)])) ?
                           reg662 : reg660) ?
                       $unsigned(((-reg684[(1'h1):(1'h1)]) << $signed(forvar665[(1'h0):(1'h0)]))) : ($unsigned(reg676) ?
                           (reg651 + {(forvar653 ^~ (8'ha2))}) : (({wire633} <<< $signed(reg679)) ?
                               ((wire630 || reg669) || reg669[(3'h5):(1'h1)]) : (reg655[(3'h5):(1'h1)] ~^ (wire661 ?
                                   reg691 : reg681)))));
  assign wire699 = (8'hb2);
  assign wire700 = reg688[(4'h9):(2'h2)];
  assign wire701 = reg692;
  always
    @(posedge clk) begin
      reg702 = $signed(wire699[(1'h0):(1'h0)]);
      for (forvar703 = (1'h0); (forvar703 < (2'h3)); forvar703 = (forvar703 + (1'h1)))
        begin
          reg704 <= $signed($unsigned((~^$unsigned((reg660 - reg663)))));
        end
    end
  assign wire705 = (^~$signed(reg693));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module788
#( parameter param838 = (((^({(8'hab), (8'ha8)} < (8'h9c))) ^~ ((~&((8'hbf) == (8'hb6))) | (((8'ha7) ? (8'hbd) : (7'h42)) + (-(8'ha8))))) ^~ (((((8'haa) ^ (8'ha0)) != ((8'ha6) ? (8'hae) : (8'ha9))) ? {(!(8'hab)), ((8'hbf) & (8'h9d))} : ((|(8'ha9)) ? ((8'hb9) ? (8'ha7) : (8'hbe)) : ((8'ha8) ^ (8'haa)))) ? {(8'had), (((7'h41) - (8'ha8)) >>> (|(8'ha3)))} : (-{{(7'h44), (7'h40)}, ((8'hbd) && (8'hbf))})))
, parameter param839 = ((^~(((param838 ^ param838) ? (8'h9c) : (|param838)) ^~ param838)) ? param838 : (~|param838)) )
(y, clk, wire793, wire792, wire791, wire790, wire789);
  output wire [(32'h1ee):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire793;
  input wire signed [(2'h2):(1'h0)] wire792;
  input wire [(2'h2):(1'h0)] wire791;
  input wire signed [(4'he):(1'h0)] wire790;
  input wire [(2'h3):(1'h0)] wire789;
  reg [(4'hc):(1'h0)] reg837 = (1'h0);
  reg [(2'h3):(1'h0)] reg836 = (1'h0);
  reg [(3'h6):(1'h0)] reg835 = (1'h0);
  reg [(3'h5):(1'h0)] reg834 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg833 = (1'h0);
  reg [(4'he):(1'h0)] reg832 = (1'h0);
  reg signed [(4'he):(1'h0)] reg831 = (1'h0);
  reg [(4'hd):(1'h0)] reg830 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg829 = (1'h0);
  reg [(4'hf):(1'h0)] reg828 = (1'h0);
  reg [(3'h5):(1'h0)] reg827 = (1'h0);
  wire [(4'ha):(1'h0)] wire826;
  reg signed [(4'h8):(1'h0)] reg825 = (1'h0);
  reg [(3'h7):(1'h0)] reg824 = (1'h0);
  reg [(4'h9):(1'h0)] forvar823 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg822 = (1'h0);
  reg [(4'hb):(1'h0)] reg821 = (1'h0);
  reg [(4'he):(1'h0)] reg820 = (1'h0);
  reg [(4'hc):(1'h0)] reg819 = (1'h0);
  reg [(4'hb):(1'h0)] forvar818 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar817 = (1'h0);
  reg [(3'h7):(1'h0)] reg816 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg815 = (1'h0);
  reg [(3'h7):(1'h0)] reg814 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg813 = (1'h0);
  reg [(4'hc):(1'h0)] reg812 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar811 = (1'h0);
  reg [(5'h13):(1'h0)] forvar810 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg809 = (1'h0);
  reg [(5'h10):(1'h0)] reg808 = (1'h0);
  reg [(4'h8):(1'h0)] forvar807 = (1'h0);
  wire [(4'h8):(1'h0)] wire806;
  wire signed [(3'h7):(1'h0)] wire805;
  reg signed [(4'hd):(1'h0)] reg804 = (1'h0);
  wire [(4'hc):(1'h0)] wire803;
  reg signed [(4'hd):(1'h0)] reg802 = (1'h0);
  reg [(5'h15):(1'h0)] reg801 = (1'h0);
  reg [(4'h8):(1'h0)] reg800 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg799 = (1'h0);
  reg [(5'h12):(1'h0)] reg798 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire797;
  wire signed [(5'h10):(1'h0)] wire796;
  wire signed [(5'h10):(1'h0)] wire795;
  wire signed [(5'h11):(1'h0)] wire794;
  assign y = {reg837,
                 reg836,
                 reg835,
                 reg834,
                 reg833,
                 reg832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 reg827,
                 wire826,
                 reg825,
                 reg824,
                 forvar823,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 forvar818,
                 forvar817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 reg812,
                 forvar811,
                 forvar810,
                 reg809,
                 reg808,
                 forvar807,
                 wire806,
                 wire805,
                 reg804,
                 wire803,
                 reg802,
                 reg801,
                 reg800,
                 reg799,
                 reg798,
                 wire797,
                 wire796,
                 wire795,
                 wire794,
                 (1'h0)};
  assign wire794 = $signed({$signed({wire792, wire790[(4'hc):(1'h0)]}),
                       (((wire790 && wire790) ?
                           (~^wire793) : ((8'haf) <= wire793)) || $signed({wire791,
                           wire793}))});
  assign wire795 = (wire792 ?
                       ((wire791[(2'h2):(2'h2)] >>> $unsigned((wire791 || (8'hb6)))) ?
                           (|wire790) : {{$signed(wire792),
                                   (wire792 ? wire794 : wire790)},
                               (&$unsigned(wire790))}) : wire790);
  assign wire796 = $unsigned(wire793);
  assign wire797 = $unsigned($unsigned(($unsigned((~&wire791)) ^~ $signed((wire791 << (8'hae))))));
  always
    @(posedge clk) begin
      reg798 <= (^(|$unsigned(((+wire793) * (^wire793)))));
      reg799 <= wire795[(4'hf):(4'hc)];
      reg800 <= ({(($unsigned(wire790) ? wire790 : wire795) ?
              ($signed(reg799) ?
                  (^~wire789) : $signed(reg798)) : $unsigned({wire797,
                  wire791}))} > wire789[(1'h0):(1'h0)]);
      reg801 <= ((wire797[(3'h6):(2'h3)] ?
          (^(|(wire789 && wire789))) : (8'ha2)) ^~ {($unsigned($unsigned(wire791)) ?
              $unsigned(reg798[(4'he):(3'h4)]) : reg799)});
      reg802 <= reg800[(2'h3):(2'h2)];
    end
  assign wire803 = (((reg798[(4'hb):(3'h5)] << ($unsigned(wire797) ?
                           (reg802 ?
                               reg798 : reg799) : $unsigned(wire796))) <<< wire792) ?
                       $unsigned($signed($unsigned((reg798 * (7'h43))))) : ((&((wire795 ?
                                   wire792 : (8'hb8)) ?
                               {reg799, wire797} : (&reg801))) ?
                           $unsigned((8'h9f)) : {(8'hb9), (~$signed(reg799))}));
  always
    @(posedge clk) begin
      reg804 = wire795;
    end
  assign wire805 = wire795;
  assign wire806 = $unsigned($signed((8'ha8)));
  always
    @(posedge clk) begin
      for (forvar807 = (1'h0); (forvar807 < (1'h0)); forvar807 = (forvar807 + (1'h1)))
        begin
          reg808 = reg798[(5'h10):(1'h1)];
          reg809 <= ((-$signed(($unsigned(wire793) & (wire791 ?
                  wire805 : reg800)))) ?
              wire794 : $unsigned(reg804));
        end
      for (forvar810 = (1'h0); (forvar810 < (1'h0)); forvar810 = (forvar810 + (1'h1)))
        begin
          for (forvar811 = (1'h0); (forvar811 < (3'h4)); forvar811 = (forvar811 + (1'h1)))
            begin
              reg812 <= wire805;
              reg813 <= (wire791 && $signed($unsigned($unsigned((wire797 ?
                  forvar807 : (8'hb2))))));
              reg814 = reg799;
            end
        end
      reg815 <= $unsigned(((((&forvar811) ?
          {reg813} : forvar811[(3'h7):(2'h3)]) ^~ $unsigned((reg812 ?
          wire795 : wire796))) ^ (^{(~reg813), $signed(wire796)})));
      reg816 <= (~$signed((~^$signed((wire796 && wire796)))));
      for (forvar817 = (1'h0); (forvar817 < (3'h4)); forvar817 = (forvar817 + (1'h1)))
        begin
          for (forvar818 = (1'h0); (forvar818 < (2'h3)); forvar818 = (forvar818 + (1'h1)))
            begin
              reg819 = {(wire806 ?
                      $unsigned($unsigned((~^wire791))) : (&$signed($signed(reg812))))};
              reg820 <= ((~$signed((wire806 ?
                  (!(8'h9d)) : wire794[(4'h9):(4'h9)]))) > (|((&forvar807) ?
                  reg802[(2'h2):(1'h1)] : $signed((8'hbf)))));
            end
          reg821 <= {reg801[(1'h0):(1'h0)]};
          reg822 = reg808[(2'h3):(1'h0)];
          for (forvar823 = (1'h0); (forvar823 < (1'h1)); forvar823 = (forvar823 + (1'h1)))
            begin
              reg824 = $signed($unsigned({($unsigned(wire793) != (~reg808)),
                  wire794}));
            end
          reg825 = (-$signed(reg809));
        end
    end
  assign wire826 = $signed((~&(8'hba)));
  always
    @(posedge clk) begin
      reg827 <= reg822;
      reg828 <= reg814;
    end
  always
    @(posedge clk) begin
      reg829 <= (|$unsigned(reg825[(3'h4):(3'h4)]));
      reg830 <= $unsigned($unsigned(reg815[(3'h4):(2'h2)]));
      reg831 <= (reg799 & $signed((wire805[(3'h4):(1'h1)] >= (7'h42))));
      reg832 <= ($signed(({$unsigned(reg820), (reg799 ? reg828 : reg825)} ?
              ($unsigned((8'ha1)) >>> (wire806 + reg828)) : (((8'hb8) ?
                      reg800 : reg813) ?
                  reg824[(2'h3):(1'h0)] : $unsigned(wire803)))) ?
          $signed((~|forvar810[(2'h2):(1'h0)])) : ($signed((~&wire805)) ?
              $signed((reg820[(4'ha):(3'h6)] ?
                  $unsigned(wire826) : reg799)) : (~$unsigned($signed(wire790)))));
    end
  always
    @(posedge clk) begin
      reg833 <= (~|wire789);
    end
  always
    @(posedge clk) begin
      reg834 = ({(^forvar818),
          $unsigned(($unsigned(wire805) - reg801[(3'h5):(2'h3)]))} & (-reg808));
      reg835 = {(+$unsigned($unsigned((~|wire796)))),
          {(reg813 << $signed(((8'hb5) ? wire797 : reg814))),
              ($unsigned(reg813[(1'h0):(1'h0)]) ?
                  $unsigned(reg825) : wire791)}};
      reg836 <= (&$unsigned((^reg832)));
      reg837 = {(reg799 + $unsigned((~^reg833[(4'h8):(3'h4)]))),
          ((8'ha3) ?
              (reg825[(4'h8):(4'h8)] ?
                  ((reg834 ? forvar811 : forvar823) ?
                      $unsigned(reg829) : $signed(reg799)) : ((forvar818 < wire826) <= reg813)) : (^~(~^wire790)))};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1133  (y, clk, wire1138, wire1137, wire1136, wire1135, wire1134);
  output wire [(32'h4a8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire1138;
  input wire [(5'h12):(1'h0)] wire1137;
  input wire [(4'h9):(1'h0)] wire1136;
  input wire signed [(5'h15):(1'h0)] wire1135;
  input wire signed [(5'h14):(1'h0)] wire1134;
  wire [(2'h2):(1'h0)] wire1687;
  wire signed [(5'h10):(1'h0)] wire1652;
  wire signed [(5'h14):(1'h0)] wire1651;
  wire [(4'he):(1'h0)] wire1650;
  reg signed [(4'h9):(1'h0)] reg1649 = (1'h0);
  reg [(5'h13):(1'h0)] reg1648 = (1'h0);
  reg [(3'h6):(1'h0)] reg1647 = (1'h0);
  reg [(5'h10):(1'h0)] reg1646 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1645;
  reg [(5'h10):(1'h0)] reg1644 = (1'h0);
  reg [(5'h10):(1'h0)] reg1643 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1642 = (1'h0);
  reg [(2'h2):(1'h0)] reg1641 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1640 = (1'h0);
  reg [(4'h8):(1'h0)] reg1639 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1638 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1637 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1636 = (1'h0);
  reg [(5'h11):(1'h0)] reg1635 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1634 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1633 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1632 = (1'h0);
  reg [(3'h5):(1'h0)] reg1631 = (1'h0);
  wire [(4'hc):(1'h0)] wire1629;
  reg signed [(5'h10):(1'h0)] reg1166 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1165 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1164 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1163 = (1'h0);
  reg [(4'h8):(1'h0)] reg1162 = (1'h0);
  reg [(5'h14):(1'h0)] reg1161 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1160 = (1'h0);
  reg [(4'hc):(1'h0)] reg1159 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1158 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1157 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1156 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire1155;
  reg signed [(4'he):(1'h0)] reg1154 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1153 = (1'h0);
  reg [(3'h7):(1'h0)] reg1152 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1151 = (1'h0);
  reg [(4'h8):(1'h0)] reg1150 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1149 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1148 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1147 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1146 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1145 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1144 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1143 = (1'h0);
  reg [(3'h6):(1'h0)] reg1142 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1141 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire1140;
  wire [(5'h10):(1'h0)] wire1139;
  reg signed [(3'h4):(1'h0)] reg1689 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1690 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1691 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1692 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1693 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1694 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1695 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1696 = (1'h0);
  reg [(5'h15):(1'h0)] reg1697 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1698 = (1'h0);
  reg [(4'hc):(1'h0)] reg1699 = (1'h0);
  reg [(3'h5):(1'h0)] reg1700 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1701 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1698 = (1'h0);
  wire [(5'h12):(1'h0)] wire1890;
  wire [(4'hd):(1'h0)] wire1892;
  reg [(5'h11):(1'h0)] reg1893 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1894 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1895 = (1'h0);
  reg [(4'h8):(1'h0)] reg1896 = (1'h0);
  reg [(4'hf):(1'h0)] reg1897 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1898 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1899 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1900 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1901 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1902 = (1'h0);
  reg [(4'he):(1'h0)] reg1903 = (1'h0);
  reg [(5'h11):(1'h0)] reg1904 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1905 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1906 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1907 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1908 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1909 = (1'h0);
  reg [(4'ha):(1'h0)] reg1910 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1911 = (1'h0);
  reg [(4'h9):(1'h0)] reg1912 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1913 = (1'h0);
  reg [(4'ha):(1'h0)] reg1914 = (1'h0);
  reg [(4'ha):(1'h0)] reg1915 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1916 = (1'h0);
  reg [(4'h8):(1'h0)] reg1917 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1918 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire2663;
  assign y = {wire1687,
                 wire1652,
                 wire1651,
                 wire1650,
                 reg1649,
                 reg1648,
                 reg1647,
                 reg1646,
                 wire1645,
                 reg1644,
                 reg1643,
                 reg1642,
                 reg1641,
                 reg1640,
                 reg1639,
                 reg1638,
                 forvar1637,
                 reg1636,
                 reg1635,
                 forvar1634,
                 reg1633,
                 reg1632,
                 reg1631,
                 wire1629,
                 reg1166,
                 reg1165,
                 reg1164,
                 reg1163,
                 reg1162,
                 reg1161,
                 reg1160,
                 reg1159,
                 reg1158,
                 forvar1157,
                 reg1156,
                 wire1155,
                 reg1154,
                 reg1153,
                 reg1152,
                 reg1151,
                 reg1150,
                 forvar1149,
                 reg1148,
                 reg1147,
                 reg1146,
                 reg1145,
                 reg1144,
                 forvar1143,
                 reg1142,
                 reg1141,
                 wire1140,
                 wire1139,
                 reg1689,
                 forvar1690,
                 reg1691,
                 forvar1692,
                 reg1693,
                 reg1694,
                 reg1695,
                 reg1696,
                 reg1697,
                 forvar1698,
                 reg1699,
                 reg1700,
                 reg1701,
                 reg1698,
                 wire1890,
                 wire1892,
                 reg1893,
                 forvar1894,
                 reg1895,
                 reg1896,
                 reg1897,
                 reg1898,
                 reg1899,
                 reg1900,
                 forvar1901,
                 reg1902,
                 reg1903,
                 reg1904,
                 forvar1905,
                 forvar1906,
                 reg1907,
                 forvar1908,
                 reg1909,
                 reg1910,
                 reg1911,
                 reg1912,
                 forvar1913,
                 reg1914,
                 reg1915,
                 reg1916,
                 reg1917,
                 reg1918,
                 wire2663,
                 (1'h0)};
  assign wire1139 = {wire1134[(2'h2):(1'h1)]};
  assign wire1140 = $unsigned((wire1138 < (($signed(wire1134) ?
                            (wire1139 ^ wire1136) : (wire1139 <<< (8'hb6))) ?
                        wire1134[(2'h3):(1'h1)] : (+$unsigned(wire1136)))));
  always
    @(posedge clk) begin
      reg1141 = (((($unsigned(wire1135) * $signed(wire1139)) ?
              (&$unsigned(wire1139)) : $signed({wire1140, wire1140})) ?
          wire1135[(3'h7):(2'h2)] : ((((8'hbd) ?
                  wire1138 : wire1136) ~^ (wire1134 ? wire1139 : wire1134)) ?
              $unsigned({wire1134}) : ((-wire1139) ?
                  $signed((8'hbb)) : wire1135[(3'h6):(3'h4)]))) + {$unsigned($unsigned((~^wire1139)))});
      reg1142 = (^~wire1140[(3'h4):(3'h4)]);
      for (forvar1143 = (1'h0); (forvar1143 < (3'h4)); forvar1143 = (forvar1143 + (1'h1)))
        begin
          reg1144 <= (wire1138[(3'h4):(1'h0)] ?
              ($signed(wire1134[(4'h9):(3'h7)]) > $unsigned(wire1139)) : (-(({(8'h9e)} >>> $signed(wire1140)) ^~ $unsigned($signed(reg1142)))));
          reg1145 <= ((-($unsigned((wire1137 > forvar1143)) ?
                  ((forvar1143 ~^ wire1139) ~^ (wire1135 ?
                      reg1144 : reg1142)) : (wire1136[(2'h2):(1'h1)] <= $signed(wire1134)))) ?
              $unsigned((|$signed(wire1135))) : ((($signed(wire1135) ?
                      $signed(wire1139) : (wire1138 ~^ (8'hbc))) ?
                  $signed($unsigned(wire1139)) : {wire1134}) > wire1137));
          reg1146 <= ($unsigned($unsigned($unsigned((wire1138 ?
              wire1137 : wire1137)))) - (wire1134[(3'h4):(2'h2)] > wire1137));
          reg1147 <= (~|$unsigned(({(wire1140 ? reg1141 : reg1144), wire1140} ?
              $unsigned(reg1142) : $signed($unsigned(wire1138)))));
          reg1148 <= ({reg1145, $signed((|{(8'ha9), reg1145}))} ?
              reg1147[(4'h8):(4'h8)] : ((!wire1135) ?
                  ((forvar1143[(3'h7):(3'h5)] ?
                      (!reg1142) : $signed(wire1138)) & $signed((reg1144 ?
                      wire1140 : reg1146))) : ({{reg1144}, (^wire1134)} ?
                      (+$unsigned(wire1137)) : $signed($unsigned(reg1146)))));
        end
      for (forvar1149 = (1'h0); (forvar1149 < (3'h4)); forvar1149 = (forvar1149 + (1'h1)))
        begin
          reg1150 = wire1138;
          reg1151 <= (($signed(wire1138) ?
              reg1142[(3'h6):(1'h1)] : ($signed({reg1142}) ^~ ($signed(reg1145) == ((8'hbb) <<< (8'h9f))))) + ((wire1134[(4'he):(2'h3)] * (wire1137[(4'he):(3'h6)] | (~|reg1144))) != wire1136[(3'h7):(2'h3)]));
          reg1152 = $signed((^~{(reg1146[(3'h5):(3'h5)] ?
                  {reg1147} : $unsigned(reg1141)),
              ((wire1137 << wire1140) ?
                  (wire1138 ? wire1137 : (8'ha0)) : ((8'ha3) ?
                      forvar1143 : wire1140))}));
          reg1153 = (wire1140[(2'h3):(1'h1)] || reg1142[(3'h6):(1'h0)]);
        end
      reg1154 <= (~^{(reg1151 != (((8'hb9) || (8'hba)) ?
              (wire1138 >>> reg1148) : (reg1145 ~^ reg1153))),
          $signed((~|$unsigned((8'ha6))))});
    end
  assign wire1155 = wire1134[(5'h10):(3'h5)];
  always
    @(posedge clk) begin
      reg1156 = {($signed(((forvar1143 ^~ (7'h40)) ?
                  wire1137[(1'h1):(1'h1)] : {reg1147})) ?
              (~|{(~reg1145), reg1152}) : (8'hb7))};
      for (forvar1157 = (1'h0); (forvar1157 < (1'h1)); forvar1157 = (forvar1157 + (1'h1)))
        begin
          reg1158 <= $unsigned((+$unsigned($unsigned((wire1135 < reg1146)))));
          reg1159 <= (forvar1157 + (^~reg1146));
          reg1160 <= forvar1149;
          reg1161 <= reg1151;
        end
      reg1162 <= $unsigned(((~|$signed($unsigned(reg1158))) ?
          {wire1137} : forvar1157));
    end
  always
    @(posedge clk) begin
      reg1163 = ((~^wire1134) ?
          reg1144[(1'h0):(1'h0)] : ($unsigned(forvar1157) == ({(wire1137 ^ reg1145)} ?
              forvar1149[(4'ha):(4'h9)] : $signed($signed(wire1138)))));
      reg1164 <= $unsigned($unsigned(({(reg1146 != (8'hb7))} ?
          $unsigned((-reg1144)) : wire1137[(3'h7):(2'h3)])));
      reg1165 <= $signed({($unsigned({wire1135}) ?
              reg1141[(3'h7):(2'h2)] : (~$signed(reg1161))),
          $signed((wire1136 >= {forvar1149, (8'hba)}))});
      reg1166 = ((~&(^~reg1160[(3'h7):(2'h3)])) - reg1142);
    end
  module1167 modinst1630 (wire1629, clk, reg1163, reg1147, reg1150, wire1136);
  always
    @(posedge clk) begin
      reg1631 <= ((8'ha4) <= (8'ha4));
      reg1632 <= wire1134;
      reg1633 <= {$unsigned((-(((8'ha2) >>> (8'h9d)) ?
              wire1137[(3'h5):(3'h4)] : (7'h42))))};
    end
  always
    @(posedge clk) begin
      for (forvar1634 = (1'h0); (forvar1634 < (3'h4)); forvar1634 = (forvar1634 + (1'h1)))
        begin
          reg1635 <= ({{{(reg1631 ? reg1159 : reg1164), $signed(wire1629)},
                  $signed((reg1631 ? reg1631 : reg1166))},
              (-(8'h9c))} - ({$unsigned((reg1145 ?
                  wire1138 : forvar1634))} >>> reg1152[(2'h2):(1'h0)]));
          reg1636 = reg1145[(3'h7):(3'h5)];
          for (forvar1637 = (1'h0); (forvar1637 < (2'h3)); forvar1637 = (forvar1637 + (1'h1)))
            begin
              reg1638 <= (|$signed($unsigned(({reg1144,
                  (8'hba)} || $unsigned(reg1161)))));
              reg1639 = (($unsigned((~^(reg1635 & reg1162))) ?
                  {reg1152,
                      $unsigned(reg1151[(4'h8):(2'h3)])} : reg1632[(2'h3):(1'h0)]) - ($unsigned(reg1162) >> $signed($unsigned(wire1139))));
              reg1640 <= wire1138;
              reg1641 = wire1136[(4'h8):(3'h7)];
            end
          reg1642 <= ($signed($signed($unsigned((~&forvar1143)))) <<< wire1155[(4'h9):(3'h5)]);
          reg1643 = $signed(reg1146);
        end
      reg1644 <= (wire1139 ^ (reg1147[(3'h4):(2'h3)] ?
          {reg1642[(3'h4):(1'h1)],
              $unsigned((reg1154 && (8'h9d)))} : $unsigned((~(8'hb1)))));
    end
  assign wire1645 = $signed(reg1639[(4'h8):(3'h5)]);
  always
    @(posedge clk) begin
      reg1646 <= forvar1634[(3'h4):(2'h2)];
      reg1647 = reg1147;
      reg1648 = $unsigned(($signed(($signed(wire1134) || $unsigned(wire1139))) ^ reg1156[(3'h6):(1'h1)]));
      reg1649 = reg1162[(3'h5):(1'h1)];
    end
  assign wire1650 = (reg1638 ? reg1141 : (|$unsigned((~^(reg1632 | (7'h43))))));
  assign wire1651 = $unsigned(((8'hb7) >> (8'hb6)));
  assign wire1652 = (|$unsigned(reg1633));
  module1653 modinst1688 (.wire1656(reg1162), .wire1654(reg1156), .y(wire1687), .wire1658(reg1145), .wire1655(wire1645), .wire1657(reg1633), .clk(clk));
  always
    @(posedge clk) begin
      reg1689 <= $signed({$unsigned(({reg1646, reg1161} ~^ (wire1645 ?
              reg1158 : wire1650)))});
      for (forvar1690 = (1'h0); (forvar1690 < (1'h0)); forvar1690 = (forvar1690 + (1'h1)))
        begin
          reg1691 <= {reg1158[(1'h0):(1'h0)],
              (reg1642[(2'h2):(2'h2)] ?
                  (((8'ha2) ?
                      forvar1149[(4'he):(1'h0)] : (reg1643 <<< wire1629)) ~^ (^~{reg1161,
                      (8'hb5)})) : $unsigned((^~(&reg1642))))};
          for (forvar1692 = (1'h0); (forvar1692 < (1'h0)); forvar1692 = (forvar1692 + (1'h1)))
            begin
              reg1693 = $signed(((-((reg1642 ^~ (8'haf)) > $unsigned(reg1648))) ?
                  (!{wire1140[(1'h1):(1'h0)],
                      {reg1156}}) : $unsigned({(wire1136 == reg1160)})));
              reg1694 = $signed(((8'ha8) ?
                  {($signed(reg1646) & reg1164),
                      ($unsigned(reg1693) * ((8'hac) && wire1140))} : $signed(reg1632[(1'h0):(1'h0)])));
            end
          reg1695 = ($unsigned($unsigned((^~{forvar1149}))) ?
              (8'hae) : $signed((wire1136[(3'h6):(1'h1)] ?
                  ((!(7'h43)) ?
                      $signed(reg1689) : $signed(reg1154)) : $signed((!(8'ha1))))));
          reg1696 = $unsigned(((~|(reg1695 ? $signed(reg1146) : {reg1643})) ?
              (|(reg1146 ? wire1650 : (-reg1644))) : reg1165));
          reg1697 <= ((^(~&(((8'ha0) ? reg1646 : wire1134) ?
                  (reg1145 ? wire1134 : (8'hb8)) : $unsigned(reg1142)))) ?
              reg1695 : ((($unsigned(reg1141) ?
                      $signed(reg1649) : wire1629) ~^ (&(reg1635 != reg1144))) ?
                  (-(^(+reg1640))) : (8'hbb)));
        end
      if ($signed($signed($signed(((wire1650 & wire1137) && {reg1158})))))
        begin
          for (forvar1698 = (1'h0); (forvar1698 < (1'h1)); forvar1698 = (forvar1698 + (1'h1)))
            begin
              reg1699 <= ((((+(&wire1650)) ?
                          ((^wire1629) ?
                              {forvar1637, reg1159} : {wire1137,
                                  reg1159}) : $unsigned($signed(wire1629))) ?
                      {$unsigned(wire1650)} : (reg1158 ?
                          {$signed(reg1643),
                              $signed(forvar1690)} : $unsigned((&(8'hb1))))) ?
                  ($signed($signed((reg1153 ?
                      reg1162 : reg1151))) ^~ reg1643) : $signed(reg1631[(2'h3):(2'h3)]));
              reg1700 <= $signed({reg1146[(3'h7):(3'h7)],
                  $unsigned(wire1135[(4'h9):(3'h4)])});
              reg1701 <= ($unsigned(reg1162[(3'h5):(3'h4)]) && $signed(reg1151[(3'h5):(1'h0)]));
            end
        end
      else
        begin
          reg1698 <= (~^$unsigned(reg1152[(3'h4):(2'h3)]));
          reg1699 = {$signed({($unsigned(reg1643) >= reg1648[(2'h2):(1'h1)]),
                  ($unsigned(wire1136) ? reg1147 : $unsigned(reg1144))}),
              reg1696[(3'h5):(3'h5)]};
        end
    end
  module1702 modinst1891 (.wire1706(reg1648), .y(wire1890), .wire1704(wire1138), .wire1703(wire1652), .clk(clk), .wire1705(reg1154));
  assign wire1892 = (reg1147 ?
                        $unsigned($signed(((wire1140 ?
                            (8'hb8) : reg1696) >> $unsigned(forvar1690)))) : (~^((wire1890[(5'h10):(5'h10)] > $signed((8'hae))) ?
                            $unsigned((8'hac)) : reg1640[(4'h8):(2'h2)])));
  always
    @(posedge clk) begin
      reg1893 = (~^wire1890[(1'h0):(1'h0)]);
      for (forvar1894 = (1'h0); (forvar1894 < (2'h2)); forvar1894 = (forvar1894 + (1'h1)))
        begin
          reg1895 <= (+(|{(-$signed(wire1651)),
              $unsigned(wire1651[(4'hc):(4'h8)])}));
          reg1896 <= $unsigned(forvar1157);
          reg1897 = ((reg1895[(5'h11):(1'h0)] || (8'hbb)) ?
              {$signed(($unsigned(reg1166) ?
                      (!reg1642) : wire1650[(3'h6):(1'h1)]))} : (reg1640 + $unsigned((forvar1149 ^~ (8'hb9)))));
          reg1898 = reg1701[(1'h1):(1'h1)];
        end
    end
  always
    @(posedge clk) begin
      reg1899 <= $unsigned(reg1145[(2'h2):(2'h2)]);
      reg1900 <= {($unsigned(reg1693) == (wire1892 ?
              (wire1134 && $unsigned((8'hbf))) : (8'h9e))),
          ({$signed((reg1631 > reg1635))} ?
              (((wire1645 << reg1145) < $signed((8'hac))) ?
                  $unsigned((reg1631 <<< forvar1698)) : (~|$signed(reg1160))) : $unsigned($signed($unsigned(reg1166))))};
      for (forvar1901 = (1'h0); (forvar1901 < (3'h4)); forvar1901 = (forvar1901 + (1'h1)))
        begin
          reg1902 = (reg1161 - wire1651);
          reg1903 <= (reg1147 && (^~((8'ha1) ?
              reg1145[(5'h12):(3'h6)] : (|(reg1164 & (7'h41))))));
          reg1904 <= reg1903;
        end
      for (forvar1905 = (1'h0); (forvar1905 < (1'h1)); forvar1905 = (forvar1905 + (1'h1)))
        begin
          for (forvar1906 = (1'h0); (forvar1906 < (1'h1)); forvar1906 = (forvar1906 + (1'h1)))
            begin
              reg1907 = $unsigned($unsigned($unsigned((~reg1147[(5'h12):(4'h9)]))));
            end
          for (forvar1908 = (1'h0); (forvar1908 < (3'h4)); forvar1908 = (forvar1908 + (1'h1)))
            begin
              reg1909 <= $unsigned(reg1154);
              reg1910 <= forvar1698;
            end
          reg1911 = {$signed((8'hbf)), reg1647};
          reg1912 <= $unsigned($signed(wire1138));
          for (forvar1913 = (1'h0); (forvar1913 < (2'h2)); forvar1913 = (forvar1913 + (1'h1)))
            begin
              reg1914 <= (^~{$signed(($unsigned(reg1701) ?
                      wire1138 : $signed(wire1155))),
                  (|((reg1693 ? reg1158 : (8'h9e)) ?
                      (forvar1908 < (8'hb9)) : {wire1155}))});
              reg1915 = reg1144[(1'h1):(1'h0)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg1916 <= (~^(((8'h9c) ?
          $signed((reg1699 ?
              reg1909 : reg1159)) : $unsigned(reg1695[(2'h2):(1'h1)])) - reg1640[(1'h1):(1'h1)]));
      reg1917 <= ((reg1151[(2'h3):(2'h2)] <<< (reg1693[(2'h3):(2'h2)] ?
              $signed($unsigned((8'hb3))) : (reg1697[(1'h0):(1'h0)] | (reg1648 && forvar1637)))) ?
          reg1910[(3'h4):(2'h2)] : wire1652[(4'hb):(2'h3)]);
      reg1918 <= reg1898;
    end
  module1919 modinst2664 (wire2663, clk, reg1896, reg1147, wire1134, reg1911, wire1651);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module906
#( parameter param1111 = {(&(!((~&(8'hb1)) * ((8'ha2) == (8'ha3))))), {((((7'h44) - (8'hbe)) >>> ((8'h9d) >>> (8'haa))) ? (8'ha3) : (((8'ha6) > (8'hb4)) + ((8'hbf) ? (8'haf) : (8'hb5)))), ({((8'ha4) ? (8'hbc) : (7'h44))} ? (~((8'hb6) ^~ (8'hbe))) : ((8'ha3) * (-(7'h41))))}} )
(y, clk, wire910, wire909, wire908, wire907);
  output wire [(32'h18b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire910;
  input wire [(2'h3):(1'h0)] wire909;
  input wire [(5'h13):(1'h0)] wire908;
  input wire [(4'hf):(1'h0)] wire907;
  wire signed [(3'h6):(1'h0)] wire1110;
  wire [(4'hc):(1'h0)] wire1109;
  reg signed [(5'h12):(1'h0)] reg1108 = (1'h0);
  reg [(4'hc):(1'h0)] reg1107 = (1'h0);
  reg [(3'h5):(1'h0)] reg1106 = (1'h0);
  reg [(2'h2):(1'h0)] reg1105 = (1'h0);
  reg [(5'h14):(1'h0)] reg1104 = (1'h0);
  reg [(4'hb):(1'h0)] reg1103 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1102 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1101 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire1100;
  reg [(5'h14):(1'h0)] reg1099 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1098 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1097 = (1'h0);
  wire [(2'h2):(1'h0)] wire1095;
  wire [(4'hd):(1'h0)] wire964;
  reg signed [(3'h6):(1'h0)] reg963 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg962 = (1'h0);
  reg [(4'he):(1'h0)] reg961 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar960 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire958;
  reg [(4'ha):(1'h0)] reg924 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg923 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg922 = (1'h0);
  wire [(2'h2):(1'h0)] wire921;
  wire signed [(5'h14):(1'h0)] wire920;
  reg [(5'h12):(1'h0)] reg919 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg918 = (1'h0);
  wire [(4'h9):(1'h0)] wire917;
  reg signed [(5'h10):(1'h0)] reg916 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg915 = (1'h0);
  reg [(4'hc):(1'h0)] reg914 = (1'h0);
  reg [(4'hc):(1'h0)] reg913 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg912 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar911 = (1'h0);
  assign y = {wire1110,
                 wire1109,
                 reg1108,
                 reg1107,
                 reg1106,
                 reg1105,
                 reg1104,
                 reg1103,
                 reg1102,
                 reg1101,
                 wire1100,
                 reg1099,
                 reg1098,
                 reg1097,
                 wire1095,
                 wire964,
                 reg963,
                 reg962,
                 reg961,
                 forvar960,
                 wire958,
                 reg924,
                 reg923,
                 reg922,
                 wire921,
                 wire920,
                 reg919,
                 reg918,
                 wire917,
                 reg916,
                 reg915,
                 reg914,
                 reg913,
                 reg912,
                 forvar911,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar911 = (1'h0); (forvar911 < (3'h4)); forvar911 = (forvar911 + (1'h1)))
        begin
          reg912 <= wire908[(5'h10):(4'hb)];
          reg913 <= $signed(reg912);
        end
      reg914 <= forvar911;
      reg915 <= (~^$signed((wire907[(4'hb):(4'h8)] | ((reg914 | wire907) & (-reg913)))));
      reg916 <= wire909;
    end
  assign wire917 = $unsigned((+(({wire910} > (forvar911 ^~ wire907)) ?
                       (8'hac) : $unsigned($unsigned((7'h43))))));
  always
    @(posedge clk) begin
      reg918 = wire909;
      reg919 <= (^~$unsigned(wire909[(2'h2):(1'h0)]));
    end
  assign wire920 = ($signed(reg916) ?
                       ((((~&(8'hbb)) >>> wire908) >= (((8'hb2) ?
                           wire917 : (8'ha0)) ~^ (wire910 >= forvar911))) | $signed($signed($unsigned(wire917)))) : (8'hab));
  assign wire921 = wire907;
  always
    @(posedge clk) begin
      reg922 = $unsigned($signed({forvar911}));
      reg923 <= (((-{((8'hb2) ? reg912 : wire920),
              (wire920 <<< wire920)}) + $unsigned((^(wire908 < wire921)))) ?
          ((!($unsigned((8'h9e)) ? (wire920 ? reg915 : forvar911) : reg916)) ?
              reg914 : {((!wire910) ?
                      $signed(reg913) : wire909[(1'h0):(1'h0)])}) : reg914[(2'h3):(2'h2)]);
      reg924 <= ($unsigned($unsigned((reg915[(3'h4):(1'h0)] ?
          $unsigned(wire908) : $signed((8'ha4))))) + ($signed(wire907) << ((~^(wire910 ?
              reg918 : reg922)) ?
          ((wire908 ? reg913 : wire908) ?
              (~|reg915) : (7'h42)) : wire920[(1'h1):(1'h1)])));
    end
  module925 modinst959 (wire958, clk, wire908, reg913, reg924, wire920);
  always
    @(posedge clk) begin
      for (forvar960 = (1'h0); (forvar960 < (2'h3)); forvar960 = (forvar960 + (1'h1)))
        begin
          reg961 <= (!wire917);
        end
      reg962 <= reg913;
      reg963 <= {wire910[(1'h1):(1'h0)], $unsigned((&reg923[(1'h1):(1'h1)]))};
    end
  assign wire964 = {reg924, wire908[(3'h4):(2'h3)]};
  module965 modinst1096 (wire1095, clk, reg912, reg919, wire910, reg922);
  always
    @(posedge clk) begin
      reg1097 <= ((~^(~^$signed((^(8'hb4))))) || (^~$unsigned((^~(-reg916)))));
      reg1098 <= $signed((~&$signed((|(forvar911 >= reg923)))));
      reg1099 <= (($signed(($signed(reg922) ^ reg918[(4'hd):(2'h3)])) ?
              (^~wire917) : reg963[(3'h4):(1'h1)]) ?
          ($signed($signed((+reg913))) ?
              ($signed(forvar911) ?
                  ({wire920} ?
                      $signed(reg922) : wire920[(3'h6):(1'h0)]) : ({wire907,
                          reg924} ?
                      wire1095 : $unsigned((8'hb2)))) : reg922) : (($unsigned((reg918 ?
                  reg918 : wire964)) ?
              {reg923, {wire1095, reg963}} : (wire909[(1'h1):(1'h1)] ?
                  $signed(wire917) : $unsigned(forvar960))) != ($signed($unsigned(reg1097)) == {((8'hb5) ?
                  wire910 : reg922)})));
    end
  assign wire1100 = ($signed((8'hb3)) ? {reg916[(4'hd):(4'hb)]} : reg1099);
  always
    @(posedge clk) begin
      reg1101 = (!(8'ha5));
      reg1102 <= ((8'hbd) >>> reg961);
      reg1103 = ($unsigned(wire907[(3'h7):(3'h4)]) * (~|({(&reg919)} & (reg1102[(1'h0):(1'h0)] ?
          $signed(forvar960) : reg1102))));
      reg1104 = wire920;
      reg1105 = ((~reg961[(1'h1):(1'h0)]) > wire921);
    end
  always
    @(posedge clk) begin
      reg1106 <= forvar911[(1'h0):(1'h0)];
      reg1107 <= $unsigned($signed((({reg924} ^ (~reg918)) <= $unsigned($unsigned(wire909)))));
      reg1108 <= reg912[(5'h12):(3'h5)];
    end
  assign wire1109 = reg1097;
  assign wire1110 = $unsigned((reg913 ? reg1107[(3'h6):(1'h1)] : reg916));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module965
#( parameter param1093 = (((~{((8'h9e) ? (8'hbe) : (8'ha6)), ((8'ha4) | (8'hb6))}) ? (~|(((8'hb0) >> (8'hbc)) | (~&(8'ha5)))) : (~&((~|(8'hbb)) || ((8'ha2) ? (7'h43) : (8'hbd))))) ~^ ((((+(8'hbd)) + (8'hb6)) ? (((7'h44) ? (7'h44) : (8'ha1)) * {(8'hb2)}) : (^((8'haa) ? (8'hab) : (7'h42)))) ? (^~({(8'hb0)} >>> {(7'h42)})) : ((^~((8'hbf) ? (8'ha4) : (8'hb9))) >>> ({(8'hbf)} ? ((8'hac) > (8'hb9)) : (~(8'hb4))))))
, parameter param1094 = (~|{((7'h40) != {(!param1093)}), ((~|(!param1093)) << param1093)}) )
(y, clk, wire969, wire968, wire967, wire966);
  output wire [(32'h30a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire969;
  input wire [(5'h12):(1'h0)] wire968;
  input wire signed [(3'h6):(1'h0)] wire967;
  input wire [(3'h6):(1'h0)] wire966;
  reg signed [(3'h5):(1'h0)] reg1092 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1091 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1090 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1089 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1088 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1087 = (1'h0);
  reg [(5'h11):(1'h0)] reg1086 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1085 = (1'h0);
  reg [(4'hc):(1'h0)] reg1084 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1083 = (1'h0);
  reg [(2'h3):(1'h0)] reg1082 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1081 = (1'h0);
  reg [(3'h4):(1'h0)] reg1080 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1079;
  reg [(4'hf):(1'h0)] reg1078 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire1076;
  wire signed [(4'hc):(1'h0)] wire1019;
  wire signed [(4'hf):(1'h0)] wire1018;
  wire signed [(5'h10):(1'h0)] wire1017;
  wire signed [(4'he):(1'h0)] wire1016;
  reg signed [(5'h10):(1'h0)] reg1015 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1014 = (1'h0);
  reg [(4'he):(1'h0)] forvar1013 = (1'h0);
  reg [(2'h3):(1'h0)] reg1012 = (1'h0);
  reg [(2'h3):(1'h0)] reg1011 = (1'h0);
  reg [(4'ha):(1'h0)] reg1010 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1009 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1008 = (1'h0);
  reg [(4'hb):(1'h0)] reg1007 = (1'h0);
  reg [(4'hf):(1'h0)] reg1006 = (1'h0);
  reg [(5'h12):(1'h0)] reg1005 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1004 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire1003;
  reg signed [(4'hb):(1'h0)] reg1002 = (1'h0);
  reg [(3'h7):(1'h0)] reg1001 = (1'h0);
  reg [(3'h4):(1'h0)] reg1000 = (1'h0);
  reg [(5'h15):(1'h0)] reg999 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg998 = (1'h0);
  reg [(4'ha):(1'h0)] forvar997 = (1'h0);
  reg [(4'he):(1'h0)] reg996 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg995 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar994 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg993 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg992 = (1'h0);
  wire [(5'h13):(1'h0)] wire991;
  wire [(4'hb):(1'h0)] wire990;
  reg [(2'h2):(1'h0)] reg989 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg988 = (1'h0);
  reg [(5'h10):(1'h0)] reg987 = (1'h0);
  reg signed [(4'he):(1'h0)] reg986 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg985 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg984 = (1'h0);
  reg [(4'he):(1'h0)] reg983 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar982 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg981 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg980 = (1'h0);
  reg [(3'h4):(1'h0)] forvar979 = (1'h0);
  reg [(4'h9):(1'h0)] reg978 = (1'h0);
  reg [(5'h15):(1'h0)] reg977 = (1'h0);
  reg [(4'hc):(1'h0)] reg976 = (1'h0);
  reg [(3'h6):(1'h0)] reg975 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar974 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg973 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg972 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg971 = (1'h0);
  reg [(4'hb):(1'h0)] forvar970 = (1'h0);
  assign y = {reg1092,
                 reg1091,
                 reg1090,
                 reg1089,
                 forvar1088,
                 reg1087,
                 reg1086,
                 reg1085,
                 reg1084,
                 forvar1083,
                 reg1082,
                 forvar1081,
                 reg1080,
                 wire1079,
                 reg1078,
                 wire1076,
                 wire1019,
                 wire1018,
                 wire1017,
                 wire1016,
                 reg1015,
                 reg1014,
                 forvar1013,
                 reg1012,
                 reg1011,
                 reg1010,
                 forvar1009,
                 forvar1008,
                 reg1007,
                 reg1006,
                 reg1005,
                 reg1004,
                 wire1003,
                 reg1002,
                 reg1001,
                 reg1000,
                 reg999,
                 reg998,
                 forvar997,
                 reg996,
                 reg995,
                 forvar994,
                 reg993,
                 reg992,
                 wire991,
                 wire990,
                 reg989,
                 reg988,
                 reg987,
                 reg986,
                 reg985,
                 reg984,
                 reg983,
                 forvar982,
                 reg981,
                 reg980,
                 forvar979,
                 reg978,
                 reg977,
                 reg976,
                 reg975,
                 forvar974,
                 reg973,
                 reg972,
                 reg971,
                 forvar970,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar970 = (1'h0); (forvar970 < (1'h1)); forvar970 = (forvar970 + (1'h1)))
        begin
          reg971 <= (^~$unsigned($unsigned((&$signed((8'hbb))))));
          reg972 <= {(((^(wire966 * (8'hb0))) <<< ((|reg971) ?
                      $signed(wire966) : {wire966, wire968})) ?
                  ($signed(((8'h9f) + wire968)) >= ({wire966, wire969} ?
                      wire969 : wire968)) : (wire967 ?
                      $unsigned(reg971[(2'h2):(1'h1)]) : $signed((wire969 ?
                          wire969 : (8'ha5))))),
              (forvar970 ?
                  (+$unsigned((forvar970 + wire968))) : $unsigned(reg971))};
          reg973 <= $signed($unsigned(wire968[(4'h8):(1'h0)]));
          for (forvar974 = (1'h0); (forvar974 < (2'h3)); forvar974 = (forvar974 + (1'h1)))
            begin
              reg975 <= {reg971,
                  ((($signed(forvar970) || $unsigned(reg971)) ?
                      ((forvar974 >> wire967) ?
                          (wire969 ? (8'hbc) : reg973) : (reg971 ?
                              reg973 : forvar970)) : $unsigned((wire967 ?
                          forvar970 : wire969))) << $unsigned($signed(((8'hac) >>> wire966))))};
              reg976 <= (8'h9d);
              reg977 = $signed((-({(wire969 ? wire969 : reg975),
                  (reg972 ? forvar970 : wire969)} & wire969)));
            end
        end
      reg978 <= $signed((($unsigned(reg971) < {(reg971 ? (8'hbb) : forvar974),
              wire969}) ?
          (wire969[(2'h3):(2'h2)] ^ reg971) : (($unsigned(forvar974) ?
              $unsigned(wire967) : {wire968,
                  (8'h9c)}) >>> (~|$unsigned((8'ha3))))));
      for (forvar979 = (1'h0); (forvar979 < (3'h4)); forvar979 = (forvar979 + (1'h1)))
        begin
          reg980 <= reg975[(2'h3):(1'h1)];
          reg981 <= (8'h9c);
          for (forvar982 = (1'h0); (forvar982 < (2'h3)); forvar982 = (forvar982 + (1'h1)))
            begin
              reg983 <= wire968;
              reg984 <= wire969;
              reg985 <= (wire969[(4'hf):(4'hb)] | $unsigned($signed((+(reg978 ?
                  reg972 : (8'hb1))))));
              reg986 <= $signed(reg978);
            end
          reg987 <= (8'ha9);
        end
      reg988 <= $unsigned($unsigned(forvar970[(4'ha):(2'h3)]));
      reg989 <= (8'hb9);
    end
  assign wire990 = reg971;
  assign wire991 = reg988[(3'h4):(1'h1)];
  always
    @(posedge clk) begin
      reg992 = (((8'hbd) >= reg988[(2'h2):(2'h2)]) & (wire991 - $unsigned($signed(forvar979))));
      reg993 <= reg988[(1'h1):(1'h1)];
      for (forvar994 = (1'h0); (forvar994 < (1'h1)); forvar994 = (forvar994 + (1'h1)))
        begin
          reg995 = reg987[(1'h1):(1'h0)];
          reg996 = {((+reg971[(1'h0):(1'h0)]) ?
                  ($unsigned($signed((8'had))) <<< (^~{forvar982})) : $signed((8'hb9))),
              $unsigned({$signed($unsigned(reg976)), (~&$signed(reg987))})};
          for (forvar997 = (1'h0); (forvar997 < (1'h1)); forvar997 = (forvar997 + (1'h1)))
            begin
              reg998 = reg985[(5'h11):(4'ha)];
              reg999 <= reg983[(4'hb):(3'h4)];
              reg1000 <= $signed(forvar982[(3'h5):(1'h0)]);
            end
          reg1001 <= wire969;
        end
      reg1002 <= $unsigned(reg984);
    end
  assign wire1003 = {(({$signed(reg985), $unsigned(reg976)} ?
                            $signed((~|reg975)) : reg978[(1'h1):(1'h0)]) ^~ reg986),
                        {reg1002[(1'h0):(1'h0)],
                            $signed(forvar994[(4'h8):(2'h3)])}};
  always
    @(posedge clk) begin
      reg1004 <= (&(~^($unsigned(reg984[(5'h13):(2'h2)]) ?
          $signed($signed((8'ha8))) : reg1001)));
      reg1005 <= ($unsigned($unsigned((&reg971))) < {($signed(reg996) ?
              {((8'hb0) >> reg983)} : $unsigned($unsigned(reg984))),
          $unsigned($unsigned($signed((8'hb1))))});
      reg1006 <= $unsigned((reg985[(3'h4):(2'h2)] ?
          $signed((~^{forvar982})) : reg978));
      reg1007 <= wire991[(5'h10):(5'h10)];
      for (forvar1008 = (1'h0); (forvar1008 < (1'h1)); forvar1008 = (forvar1008 + (1'h1)))
        begin
          for (forvar1009 = (1'h0); (forvar1009 < (3'h4)); forvar1009 = (forvar1009 + (1'h1)))
            begin
              reg1010 <= ((-(($unsigned(forvar1009) | wire966[(1'h0):(1'h0)]) ^ wire1003)) << {{reg981[(2'h3):(2'h2)],
                      ((reg973 || reg1002) ?
                          ((8'ha0) <<< reg1000) : (reg973 ^ reg1000))},
                  reg986[(3'h5):(3'h4)]});
            end
          reg1011 <= (&{((|(|reg975)) >>> reg976[(3'h4):(2'h2)]),
              $unsigned((&(reg1004 ? reg1007 : forvar979)))});
          reg1012 = (((8'hb9) ?
              wire991 : $unsigned(((^~reg1005) ?
                  $unsigned(wire967) : (forvar982 ?
                      (8'hae) : reg988)))) ^ ((($unsigned((8'hb5)) ?
              wire969[(3'h6):(2'h3)] : (reg1006 >= reg1006)) ^~ ($unsigned(reg993) ?
              (~reg986) : forvar994)) <= $signed($unsigned(reg1002))));
          for (forvar1013 = (1'h0); (forvar1013 < (3'h4)); forvar1013 = (forvar1013 + (1'h1)))
            begin
              reg1014 <= (forvar982 <= (&$signed($unsigned(reg999))));
            end
          reg1015 <= (^((!($signed(reg972) != (reg985 < (8'hbf)))) ?
              $unsigned((reg984 ?
                  $unsigned((8'hae)) : $signed(reg980))) : $unsigned((8'hbc))));
        end
    end
  assign wire1016 = reg973;
  assign wire1017 = ((~&(($unsigned((7'h42)) ?
                                reg975[(2'h2):(1'h0)] : (reg1015 ?
                                    reg978 : forvar970)) ?
                            $signed(forvar997[(3'h7):(2'h3)]) : ({reg976} ?
                                {(8'hbe), wire991} : {(8'ha4)}))) ?
                        (reg981[(4'h9):(4'h9)] ?
                            (-(|(|reg1014))) : ((wire969 ?
                                (!wire968) : (reg989 ^~ reg995)) < reg1010[(4'h8):(3'h5)])) : wire990[(1'h1):(1'h1)]);
  assign wire1018 = reg971[(1'h0):(1'h0)];
  assign wire1019 = $unsigned((~reg1010));
  module1020 modinst1077 (wire1076, clk, reg975, reg999, reg998, reg995);
  always
    @(posedge clk) begin
      reg1078 = wire1016;
    end
  assign wire1079 = {forvar979[(1'h1):(1'h1)], reg985[(4'h8):(3'h6)]};
  always
    @(posedge clk) begin
      reg1080 <= wire990[(4'hb):(3'h6)];
      for (forvar1081 = (1'h0); (forvar1081 < (2'h2)); forvar1081 = (forvar1081 + (1'h1)))
        begin
          reg1082 <= $unsigned(((~&forvar1081) | reg1011));
          for (forvar1083 = (1'h0); (forvar1083 < (2'h2)); forvar1083 = (forvar1083 + (1'h1)))
            begin
              reg1084 <= $unsigned($unsigned(forvar979));
              reg1085 = ((~|((+reg986) & wire1003)) >> $unsigned((((wire1003 ?
                      reg987 : reg989) <= (reg987 ? reg971 : reg975)) ?
                  reg983[(3'h6):(2'h3)] : {((8'hb5) ? reg971 : reg993)})));
              reg1086 <= reg986;
            end
          reg1087 <= (reg1002[(2'h2):(1'h0)] << (~|reg1004));
          for (forvar1088 = (1'h0); (forvar1088 < (2'h3)); forvar1088 = (forvar1088 + (1'h1)))
            begin
              reg1089 <= ({reg1014[(3'h5):(1'h0)],
                      $signed((wire1076[(4'hf):(1'h1)] < reg978))} ?
                  reg1078 : {((wire968 & $unsigned(reg972)) ?
                          ({reg1014} > $signed(forvar979)) : $unsigned((&reg1085))),
                      $signed(((reg1012 ? wire1019 : forvar970) ?
                          $signed(forvar1083) : (reg984 ?
                              reg1015 : reg1012)))});
            end
        end
      reg1090 <= (~|($unsigned(reg976[(4'hc):(3'h5)]) && reg1087));
      reg1091 <= ($unsigned($unsigned($signed(reg1078[(1'h1):(1'h1)]))) ^ $signed($unsigned((&(8'hbd)))));
    end
  always
    @(posedge clk) begin
      reg1092 <= $signed(wire991[(3'h4):(3'h4)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module925  (y, clk, wire929, wire928, wire927, wire926);
  output wire [(32'h16d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire929;
  input wire [(2'h2):(1'h0)] wire928;
  input wire signed [(4'ha):(1'h0)] wire927;
  input wire [(5'h14):(1'h0)] wire926;
  reg signed [(4'he):(1'h0)] reg957 = (1'h0);
  reg [(3'h5):(1'h0)] reg956 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg955 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg954 = (1'h0);
  reg [(2'h3):(1'h0)] reg953 = (1'h0);
  reg [(3'h4):(1'h0)] reg952 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg951 = (1'h0);
  reg [(5'h13):(1'h0)] forvar950 = (1'h0);
  reg [(5'h10):(1'h0)] reg949 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg948 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg947 = (1'h0);
  reg [(5'h15):(1'h0)] reg946 = (1'h0);
  reg [(5'h13):(1'h0)] forvar945 = (1'h0);
  reg [(3'h6):(1'h0)] reg944 = (1'h0);
  reg [(5'h15):(1'h0)] forvar943 = (1'h0);
  reg [(4'ha):(1'h0)] reg942 = (1'h0);
  reg [(4'hb):(1'h0)] reg941 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg940 = (1'h0);
  reg [(4'hf):(1'h0)] reg939 = (1'h0);
  reg [(4'hc):(1'h0)] reg938 = (1'h0);
  wire [(2'h3):(1'h0)] wire937;
  wire [(4'hb):(1'h0)] wire936;
  reg [(5'h13):(1'h0)] reg935 = (1'h0);
  reg [(4'hf):(1'h0)] reg934 = (1'h0);
  reg [(5'h15):(1'h0)] reg933 = (1'h0);
  wire [(4'h8):(1'h0)] wire932;
  wire signed [(5'h11):(1'h0)] wire931;
  wire [(5'h13):(1'h0)] wire930;
  assign y = {reg957,
                 reg956,
                 reg955,
                 reg954,
                 reg953,
                 reg952,
                 reg951,
                 forvar950,
                 reg949,
                 reg948,
                 reg947,
                 reg946,
                 forvar945,
                 reg944,
                 forvar943,
                 reg942,
                 reg941,
                 reg940,
                 reg939,
                 reg938,
                 wire937,
                 wire936,
                 reg935,
                 reg934,
                 reg933,
                 wire932,
                 wire931,
                 wire930,
                 (1'h0)};
  assign wire930 = (($signed({(wire929 ? wire926 : wire929),
                               $signed(wire929)}) ?
                           wire927 : wire926) ?
                       (((~|(wire928 >>> wire927)) ?
                           wire927 : (((8'hae) <= wire927) ^ $unsigned(wire927))) * (wire928 * wire926)) : ((wire927[(2'h2):(1'h0)] >>> wire927[(1'h1):(1'h1)]) && wire927));
  assign wire931 = $signed($signed({wire929[(2'h2):(1'h1)],
                       ((^~wire929) ?
                           wire929[(3'h6):(1'h1)] : $signed((8'h9c)))}));
  assign wire932 = $unsigned(((8'h9d) ?
                       $signed(((8'haf) > $signed(wire928))) : (wire930[(2'h3):(2'h2)] <= wire927[(3'h4):(3'h4)])));
  always
    @(posedge clk) begin
      reg933 <= ({((((8'ha7) ? wire932 : wire931) ?
                  (~wire931) : wire929) ~^ $unsigned((wire931 | wire932))),
              $unsigned(wire928[(1'h1):(1'h1)])} ?
          ((wire931[(1'h1):(1'h1)] ? wire930 : wire932[(3'h7):(2'h2)]) ?
              $signed((^~$unsigned(wire927))) : (8'hae)) : $signed($signed(wire929[(2'h2):(1'h0)])));
    end
  always
    @(posedge clk) begin
      reg934 <= wire927[(1'h1):(1'h1)];
    end
  always
    @(posedge clk) begin
      reg935 <= {wire931,
          ({wire927[(2'h2):(1'h0)], wire927[(4'h8):(2'h2)]} ?
              $unsigned((wire930 >>> (^wire930))) : $signed($signed((reg934 >= wire930))))};
    end
  assign wire936 = $signed((({wire930} ?
                           $unsigned($signed(wire931)) : (+reg934)) ?
                       wire931[(2'h2):(1'h0)] : (($unsigned(wire926) ?
                               (|reg934) : (-wire927)) ?
                           $signed((~&wire929)) : (^~(^~(8'hbb))))));
  assign wire937 = (+(8'hae));
  always
    @(posedge clk) begin
      reg938 = $unsigned((~^wire926[(4'hb):(3'h6)]));
      reg939 <= wire926;
      reg940 <= wire936[(4'h8):(4'h8)];
    end
  always
    @(posedge clk) begin
      reg941 = reg938;
      reg942 = reg941;
      for (forvar943 = (1'h0); (forvar943 < (1'h0)); forvar943 = (forvar943 + (1'h1)))
        begin
          reg944 = (((reg942[(4'h9):(3'h4)] ^ $signed(wire928[(1'h0):(1'h0)])) & {(~{reg940}),
              ((reg935 ? (8'ha8) : reg942) ?
                  reg934 : wire930)}) || ($signed(reg942) >> (~|{$unsigned(wire928),
              reg935[(5'h13):(1'h1)]})));
          for (forvar945 = (1'h0); (forvar945 < (2'h3)); forvar945 = (forvar945 + (1'h1)))
            begin
              reg946 <= $signed($signed((-((~^reg934) * wire929))));
              reg947 <= ($signed(wire926) + reg938[(2'h2):(1'h1)]);
              reg948 <= ($signed($unsigned((reg947[(1'h1):(1'h0)] >> forvar943))) <<< ($signed($unsigned({wire936,
                      reg938})) ?
                  (reg941 ? $signed((~&reg939)) : wire926) : (8'hae)));
            end
          reg949 <= reg946;
          for (forvar950 = (1'h0); (forvar950 < (2'h3)); forvar950 = (forvar950 + (1'h1)))
            begin
              reg951 <= $unsigned(((|wire927) - $unsigned((~|{reg940,
                  forvar945}))));
              reg952 <= ((((^~{reg948}) ?
                  reg933 : ($unsigned(reg934) ?
                      (^reg951) : (wire937 ~^ forvar945))) == ($signed({reg944}) ?
                  $unsigned((~|reg946)) : $signed((reg938 < forvar943)))) ^ ($signed({reg934[(2'h3):(2'h3)]}) ?
                  {(|(reg934 ? (8'hbb) : reg934)), (+reg951)} : wire928));
              reg953 <= forvar950[(5'h10):(3'h6)];
              reg954 <= forvar950;
              reg955 <= $unsigned($unsigned((~(^~{reg941, wire928}))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg956 = ({(((^~reg944) ?
                  {wire927, reg942} : (wire929 ? forvar950 : (8'hb0))) ?
              $signed($unsigned(reg949)) : ($signed(wire926) ?
                  $unsigned((8'hb2)) : (^~reg947))),
          $signed($signed((&wire928)))} > forvar945);
      reg957 <= (^~reg941);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1020  (y, clk, wire1024, wire1023, wire1022, wire1021);
  output wire [(32'h139):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire1024;
  input wire signed [(4'he):(1'h0)] wire1023;
  input wire [(3'h5):(1'h0)] wire1022;
  input wire signed [(5'h13):(1'h0)] wire1021;
  wire [(4'hf):(1'h0)] wire1075;
  reg [(3'h5):(1'h0)] reg1074 = (1'h0);
  reg [(4'he):(1'h0)] reg1073 = (1'h0);
  reg [(4'hf):(1'h0)] reg1072 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1071 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1070 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1069 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1068 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1067 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1066 = (1'h0);
  reg [(3'h4):(1'h0)] reg1065 = (1'h0);
  reg [(5'h15):(1'h0)] reg1064 = (1'h0);
  reg [(2'h2):(1'h0)] reg1063 = (1'h0);
  reg [(4'hb):(1'h0)] reg1062 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1061 = (1'h0);
  wire [(5'h13):(1'h0)] wire1060;
  wire signed [(5'h13):(1'h0)] wire1058;
  wire [(4'h8):(1'h0)] wire1033;
  reg [(3'h4):(1'h0)] reg1032 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1031 = (1'h0);
  reg [(4'hd):(1'h0)] reg1030 = (1'h0);
  reg [(5'h12):(1'h0)] reg1029 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1028 = (1'h0);
  reg [(5'h11):(1'h0)] reg1027 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1026 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1025 = (1'h0);
  assign y = {wire1075,
                 reg1074,
                 reg1073,
                 reg1072,
                 reg1071,
                 reg1070,
                 reg1069,
                 reg1068,
                 forvar1067,
                 forvar1066,
                 reg1065,
                 reg1064,
                 reg1063,
                 reg1062,
                 forvar1061,
                 wire1060,
                 wire1058,
                 wire1033,
                 reg1032,
                 reg1031,
                 reg1030,
                 reg1029,
                 reg1028,
                 reg1027,
                 forvar1026,
                 reg1025,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1025 <= {(8'ha7), $signed($unsigned({wire1022[(1'h0):(1'h0)]}))};
      for (forvar1026 = (1'h0); (forvar1026 < (1'h1)); forvar1026 = (forvar1026 + (1'h1)))
        begin
          reg1027 = forvar1026[(3'h7):(2'h3)];
          reg1028 <= ((8'h9f) ?
              $signed(($unsigned(wire1021[(1'h0):(1'h0)]) & ({wire1023} - wire1021[(3'h6):(3'h6)]))) : (forvar1026 || $signed($signed(forvar1026[(1'h1):(1'h1)]))));
          reg1029 = $unsigned($unsigned({$signed($unsigned(reg1027))}));
          reg1030 <= $signed($unsigned($unsigned((reg1025[(5'h10):(2'h3)] + {reg1029,
              reg1027}))));
        end
      reg1031 <= $signed(reg1028[(2'h3):(2'h2)]);
      reg1032 = (reg1028 ?
          {($unsigned(forvar1026[(5'h10):(1'h1)]) - ((reg1030 >= forvar1026) | $unsigned(reg1029)))} : wire1023[(4'hc):(2'h3)]);
    end
  assign wire1033 = reg1028;
  module1034 modinst1059 (.wire1036(reg1031), .wire1035(reg1029), .clk(clk), .wire1038(reg1027), .y(wire1058), .wire1037(forvar1026));
  assign wire1060 = (+wire1022);
  always
    @(posedge clk) begin
      for (forvar1061 = (1'h0); (forvar1061 < (2'h2)); forvar1061 = (forvar1061 + (1'h1)))
        begin
          reg1062 <= ($unsigned({((wire1060 + reg1030) ?
                      wire1033 : $signed(wire1023))}) ?
              {(~reg1027)} : reg1029[(4'ha):(1'h0)]);
          reg1063 = $signed(((~($signed(reg1032) > wire1023)) <<< (&$unsigned(wire1022))));
          reg1064 <= $unsigned(wire1023[(3'h5):(1'h0)]);
          reg1065 <= $signed($signed({wire1058[(4'he):(4'ha)],
              forvar1061[(1'h0):(1'h0)]}));
        end
      for (forvar1066 = (1'h0); (forvar1066 < (2'h2)); forvar1066 = (forvar1066 + (1'h1)))
        begin
          for (forvar1067 = (1'h0); (forvar1067 < (1'h0)); forvar1067 = (forvar1067 + (1'h1)))
            begin
              reg1068 <= (!$signed($signed({wire1033,
                  (wire1033 ? reg1063 : (8'hb4))})));
              reg1069 = (^~$signed($unsigned($unsigned(wire1058))));
              reg1070 <= $unsigned(reg1029);
            end
          reg1071 = {(~|$unsigned((~^$unsigned(wire1021))))};
          reg1072 <= $unsigned($signed(reg1027));
          reg1073 <= {{reg1062}, {$signed((reg1030 != forvar1066))}};
        end
      reg1074 = (reg1062 ?
          reg1064 : ((reg1027 ?
                  ((reg1069 ? reg1071 : reg1030) ?
                      (&forvar1066) : (reg1071 ^~ reg1068)) : ($unsigned(reg1072) <<< reg1068[(5'h10):(4'hf)])) ?
              $unsigned(((8'ha7) * ((8'h9c) ? wire1058 : reg1025))) : reg1030));
    end
  assign wire1075 = reg1068[(2'h2):(2'h2)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1034  (y, clk, wire1038, wire1037, wire1036, wire1035);
  output wire [(32'he7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire1038;
  input wire signed [(3'h4):(1'h0)] wire1037;
  input wire [(4'ha):(1'h0)] wire1036;
  input wire [(5'h12):(1'h0)] wire1035;
  wire signed [(5'h12):(1'h0)] wire1057;
  wire signed [(4'he):(1'h0)] wire1056;
  reg [(2'h2):(1'h0)] reg1055 = (1'h0);
  reg [(4'hd):(1'h0)] reg1054 = (1'h0);
  reg [(4'hf):(1'h0)] reg1053 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1052 = (1'h0);
  reg [(4'hf):(1'h0)] reg1051 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1050 = (1'h0);
  reg [(5'h10):(1'h0)] reg1049 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1048 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1047 = (1'h0);
  reg [(2'h3):(1'h0)] reg1046 = (1'h0);
  reg [(4'hd):(1'h0)] reg1045 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1044 = (1'h0);
  reg [(3'h4):(1'h0)] reg1043 = (1'h0);
  wire [(4'ha):(1'h0)] wire1042;
  wire signed [(5'h10):(1'h0)] wire1041;
  reg signed [(5'h12):(1'h0)] reg1040 = (1'h0);
  reg [(5'h15):(1'h0)] reg1039 = (1'h0);
  assign y = {wire1057,
                 wire1056,
                 reg1055,
                 reg1054,
                 reg1053,
                 forvar1052,
                 reg1051,
                 reg1050,
                 reg1049,
                 reg1048,
                 reg1047,
                 reg1046,
                 reg1045,
                 reg1044,
                 reg1043,
                 wire1042,
                 wire1041,
                 reg1040,
                 reg1039,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1039 <= ($unsigned(wire1037) ?
          $signed({(-$unsigned((8'hb5)))}) : wire1038);
      reg1040 <= ($signed(wire1035[(4'hb):(2'h2)]) & $unsigned(wire1035[(3'h6):(3'h4)]));
    end
  assign wire1041 = $unsigned(($signed($signed((wire1036 ?
                        wire1037 : reg1039))) << $unsigned((+wire1035[(2'h2):(1'h0)]))));
  assign wire1042 = $unsigned(wire1041[(3'h5):(1'h0)]);
  always
    @(posedge clk) begin
      reg1043 <= {{wire1038[(4'h8):(3'h7)], wire1035},
          $unsigned((&$signed((~&wire1036))))};
      reg1044 = wire1037;
      reg1045 <= $signed((7'h42));
      reg1046 <= $signed(wire1036);
      reg1047 <= ($signed(((~|$unsigned((8'haa))) >> reg1046)) + (($signed((~|wire1037)) ?
          ($unsigned(reg1043) ?
              $unsigned(reg1040) : {wire1038}) : $unsigned({reg1045,
              (8'ha1)})) < (&{(^~wire1035)})));
    end
  always
    @(posedge clk) begin
      reg1048 = $unsigned((wire1041[(4'hf):(1'h0)] & (~^reg1047[(4'h8):(1'h1)])));
      reg1049 <= $unsigned((wire1037[(1'h1):(1'h1)] ^ $signed(((wire1038 >>> wire1036) ?
          $unsigned(reg1039) : reg1047))));
      reg1050 <= (-$signed(wire1035[(4'hc):(2'h3)]));
      reg1051 = reg1045;
      for (forvar1052 = (1'h0); (forvar1052 < (2'h2)); forvar1052 = (forvar1052 + (1'h1)))
        begin
          reg1053 <= reg1047;
          reg1054 <= ($signed((-reg1049)) ?
              (^{(~^wire1041)}) : $unsigned($signed($unsigned((wire1037 | wire1041)))));
          reg1055 <= reg1045;
        end
    end
  assign wire1056 = {(~&(-(8'ha2))),
                        ($unsigned($unsigned((|reg1045))) > {$signed({reg1045,
                                (8'hb5)})})};
  assign wire1057 = (($unsigned((&{reg1040, reg1054})) ?
                            (~{$unsigned(wire1042),
                                $unsigned(reg1051)}) : reg1044[(1'h1):(1'h1)]) ?
                        reg1049 : reg1047[(2'h3):(1'h1)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1919  (y, clk, wire1924, wire1923, wire1922, wire1921, wire1920);
  output wire [(32'h1dd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire1924;
  input wire [(5'h15):(1'h0)] wire1923;
  input wire signed [(5'h14):(1'h0)] wire1922;
  input wire signed [(4'hf):(1'h0)] wire1921;
  input wire signed [(5'h14):(1'h0)] wire1920;
  wire signed [(4'he):(1'h0)] wire2662;
  reg [(3'h4):(1'h0)] reg2661 = (1'h0);
  reg [(3'h4):(1'h0)] reg2660 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2659 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2658 = (1'h0);
  reg [(4'hf):(1'h0)] reg2657 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2656 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2655 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2654 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2653 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2652 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2651 = (1'h0);
  reg [(4'hd):(1'h0)] reg2650 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2649 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2648 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2647 = (1'h0);
  reg [(4'h9):(1'h0)] reg2646 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2645 = (1'h0);
  reg [(4'he):(1'h0)] forvar2644 = (1'h0);
  reg [(5'h12):(1'h0)] reg2643 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar2642 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2641 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2640 = (1'h0);
  reg [(3'h7):(1'h0)] reg2639 = (1'h0);
  reg [(4'hb):(1'h0)] reg2638 = (1'h0);
  reg [(5'h15):(1'h0)] reg2637 = (1'h0);
  reg [(3'h5):(1'h0)] reg2636 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2635 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2634 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2633 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2632 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2631 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire2630;
  wire signed [(4'he):(1'h0)] wire2170;
  wire [(4'ha):(1'h0)] wire1929;
  wire signed [(5'h13):(1'h0)] wire1928;
  reg [(4'he):(1'h0)] reg1927 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1926 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1925 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire2172;
  wire signed [(5'h14):(1'h0)] wire2628;
  assign y = {wire2662,
                 reg2661,
                 reg2660,
                 reg2659,
                 reg2658,
                 reg2657,
                 reg2656,
                 forvar2655,
                 reg2654,
                 forvar2653,
                 reg2652,
                 reg2651,
                 reg2650,
                 reg2649,
                 reg2648,
                 reg2647,
                 reg2646,
                 reg2645,
                 forvar2644,
                 reg2643,
                 forvar2642,
                 reg2641,
                 forvar2640,
                 reg2639,
                 reg2638,
                 reg2637,
                 reg2636,
                 forvar2635,
                 forvar2634,
                 reg2633,
                 reg2632,
                 forvar2631,
                 wire2630,
                 wire2170,
                 wire1929,
                 wire1928,
                 reg1927,
                 reg1926,
                 reg1925,
                 wire2172,
                 wire2628,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1925 <= wire1923;
    end
  always
    @(posedge clk) begin
      reg1926 <= ((|$unsigned((-reg1925[(4'hf):(4'hf)]))) ?
          (({$signed(wire1920)} ?
              {{reg1925, (8'ha1)}, $unsigned(wire1924)} : {(wire1921 ?
                      reg1925 : reg1925),
                  (wire1922 | reg1925)}) == {wire1921,
              ((~^wire1922) ?
                  $unsigned(wire1920) : $unsigned(wire1922))}) : $unsigned(reg1925));
      reg1927 <= $unsigned((&(~|wire1924)));
    end
  assign wire1928 = wire1920;
  assign wire1929 = (&((~^($unsigned(wire1924) >>> ((8'hb1) ?
                        wire1921 : wire1924))) * $unsigned(wire1928[(3'h5):(2'h3)])));
  module1930 modinst2171 (wire2170, clk, wire1922, wire1923, reg1926, wire1920, wire1929);
  assign wire2172 = $unsigned(wire1922[(5'h13):(4'he)]);
  module2173 modinst2629 (.clk(clk), .wire2174(reg1926), .y(wire2628), .wire2175(wire1928), .wire2178(wire2172), .wire2177(reg1927), .wire2176(wire1920));
  assign wire2630 = wire1920[(4'he):(4'hd)];
  always
    @(posedge clk) begin
      for (forvar2631 = (1'h0); (forvar2631 < (3'h4)); forvar2631 = (forvar2631 + (1'h1)))
        begin
          reg2632 <= $unsigned((~&wire1924[(2'h2):(1'h0)]));
          reg2633 <= (+$signed($unsigned($signed((wire2172 + wire1921)))));
        end
      for (forvar2634 = (1'h0); (forvar2634 < (1'h1)); forvar2634 = (forvar2634 + (1'h1)))
        begin
          for (forvar2635 = (1'h0); (forvar2635 < (1'h1)); forvar2635 = (forvar2635 + (1'h1)))
            begin
              reg2636 <= reg2633;
              reg2637 <= $signed(reg2633[(3'h4):(2'h2)]);
              reg2638 <= (($unsigned(wire1928[(4'ha):(4'h8)]) ?
                  (($unsigned(reg1925) ?
                          (wire1922 ?
                              wire2172 : wire1920) : reg2636[(2'h2):(2'h2)]) ?
                      ((wire2628 || (7'h41)) ^~ (~reg2633)) : ((reg1926 ^ wire2628) ?
                          forvar2631[(2'h3):(1'h1)] : reg1927)) : ((((8'hb4) || reg1925) ?
                          $unsigned(wire1929) : $signed(wire2170)) ?
                      (&(reg2633 && forvar2635)) : ($signed((8'ha9)) << (reg2637 * reg2637)))) <= reg2637);
              reg2639 <= $unsigned($unsigned((reg1927[(4'hb):(4'ha)] | reg1926)));
            end
          for (forvar2640 = (1'h0); (forvar2640 < (3'h4)); forvar2640 = (forvar2640 + (1'h1)))
            begin
              reg2641 = $signed((+wire1922[(5'h14):(5'h11)]));
            end
          for (forvar2642 = (1'h0); (forvar2642 < (3'h4)); forvar2642 = (forvar2642 + (1'h1)))
            begin
              reg2643 <= wire1921;
            end
          for (forvar2644 = (1'h0); (forvar2644 < (3'h4)); forvar2644 = (forvar2644 + (1'h1)))
            begin
              reg2645 <= wire1921;
              reg2646 <= $signed(($signed($signed((reg2638 * wire1928))) <= ($signed(wire1924) ?
                  (((8'h9e) ? (8'h9e) : wire1928) ?
                      (&forvar2631) : $unsigned(wire1921)) : (^~(~wire2172)))));
              reg2647 <= (((reg1927 ?
                  reg2636 : ($unsigned(forvar2644) ?
                      (forvar2635 ?
                          wire2172 : reg1926) : reg2638[(4'h9):(2'h3)])) >>> reg2636[(1'h1):(1'h1)]) != $signed((|$unsigned((reg2646 ?
                  (8'hbb) : forvar2640)))));
              reg2648 <= wire2172[(4'hc):(3'h5)];
            end
        end
      reg2649 = wire1923[(4'hf):(3'h5)];
      reg2650 = {wire1920[(3'h7):(3'h7)]};
      reg2651 <= ((+$unsigned(forvar2642[(1'h0):(1'h0)])) - reg1927[(4'ha):(2'h2)]);
    end
  always
    @(posedge clk) begin
      reg2652 <= $unsigned((wire1921[(4'h9):(1'h0)] && reg2632));
      for (forvar2653 = (1'h0); (forvar2653 < (1'h1)); forvar2653 = (forvar2653 + (1'h1)))
        begin
          reg2654 <= wire2172;
          for (forvar2655 = (1'h0); (forvar2655 < (1'h1)); forvar2655 = (forvar2655 + (1'h1)))
            begin
              reg2656 <= ((!wire1924) ?
                  {$signed({reg2633, $unsigned(reg2648)}),
                      (reg2647 ~^ {wire1920[(2'h2):(2'h2)],
                          (forvar2655 ?
                              wire1929 : wire1924)})} : (wire1921 >> $unsigned(reg2650)));
              reg2657 <= (^~reg2638);
              reg2658 = $signed((+wire2630[(3'h6):(3'h5)]));
              reg2659 <= {(8'ha0)};
            end
          reg2660 <= (((7'h41) != (reg2638 ^~ (wire2170[(2'h2):(1'h1)] ?
              (wire2628 ? forvar2640 : wire2170) : {reg2648,
                  reg1927}))) || $signed(((&(wire1923 ? reg1927 : (8'ha9))) ?
              (reg2650 ?
                  (-wire2628) : $signed((8'hb7))) : reg2637[(4'hb):(3'h7)])));
        end
      reg2661 <= ({$unsigned($signed($unsigned((8'haa)))), wire2630} ?
          reg2654 : $unsigned({{wire2630}}));
    end
  assign wire2662 = forvar2653;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1702
#( parameter param1888 = ((8'ha4) ? (~^({((8'hb7) < (8'ha0)), (^~(8'hbf))} ? (|(8'h9e)) : (((8'hb1) < (8'had)) ? (-(8'h9c)) : (!(8'hab))))) : ((~^{((8'ha9) ? (8'ha2) : (8'hb6)), (8'hae)}) ? ({{(8'ha1)}} | (((8'hb6) ? (7'h42) : (8'ha8)) ? (|(8'ha6)) : ((8'h9e) ? (8'ha8) : (8'hbd)))) : ((!{(7'h44), (8'hb3)}) & (((8'haf) ? (8'ha1) : (8'ha5)) + ((8'h9d) ? (7'h43) : (8'h9c))))))
, parameter param1889 = param1888 )
(y, clk, wire1703, wire1704, wire1705, wire1706);
  output wire [(32'hb1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire1703;
  input wire signed [(4'hb):(1'h0)] wire1704;
  input wire [(4'hd):(1'h0)] wire1705;
  input wire [(5'h13):(1'h0)] wire1706;
  wire signed [(2'h2):(1'h0)] wire1887;
  reg [(5'h14):(1'h0)] reg1707 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire1708;
  reg [(5'h10):(1'h0)] reg1709 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1710 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1711 = (1'h0);
  reg [(2'h2):(1'h0)] reg1712 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1713 = (1'h0);
  reg [(5'h15):(1'h0)] reg1714 = (1'h0);
  reg [(5'h14):(1'h0)] reg1715 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1716 = (1'h0);
  reg [(4'he):(1'h0)] reg1717 = (1'h0);
  wire [(3'h6):(1'h0)] wire1885;
  assign y = {wire1887,
                 reg1707,
                 wire1708,
                 reg1709,
                 reg1710,
                 forvar1711,
                 reg1712,
                 reg1713,
                 reg1714,
                 reg1715,
                 reg1716,
                 reg1717,
                 wire1885,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1707 <= $unsigned($signed(wire1704));
    end
  assign wire1708 = $unsigned($signed(wire1703));
  always
    @(posedge clk) begin
      reg1709 = wire1705[(4'h9):(3'h4)];
      reg1710 <= $signed($signed($unsigned($signed(((8'ha3) >> wire1705)))));
      for (forvar1711 = (1'h0); (forvar1711 < (1'h1)); forvar1711 = (forvar1711 + (1'h1)))
        begin
          reg1712 <= ((|$signed(wire1706)) >> $signed(($unsigned(wire1704) >> wire1704)));
          reg1713 = wire1705[(4'hd):(2'h2)];
          reg1714 <= ({wire1704[(1'h1):(1'h0)]} & forvar1711);
          reg1715 = $signed((~(~(+((7'h40) ? reg1709 : reg1712)))));
          reg1716 = forvar1711[(4'ha):(4'h9)];
        end
      reg1717 <= ((wire1708 | wire1704) == ($signed($signed((reg1715 ?
          wire1705 : reg1709))) < wire1703[(3'h6):(1'h0)]));
    end
  module1718 modinst1886 (wire1885, clk, reg1715, wire1708, reg1710, reg1714, reg1713);
  assign wire1887 = $signed((^~{reg1710[(4'h9):(3'h6)],
                        $unsigned($unsigned(wire1706))}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1653
#( parameter param1686 = (({(-((7'h44) * (8'ha0))), (-((8'hb0) ^ (8'hb1)))} ~^ ((((8'haa) <= (8'hbc)) + (+(8'ha9))) ? (-((8'ha8) ^ (8'hb5))) : (((8'hbd) > (8'ha9)) * (-(8'h9c))))) ? ({(~((8'ha2) * (8'hbf)))} - (~&(((8'h9f) ? (8'ha3) : (8'hba)) ? ((8'hbc) || (7'h40)) : (8'ha3)))) : (((((8'ha0) ? (7'h43) : (8'ha5)) ? ((8'ha4) ? (8'hba) : (8'hab)) : ((7'h44) || (8'h9c))) >>> {(!(8'hbe)), ((8'h9c) ? (8'hbe) : (8'ha1))}) ? ({((8'hb0) ? (8'hb3) : (8'hb4))} || (((8'ha2) | (8'h9f)) ? ((8'ha5) & (8'hba)) : ((8'hae) != (7'h44)))) : {{((8'hab) ? (7'h44) : (8'ha3))}})) )
(y, clk, wire1658, wire1657, wire1656, wire1655, wire1654);
  output wire [(32'h120):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire1658;
  input wire signed [(5'h12):(1'h0)] wire1657;
  input wire [(3'h6):(1'h0)] wire1656;
  input wire signed [(4'h9):(1'h0)] wire1655;
  input wire signed [(4'h8):(1'h0)] wire1654;
  reg signed [(4'ha):(1'h0)] reg1685 = (1'h0);
  reg [(5'h15):(1'h0)] reg1684 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1683 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1682 = (1'h0);
  wire [(2'h2):(1'h0)] wire1681;
  reg signed [(4'hc):(1'h0)] reg1680 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1679 = (1'h0);
  reg [(5'h15):(1'h0)] reg1678 = (1'h0);
  reg [(5'h14):(1'h0)] reg1677 = (1'h0);
  reg [(4'hb):(1'h0)] reg1676 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1675 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1674 = (1'h0);
  reg [(4'he):(1'h0)] reg1673 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1672 = (1'h0);
  reg [(3'h6):(1'h0)] reg1671 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1670 = (1'h0);
  wire [(5'h12):(1'h0)] wire1669;
  wire signed [(2'h3):(1'h0)] wire1668;
  reg signed [(2'h3):(1'h0)] reg1667 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1666 = (1'h0);
  reg [(5'h14):(1'h0)] reg1665 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1664 = (1'h0);
  reg [(4'hf):(1'h0)] reg1663 = (1'h0);
  reg [(3'h7):(1'h0)] reg1662 = (1'h0);
  reg [(5'h12):(1'h0)] reg1661 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1660 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1659 = (1'h0);
  assign y = {reg1685,
                 reg1684,
                 reg1683,
                 reg1682,
                 wire1681,
                 reg1680,
                 reg1679,
                 reg1678,
                 reg1677,
                 reg1676,
                 reg1675,
                 reg1674,
                 reg1673,
                 forvar1672,
                 reg1671,
                 reg1670,
                 wire1669,
                 wire1668,
                 reg1667,
                 reg1666,
                 reg1665,
                 reg1664,
                 reg1663,
                 reg1662,
                 reg1661,
                 forvar1660,
                 reg1659,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1659 <= $unsigned(wire1657[(3'h4):(3'h4)]);
      if (wire1655[(3'h4):(2'h2)])
        begin
          for (forvar1660 = (1'h0); (forvar1660 < (2'h2)); forvar1660 = (forvar1660 + (1'h1)))
            begin
              reg1661 <= forvar1660;
              reg1662 <= forvar1660;
              reg1663 <= wire1658;
              reg1664 <= (($signed($signed($signed(reg1663))) == (((~^forvar1660) ?
                      $unsigned(wire1656) : {wire1657}) ?
                  ((reg1659 != wire1657) != (reg1661 - forvar1660)) : ((8'ha0) ~^ (8'hbc)))) || (^$signed(({wire1654,
                      wire1655} ?
                  (~|wire1656) : $signed(wire1656)))));
              reg1665 <= (($signed($unsigned($signed(reg1661))) ?
                  $unsigned((8'hb9)) : $unsigned(({reg1663} ?
                      wire1657[(1'h0):(1'h0)] : forvar1660[(1'h1):(1'h1)]))) | (^~(8'hbe)));
            end
          reg1666 <= ($unsigned(reg1659) ?
              wire1654 : {wire1656[(3'h5):(1'h0)]});
          reg1667 = (((8'hb2) < (($unsigned(reg1663) >>> reg1661[(3'h7):(3'h6)]) + $unsigned((reg1662 ?
                  forvar1660 : reg1662)))) ?
              wire1654[(3'h7):(2'h3)] : $signed($signed({(wire1655 << reg1666),
                  {reg1659}})));
        end
      else
        begin
          for (forvar1660 = (1'h0); (forvar1660 < (1'h0)); forvar1660 = (forvar1660 + (1'h1)))
            begin
              reg1661 <= (((8'hab) + $signed((8'ha9))) <= $unsigned($signed({(8'hb4)})));
              reg1662 = $signed($signed(reg1661[(4'h8):(2'h2)]));
              reg1663 <= {($signed(reg1662[(2'h3):(1'h1)]) ^ (reg1663[(3'h6):(3'h6)] ~^ {(reg1665 * reg1666),
                      $signed(reg1666)})),
                  reg1659};
            end
          reg1664 <= ($signed(forvar1660[(1'h1):(1'h0)]) ?
              ((8'ha1) <<< reg1666) : $unsigned((~&(!reg1663[(4'hc):(3'h7)]))));
          reg1665 <= ((8'hbc) ^ reg1665[(4'hf):(1'h0)]);
        end
    end
  assign wire1668 = reg1659;
  assign wire1669 = ($signed((^(((8'hb6) <= (8'hb7)) ~^ (~^forvar1660)))) + ((reg1659 ?
                            ((wire1656 ?
                                wire1654 : reg1661) != (reg1665 * (8'ha6))) : reg1667) ?
                        $unsigned($signed(wire1658)) : (~&((8'hbf) ?
                            {wire1668, wire1658} : $signed(wire1655)))));
  always
    @(posedge clk) begin
      reg1670 <= $unsigned($signed(((+reg1667[(1'h1):(1'h0)]) ?
          ({wire1656} ?
              $unsigned(reg1663) : (reg1666 >>> reg1663)) : $signed((|wire1668)))));
      reg1671 = wire1658;
      for (forvar1672 = (1'h0); (forvar1672 < (2'h3)); forvar1672 = (forvar1672 + (1'h1)))
        begin
          reg1673 <= wire1656;
          reg1674 <= wire1656[(3'h4):(3'h4)];
        end
      reg1675 = ((reg1664 != (!($signed((8'hb9)) + ((8'ha3) || reg1662)))) ?
          ((~^reg1674) & $unsigned(wire1656[(1'h1):(1'h1)])) : wire1668);
      reg1676 <= reg1665;
    end
  always
    @(posedge clk) begin
      reg1677 = reg1674;
      reg1678 <= forvar1672[(2'h2):(1'h1)];
      reg1679 <= ({wire1654} ?
          reg1675[(2'h2):(2'h2)] : (($signed(wire1657[(4'h8):(3'h7)]) ?
                  $signed(reg1664) : $signed(forvar1660)) ?
              $signed(reg1675[(1'h0):(1'h0)]) : wire1654));
    end
  always
    @(posedge clk) begin
      reg1680 <= (forvar1672[(2'h2):(1'h0)] ~^ $signed(wire1655));
    end
  assign wire1681 = (^$signed((7'h43)));
  always
    @(posedge clk) begin
      reg1682 <= forvar1672[(1'h1):(1'h1)];
    end
  always
    @(posedge clk) begin
      reg1683 <= (|wire1655[(3'h7):(3'h7)]);
      reg1684 <= reg1678[(3'h6):(3'h5)];
    end
  always
    @(posedge clk) begin
      reg1685 = (&reg1667);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1167  (y, clk, wire1168, wire1169, wire1170, wire1171);
  output wire [(32'h24d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire1168;
  input wire signed [(5'h14):(1'h0)] wire1169;
  input wire signed [(4'h8):(1'h0)] wire1170;
  input wire [(3'h4):(1'h0)] wire1171;
  reg signed [(5'h14):(1'h0)] reg1628 = (1'h0);
  reg [(3'h6):(1'h0)] reg1627 = (1'h0);
  reg [(3'h5):(1'h0)] reg1626 = (1'h0);
  wire [(4'h9):(1'h0)] wire1625;
  wire [(4'hf):(1'h0)] wire1623;
  wire signed [(5'h12):(1'h0)] wire1460;
  reg [(5'h13):(1'h0)] reg1459 = (1'h0);
  wire [(5'h11):(1'h0)] wire1458;
  wire [(3'h5):(1'h0)] wire1456;
  wire signed [(5'h14):(1'h0)] wire1172;
  reg [(4'hd):(1'h0)] reg1173 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1174 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1175 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1176 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1177 = (1'h0);
  reg [(3'h7):(1'h0)] reg1178 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1179 = (1'h0);
  reg [(4'h8):(1'h0)] reg1180 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1181 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1182 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1183 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1184 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1185 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1186 = (1'h0);
  reg [(3'h7):(1'h0)] reg1187 = (1'h0);
  reg [(5'h15):(1'h0)] reg1188 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1189 = (1'h0);
  reg [(3'h6):(1'h0)] reg1190 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1191 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1192 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1193 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1194 = (1'h0);
  reg [(5'h10):(1'h0)] reg1195 = (1'h0);
  reg [(5'h11):(1'h0)] reg1196 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1197 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1198 = (1'h0);
  reg [(5'h10):(1'h0)] reg1199 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1200 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1201 = (1'h0);
  reg [(3'h7):(1'h0)] reg1202 = (1'h0);
  reg [(4'hf):(1'h0)] reg1203 = (1'h0);
  reg [(5'h14):(1'h0)] reg1204 = (1'h0);
  wire [(3'h7):(1'h0)] wire1205;
  wire [(3'h5):(1'h0)] wire1206;
  wire [(2'h3):(1'h0)] wire1207;
  wire signed [(3'h4):(1'h0)] wire1313;
  assign y = {reg1628,
                 reg1627,
                 reg1626,
                 wire1625,
                 wire1623,
                 wire1460,
                 reg1459,
                 wire1458,
                 wire1456,
                 wire1172,
                 reg1173,
                 forvar1174,
                 reg1175,
                 reg1176,
                 reg1177,
                 reg1178,
                 reg1179,
                 reg1180,
                 reg1181,
                 forvar1182,
                 forvar1183,
                 reg1184,
                 reg1185,
                 reg1186,
                 reg1187,
                 reg1188,
                 forvar1189,
                 reg1190,
                 reg1191,
                 forvar1192,
                 forvar1193,
                 reg1194,
                 reg1195,
                 reg1196,
                 forvar1197,
                 reg1198,
                 reg1199,
                 forvar1200,
                 reg1201,
                 reg1202,
                 reg1203,
                 reg1204,
                 wire1205,
                 wire1206,
                 wire1207,
                 wire1313,
                 (1'h0)};
  assign wire1172 = wire1171;
  always
    @(posedge clk) begin
      reg1173 = wire1169[(5'h14):(5'h14)];
      for (forvar1174 = (1'h0); (forvar1174 < (2'h3)); forvar1174 = (forvar1174 + (1'h1)))
        begin
          reg1175 = wire1168[(4'h9):(4'h8)];
        end
      reg1176 <= $signed(reg1175);
      reg1177 = (8'hbd);
      reg1178 <= $signed($unsigned(((forvar1174 & ((8'hae) ?
          wire1168 : reg1176)) && (((8'hb7) - (8'ha1)) ?
          ((8'ha6) && reg1173) : (wire1169 ? wire1170 : reg1177)))));
    end
  always
    @(posedge clk) begin
      reg1179 <= $signed(($signed(((wire1169 <= wire1172) ?
              (forvar1174 * wire1171) : (wire1172 > wire1172))) ?
          {(8'ha5), $signed((reg1178 & (8'hbb)))} : reg1176));
    end
  always
    @(posedge clk) begin
      reg1180 = $unsigned(($unsigned(forvar1174) < $unsigned($signed(wire1169))));
      reg1181 = (reg1180 ?
          (reg1178 ?
              (-((wire1171 ?
                  wire1170 : reg1173) == (|(8'ha3)))) : ($unsigned(reg1179[(4'h8):(3'h6)]) ?
                  (~|(wire1172 ? reg1176 : (8'hb1))) : (~^(reg1180 ?
                      (7'h43) : reg1176)))) : $unsigned(forvar1174[(3'h4):(1'h1)]));
      for (forvar1182 = (1'h0); (forvar1182 < (1'h1)); forvar1182 = (forvar1182 + (1'h1)))
        begin
          for (forvar1183 = (1'h0); (forvar1183 < (2'h3)); forvar1183 = (forvar1183 + (1'h1)))
            begin
              reg1184 <= ((($signed($unsigned(wire1169)) ?
                      wire1171[(3'h4):(1'h1)] : ($unsigned(reg1175) * reg1177[(4'hf):(4'h8)])) == ($unsigned((^~reg1180)) | (^(~&forvar1182)))) ?
                  ((($unsigned(reg1179) ?
                              (wire1169 >= (8'hb5)) : (reg1176 > reg1178)) ?
                          {$signed(wire1169)} : ($unsigned((8'ha4)) ?
                              (forvar1183 ? wire1171 : (8'hbb)) : {wire1168})) ?
                      reg1178[(2'h3):(1'h1)] : ($signed(wire1169) ?
                          (^((8'haf) ?
                              forvar1174 : forvar1182)) : $signed((^(8'ha2))))) : ($signed(((|reg1177) > $unsigned(reg1177))) ?
                      (^~{reg1177[(4'hd):(4'hd)]}) : (!(~|(forvar1174 ?
                          reg1175 : reg1181)))));
              reg1185 = (reg1177 ?
                  (reg1177 > ($unsigned((wire1172 ^~ reg1173)) ?
                      (~&$unsigned(reg1184)) : (wire1171[(1'h1):(1'h1)] ?
                          (forvar1174 ? wire1169 : reg1175) : ((7'h43) ?
                              wire1172 : forvar1182)))) : $signed(reg1181));
              reg1186 = reg1181;
            end
          reg1187 <= $unsigned((8'ha1));
          reg1188 <= reg1173[(3'h7):(3'h5)];
          for (forvar1189 = (1'h0); (forvar1189 < (1'h1)); forvar1189 = (forvar1189 + (1'h1)))
            begin
              reg1190 <= (reg1173 && {(((wire1170 + wire1172) <<< forvar1189[(1'h1):(1'h0)]) ?
                      (^~reg1187[(3'h4):(2'h3)]) : (~|$signed(reg1178)))});
            end
          reg1191 <= $signed(reg1188);
        end
      for (forvar1192 = (1'h0); (forvar1192 < (3'h4)); forvar1192 = (forvar1192 + (1'h1)))
        begin
          for (forvar1193 = (1'h0); (forvar1193 < (1'h0)); forvar1193 = (forvar1193 + (1'h1)))
            begin
              reg1194 <= (~^$unsigned($signed((&(wire1172 || reg1177)))));
              reg1195 = $unsigned((&$signed($signed(reg1180[(3'h7):(3'h5)]))));
              reg1196 = (~((~|((&reg1181) ?
                      (forvar1192 ? reg1173 : reg1187) : (reg1185 ?
                          reg1185 : (8'hbd)))) ?
                  {wire1168} : $signed((forvar1182 ?
                      $signed(wire1172) : $signed(forvar1193)))));
            end
          for (forvar1197 = (1'h0); (forvar1197 < (1'h0)); forvar1197 = (forvar1197 + (1'h1)))
            begin
              reg1198 <= reg1190[(2'h2):(1'h1)];
            end
          reg1199 <= forvar1182;
          for (forvar1200 = (1'h0); (forvar1200 < (2'h2)); forvar1200 = (forvar1200 + (1'h1)))
            begin
              reg1201 <= (~($signed($signed($signed(reg1173))) ?
                  $unsigned(($signed(forvar1200) ?
                      $unsigned((8'ha7)) : reg1178)) : $signed(reg1185)));
              reg1202 <= (~$unsigned($unsigned((^reg1187[(3'h7):(3'h5)]))));
              reg1203 = reg1184[(3'h6):(3'h5)];
              reg1204 <= ($unsigned((8'ha9)) ?
                  (($signed($signed(forvar1182)) ?
                          (-((8'hbc) | wire1171)) : (~|{reg1196})) ?
                      reg1190[(2'h3):(1'h0)] : reg1202[(3'h5):(2'h3)]) : wire1170);
            end
        end
    end
  assign wire1205 = ($unsigned((|((reg1202 == reg1188) ?
                        (^(8'ha2)) : ((8'hb3) ?
                            forvar1182 : reg1203)))) ^ $unsigned(((8'hb6) ?
                        (((7'h44) ? (8'ha6) : reg1178) ?
                            {forvar1182} : (reg1203 ?
                                reg1190 : reg1184)) : $signed(reg1195))));
  assign wire1206 = reg1184;
  assign wire1207 = ($unsigned((-wire1169)) ?
                        ((forvar1193[(1'h1):(1'h0)] - (wire1169 >>> $signed(forvar1192))) <<< $signed(reg1187[(3'h4):(2'h2)])) : $unsigned(reg1198[(2'h2):(1'h1)]));
  module1208 modinst1314 (wire1313, clk, wire1172, forvar1192, forvar1200, wire1168, wire1169);
  module1315 modinst1457 (wire1456, clk, forvar1183, reg1204, forvar1174, reg1203);
  assign wire1458 = (~^wire1206);
  always
    @(posedge clk) begin
      reg1459 <= $unsigned({reg1195[(1'h1):(1'h1)], forvar1189});
    end
  assign wire1460 = wire1171[(1'h0):(1'h0)];
  module1461 modinst1624 (.wire1465(reg1175), .clk(clk), .wire1464(reg1181), .wire1462(reg1196), .wire1463(wire1169), .y(wire1623));
  assign wire1625 = (forvar1182 ?
                        $signed(((^((8'ha2) < reg1201)) ?
                            ($unsigned(reg1203) << $signed((8'hbe))) : (wire1170 <= $signed(reg1195)))) : $signed((wire1313 ?
                            ({(8'hbd), reg1186} ?
                                reg1181 : reg1196) : forvar1189[(2'h3):(2'h2)])));
  always
    @(posedge clk) begin
      reg1626 <= wire1168[(3'h4):(2'h2)];
      reg1627 = ($signed((-(wire1169[(3'h4):(2'h3)] | (reg1178 ?
              reg1187 : reg1196)))) ?
          $unsigned($unsigned(reg1194[(2'h2):(2'h2)])) : reg1196[(3'h7):(3'h7)]);
      reg1628 <= wire1171;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1461
#( parameter param1621 = (((^~((+(8'hb6)) && ((8'had) & (8'had)))) || ({(~|(8'ha7)), ((8'hb5) - (8'hbb))} ? {(&(8'haa)), {(8'h9e)}} : (((7'h42) & (8'h9e)) ? ((8'ha9) ? (8'hbf) : (8'hbf)) : (8'hb5)))) && (((+(8'h9e)) ? (!((8'ha5) ^~ (8'hbc))) : (((8'ha2) << (7'h42)) - (^~(8'h9f)))) >>> ((((8'ha9) | (8'haf)) ~^ (+(8'hbc))) >= (~^((8'hb5) - (8'ha8))))))
, parameter param1622 = ((8'hbf) ? ((|({param1621, param1621} >>> param1621)) ? (^~(+(param1621 && param1621))) : (&(8'haf))) : {((+(^~param1621)) << param1621)}) )
(y, clk, wire1465, wire1464, wire1463, wire1462);
  output wire [(32'h343):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire1465;
  input wire [(4'he):(1'h0)] wire1464;
  input wire signed [(5'h14):(1'h0)] wire1463;
  input wire [(5'h11):(1'h0)] wire1462;
  wire [(4'hb):(1'h0)] wire1620;
  wire [(5'h14):(1'h0)] wire1619;
  reg [(5'h12):(1'h0)] reg1618 = (1'h0);
  reg [(5'h12):(1'h0)] reg1617 = (1'h0);
  reg [(2'h3):(1'h0)] reg1616 = (1'h0);
  wire [(5'h14):(1'h0)] wire1615;
  wire [(4'h8):(1'h0)] wire1614;
  wire [(4'hf):(1'h0)] wire1613;
  reg signed [(4'h8):(1'h0)] reg1612 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1611 = (1'h0);
  reg [(5'h10):(1'h0)] reg1610 = (1'h0);
  reg [(5'h14):(1'h0)] reg1609 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1608 = (1'h0);
  reg [(5'h15):(1'h0)] reg1607 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1606 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1605 = (1'h0);
  reg [(4'he):(1'h0)] reg1604 = (1'h0);
  reg [(3'h6):(1'h0)] reg1603 = (1'h0);
  reg [(5'h14):(1'h0)] reg1602 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1601 = (1'h0);
  reg [(4'h8):(1'h0)] reg1600 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1599 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1598 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire1596;
  reg signed [(2'h2):(1'h0)] reg1551 = (1'h0);
  reg [(4'he):(1'h0)] reg1550 = (1'h0);
  reg [(3'h7):(1'h0)] reg1549 = (1'h0);
  reg [(3'h7):(1'h0)] reg1548 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1547 = (1'h0);
  reg [(4'hb):(1'h0)] reg1546 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1545 = (1'h0);
  reg [(5'h11):(1'h0)] reg1544 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1543 = (1'h0);
  reg [(5'h14):(1'h0)] reg1542 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1541 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1540 = (1'h0);
  reg [(2'h3):(1'h0)] reg1539 = (1'h0);
  reg [(4'hd):(1'h0)] reg1538 = (1'h0);
  reg [(4'hc):(1'h0)] reg1537 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1536 = (1'h0);
  reg [(5'h10):(1'h0)] reg1535 = (1'h0);
  reg [(2'h3):(1'h0)] reg1534 = (1'h0);
  reg [(4'hd):(1'h0)] reg1533 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1532 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1531 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1530 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1529 = (1'h0);
  reg [(3'h4):(1'h0)] reg1528 = (1'h0);
  wire [(4'h9):(1'h0)] wire1527;
  reg [(2'h3):(1'h0)] reg1526 = (1'h0);
  reg [(5'h14):(1'h0)] reg1525 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1524 = (1'h0);
  reg [(5'h13):(1'h0)] reg1523 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1522 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1521 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1520 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1519 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1518 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1517 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1516 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1515 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1514 = (1'h0);
  reg [(2'h3):(1'h0)] reg1513 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1512 = (1'h0);
  reg [(3'h4):(1'h0)] reg1511 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire1510;
  wire signed [(4'h8):(1'h0)] wire1508;
  wire signed [(5'h12):(1'h0)] wire1471;
  wire signed [(4'hd):(1'h0)] wire1470;
  reg signed [(3'h5):(1'h0)] reg1469 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1468 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1467 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1466 = (1'h0);
  assign y = {wire1620,
                 wire1619,
                 reg1618,
                 reg1617,
                 reg1616,
                 wire1615,
                 wire1614,
                 wire1613,
                 reg1612,
                 reg1611,
                 reg1610,
                 reg1609,
                 reg1608,
                 reg1607,
                 forvar1606,
                 forvar1605,
                 reg1604,
                 reg1603,
                 reg1602,
                 forvar1601,
                 reg1600,
                 reg1599,
                 reg1598,
                 wire1596,
                 reg1551,
                 reg1550,
                 reg1549,
                 reg1548,
                 forvar1547,
                 reg1546,
                 reg1545,
                 reg1544,
                 reg1543,
                 reg1542,
                 reg1541,
                 forvar1540,
                 reg1539,
                 reg1538,
                 reg1537,
                 forvar1536,
                 reg1535,
                 reg1534,
                 reg1533,
                 reg1532,
                 forvar1531,
                 reg1530,
                 forvar1529,
                 reg1528,
                 wire1527,
                 reg1526,
                 reg1525,
                 forvar1524,
                 reg1523,
                 reg1522,
                 reg1521,
                 reg1520,
                 reg1519,
                 reg1518,
                 reg1517,
                 reg1516,
                 reg1515,
                 forvar1514,
                 reg1513,
                 forvar1512,
                 reg1511,
                 wire1510,
                 wire1508,
                 wire1471,
                 wire1470,
                 reg1469,
                 reg1468,
                 forvar1467,
                 reg1466,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1466 <= {$signed(wire1462[(3'h6):(3'h5)]),
          $signed(wire1463[(5'h12):(4'ha)])};
      for (forvar1467 = (1'h0); (forvar1467 < (1'h1)); forvar1467 = (forvar1467 + (1'h1)))
        begin
          reg1468 = $unsigned((((wire1464[(4'h8):(3'h7)] < $signed((7'h44))) ?
              $unsigned($signed(reg1466)) : wire1465) == ($signed(((8'hb7) ^ wire1465)) ^~ (~&(^reg1466)))));
          reg1469 <= (forvar1467[(1'h1):(1'h0)] ?
              {(^~$signed((~wire1463)))} : reg1468);
        end
    end
  assign wire1470 = wire1462[(3'h4):(1'h1)];
  assign wire1471 = (+$unsigned((&$unsigned(reg1466))));
  module1472 modinst1509 (.clk(clk), .wire1473(wire1463), .wire1476(reg1468), .wire1475(wire1464), .wire1474(wire1471), .y(wire1508));
  assign wire1510 = wire1463;
  always
    @(posedge clk) begin
      reg1511 <= wire1470[(2'h2):(1'h0)];
      for (forvar1512 = (1'h0); (forvar1512 < (1'h0)); forvar1512 = (forvar1512 + (1'h1)))
        begin
          reg1513 <= $signed((!$signed(({wire1470, (8'hb2)} ?
              {wire1464, wire1465} : forvar1467[(1'h1):(1'h0)]))));
          for (forvar1514 = (1'h0); (forvar1514 < (3'h4)); forvar1514 = (forvar1514 + (1'h1)))
            begin
              reg1515 <= reg1466;
              reg1516 <= {(($signed(reg1469[(1'h0):(1'h0)]) || (!(wire1471 || wire1465))) ?
                      (7'h43) : {$signed(reg1466),
                          ($signed(wire1465) ^~ $unsigned(wire1462))}),
                  {$signed(reg1515[(1'h0):(1'h0)]),
                      $unsigned($unsigned(wire1462[(5'h11):(4'ha)]))}};
              reg1517 <= (!reg1516[(1'h1):(1'h1)]);
              reg1518 <= ($unsigned(wire1470[(3'h4):(1'h0)]) <<< ({wire1508[(3'h7):(2'h3)],
                      (|reg1517[(2'h3):(2'h3)])} ?
                  $signed(wire1463[(5'h12):(4'hf)]) : $signed($unsigned(forvar1514[(2'h3):(1'h1)]))));
              reg1519 <= (($signed({(wire1508 && forvar1467),
                          $unsigned(wire1508)}) ?
                      {$signed((^wire1464))} : reg1516) ?
                  ($unsigned(($signed(wire1462) >> $signed(wire1462))) >= $unsigned((~|$unsigned((8'hb9))))) : reg1517);
            end
          reg1520 <= ((reg1518[(4'he):(2'h2)] - $signed($signed((wire1465 ?
              wire1510 : (8'hb6))))) <= wire1462);
          reg1521 <= $unsigned(($unsigned(reg1511) && {wire1462,
              (forvar1512[(3'h7):(1'h0)] | (-(8'hbe)))}));
          reg1522 = ($signed({(~(+wire1470)),
              $unsigned(reg1468[(3'h4):(2'h2)])}) + (($signed(reg1513[(2'h2):(2'h2)]) ?
              ($signed(wire1463) ?
                  $unsigned((8'h9d)) : (8'ha8)) : (8'h9d)) != $signed($unsigned((reg1518 ?
              wire1510 : reg1520)))));
        end
      reg1523 <= reg1513[(2'h2):(1'h0)];
      for (forvar1524 = (1'h0); (forvar1524 < (3'h4)); forvar1524 = (forvar1524 + (1'h1)))
        begin
          reg1525 <= $unsigned((^(reg1517[(3'h4):(1'h0)] ?
              ($signed(forvar1524) ?
                  (|reg1519) : (8'ha2)) : reg1521[(3'h6):(2'h3)])));
          reg1526 <= wire1470;
        end
    end
  assign wire1527 = (wire1463[(1'h0):(1'h0)] >> (&$unsigned($signed((8'ha1)))));
  always
    @(posedge clk) begin
      reg1528 <= ((8'hb3) ?
          $signed($unsigned($signed(forvar1524[(1'h1):(1'h1)]))) : (8'hb2));
      for (forvar1529 = (1'h0); (forvar1529 < (3'h4)); forvar1529 = (forvar1529 + (1'h1)))
        begin
          reg1530 <= $signed((|forvar1529[(3'h4):(1'h1)]));
          for (forvar1531 = (1'h0); (forvar1531 < (1'h0)); forvar1531 = (forvar1531 + (1'h1)))
            begin
              reg1532 <= (-wire1463[(3'h4):(2'h3)]);
              reg1533 <= (|$unsigned((wire1462 << {forvar1514[(1'h0):(1'h0)],
                  reg1521[(2'h3):(1'h1)]})));
              reg1534 = {($unsigned($signed({reg1469})) ?
                      forvar1514[(3'h5):(3'h5)] : $signed(reg1520)),
                  $signed($unsigned({((8'hbb) >= (8'hac))}))};
            end
          reg1535 <= reg1523;
          for (forvar1536 = (1'h0); (forvar1536 < (3'h4)); forvar1536 = (forvar1536 + (1'h1)))
            begin
              reg1537 <= ((forvar1514[(1'h1):(1'h0)] ?
                  $unsigned((wire1470 ?
                      $signed(wire1508) : $signed(forvar1514))) : (-((~&forvar1531) < {wire1471,
                      reg1466}))) <<< (reg1519[(2'h3):(2'h3)] <<< ((reg1519[(2'h3):(2'h3)] ?
                  $unsigned(reg1469) : (&forvar1524)) ~^ $signed($signed(reg1530)))));
              reg1538 = {(((reg1522[(4'ha):(3'h7)] ?
                          {reg1466, reg1532} : (reg1522 ?
                              reg1511 : reg1516)) <<< forvar1536[(2'h2):(1'h1)]) ?
                      (-((forvar1536 ? reg1517 : (8'ha3)) ?
                          $unsigned(wire1463) : $unsigned(reg1466))) : (-wire1463[(4'h9):(3'h6)])),
                  $signed((+reg1516[(1'h1):(1'h0)]))};
              reg1539 <= $signed(reg1538[(1'h1):(1'h1)]);
            end
          for (forvar1540 = (1'h0); (forvar1540 < (2'h3)); forvar1540 = (forvar1540 + (1'h1)))
            begin
              reg1541 <= forvar1512[(2'h3):(2'h3)];
              reg1542 = $unsigned(((reg1513[(1'h1):(1'h1)] << (wire1471 ?
                      reg1530[(3'h7):(3'h7)] : (wire1464 ?
                          reg1468 : forvar1512))) ?
                  ((&reg1519[(1'h1):(1'h0)]) ?
                      reg1528 : forvar1514[(3'h5):(3'h5)]) : (wire1462 | reg1520[(1'h0):(1'h0)])));
              reg1543 = ({$unsigned(reg1516[(3'h4):(1'h1)])} ?
                  {{((!wire1463) ? wire1463 : forvar1512[(1'h1):(1'h1)]),
                          $unsigned({(7'h40)})},
                      $signed($signed(reg1534[(1'h1):(1'h0)]))} : {(^~forvar1529)});
              reg1544 = ($unsigned($signed((^~wire1510))) ?
                  ($signed(reg1523[(5'h13):(4'hd)]) ?
                      $unsigned($unsigned({wire1510})) : (wire1510[(4'hb):(4'ha)] & $signed($unsigned(wire1463)))) : $unsigned((&(+forvar1536))));
              reg1545 <= (^~reg1541);
            end
        end
      reg1546 = ((-(~($unsigned(reg1528) << (reg1528 ?
          reg1525 : reg1518)))) >= reg1520);
      for (forvar1547 = (1'h0); (forvar1547 < (2'h2)); forvar1547 = (forvar1547 + (1'h1)))
        begin
          reg1548 <= reg1532;
          reg1549 <= (!(!reg1523));
          reg1550 = {reg1518, wire1508[(3'h7):(2'h3)]};
        end
      reg1551 <= (^{wire1470, (8'hb7)});
    end
  module1552 modinst1597 (.wire1553(reg1546), .wire1554(reg1542), .clk(clk), .y(wire1596), .wire1556(reg1468), .wire1555(reg1525));
  always
    @(posedge clk) begin
      reg1598 <= $signed($unsigned($unsigned($signed(forvar1467[(3'h4):(1'h0)]))));
    end
  always
    @(posedge clk) begin
      reg1599 <= reg1537[(2'h3):(2'h2)];
      reg1600 = {(($signed($unsigned(reg1542)) ~^ (^$unsigned(reg1521))) ?
              reg1526[(1'h0):(1'h0)] : (^~{reg1519[(2'h2):(2'h2)],
                  $unsigned(reg1543)})),
          reg1522[(4'hf):(1'h0)]};
      for (forvar1601 = (1'h0); (forvar1601 < (3'h4)); forvar1601 = (forvar1601 + (1'h1)))
        begin
          reg1602 <= (((((+forvar1467) ?
                      (!(8'hac)) : (reg1513 > wire1463)) * {reg1543[(3'h4):(3'h4)]}) ?
                  (~^$signed((^~reg1534))) : reg1599[(1'h0):(1'h0)]) ?
              reg1518 : (-$signed(((+reg1542) ?
                  (forvar1547 ? reg1516 : (8'hba)) : (wire1470 ?
                      reg1537 : reg1533)))));
        end
      reg1603 <= (!(reg1545[(3'h5):(1'h1)] ?
          (+reg1545[(3'h4):(2'h3)]) : (((~&reg1550) + reg1600) ?
              $unsigned((~^reg1533)) : (~forvar1536[(4'hf):(4'hb)]))));
      reg1604 = ((~^(~^(^~(8'hb9)))) | reg1515[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      for (forvar1605 = (1'h0); (forvar1605 < (2'h2)); forvar1605 = (forvar1605 + (1'h1)))
        begin
          for (forvar1606 = (1'h0); (forvar1606 < (2'h2)); forvar1606 = (forvar1606 + (1'h1)))
            begin
              reg1607 <= (reg1518[(2'h3):(2'h3)] + (|reg1469));
              reg1608 <= $unsigned({$unsigned($signed(((8'had) ?
                      (8'hbe) : reg1551)))});
              reg1609 = (|(~^{({reg1544, forvar1512} <= ((8'hae) > reg1516))}));
              reg1610 <= reg1548[(3'h4):(2'h2)];
            end
        end
      reg1611 <= (-($unsigned($signed({reg1532, reg1516})) ?
          reg1608 : $unsigned($unsigned(forvar1601[(1'h0):(1'h0)]))));
      reg1612 <= ((^(~&reg1511)) ?
          (8'hb8) : ($unsigned($unsigned({reg1468})) <= forvar1547[(2'h2):(1'h1)]));
    end
  assign wire1613 = $unsigned($signed(((reg1607[(4'hf):(2'h3)] ?
                            {reg1533} : reg1599) ?
                        reg1469 : wire1463[(4'he):(4'ha)])));
  assign wire1614 = $unsigned($unsigned((8'hb1)));
  assign wire1615 = $unsigned((reg1541 >> (~|{$signed(reg1598), wire1462})));
  always
    @(posedge clk) begin
      reg1616 <= ($signed((8'hb1)) ?
          (^(-($signed(reg1469) ?
              ((8'hb3) ^~ reg1551) : (wire1463 ?
                  reg1603 : reg1520)))) : reg1522);
      reg1617 = $unsigned($signed({reg1616[(1'h1):(1'h0)]}));
      reg1618 <= (8'haf);
    end
  assign wire1619 = {reg1604[(4'hc):(1'h0)],
                        {($unsigned($unsigned((7'h40))) ^~ (reg1543 ?
                                forvar1601[(3'h6):(2'h3)] : reg1522[(4'hc):(1'h1)])),
                            (((~&(8'haa)) ?
                                (~^reg1618) : (reg1469 ?
                                    reg1515 : reg1599)) - reg1618)}};
  assign wire1620 = $signed((^reg1616[(2'h3):(1'h0)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1315
#( parameter param1454 = {({{((8'ha8) ? (7'h42) : (8'ha0))}} ? ({((7'h41) ? (8'haa) : (8'hb5))} + ((^(7'h41)) ? ((8'hbb) < (7'h41)) : (8'hb6))) : ((~((8'ha2) ~^ (8'hb4))) >> ((^(8'hb7)) ? (8'hb0) : {(7'h44)}))), (!((((8'hb2) ? (8'ha6) : (8'had)) != {(8'hbe)}) - (((8'hb9) >>> (8'hb8)) ? ((8'hbd) ? (8'hbf) : (7'h40)) : (|(7'h41)))))}
, parameter param1455 = ((8'h9e) || (&({(param1454 >= param1454)} - (param1454 ? (param1454 ? param1454 : param1454) : (param1454 > param1454))))) )
(y, clk, wire1319, wire1318, wire1317, wire1316);
  output wire [(32'h340):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire1319;
  input wire signed [(5'h14):(1'h0)] wire1318;
  input wire signed [(5'h15):(1'h0)] wire1317;
  input wire signed [(4'hf):(1'h0)] wire1316;
  reg [(5'h15):(1'h0)] reg1453 = (1'h0);
  reg [(5'h14):(1'h0)] reg1452 = (1'h0);
  reg [(4'hb):(1'h0)] reg1451 = (1'h0);
  reg [(4'hf):(1'h0)] reg1450 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1449 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1448 = (1'h0);
  reg [(5'h13):(1'h0)] reg1447 = (1'h0);
  reg [(4'hf):(1'h0)] reg1446 = (1'h0);
  reg [(3'h6):(1'h0)] reg1445 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1444 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1443 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1442 = (1'h0);
  reg [(4'hc):(1'h0)] reg1441 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1440 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1439 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1438 = (1'h0);
  reg [(3'h7):(1'h0)] reg1437 = (1'h0);
  reg [(3'h4):(1'h0)] reg1436 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1435 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1434 = (1'h0);
  reg [(3'h7):(1'h0)] reg1433 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1432 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1431 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1430 = (1'h0);
  reg [(4'hf):(1'h0)] reg1429 = (1'h0);
  reg [(5'h14):(1'h0)] reg1428 = (1'h0);
  reg [(5'h14):(1'h0)] reg1427 = (1'h0);
  reg [(4'h8):(1'h0)] reg1426 = (1'h0);
  reg [(3'h7):(1'h0)] reg1425 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1424 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1423 = (1'h0);
  reg [(5'h11):(1'h0)] reg1422 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1421 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1420 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1419 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1418 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire1417;
  wire signed [(5'h12):(1'h0)] wire1346;
  wire signed [(5'h13):(1'h0)] wire1320;
  reg signed [(4'hb):(1'h0)] reg1348 = (1'h0);
  reg [(5'h15):(1'h0)] reg1349 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1350 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1351 = (1'h0);
  reg [(5'h10):(1'h0)] reg1352 = (1'h0);
  reg [(4'hc):(1'h0)] reg1353 = (1'h0);
  reg [(5'h13):(1'h0)] reg1354 = (1'h0);
  reg [(3'h7):(1'h0)] reg1355 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1356 = (1'h0);
  reg [(4'hb):(1'h0)] reg1357 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1358 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1359 = (1'h0);
  reg [(2'h3):(1'h0)] reg1360 = (1'h0);
  reg [(4'he):(1'h0)] reg1361 = (1'h0);
  reg [(4'hc):(1'h0)] reg1362 = (1'h0);
  reg [(2'h2):(1'h0)] reg1363 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1364 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1365 = (1'h0);
  reg [(5'h15):(1'h0)] reg1366 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1367 = (1'h0);
  reg [(5'h15):(1'h0)] reg1368 = (1'h0);
  reg [(4'hc):(1'h0)] reg1369 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1370 = (1'h0);
  reg [(3'h5):(1'h0)] reg1371 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1372 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire1415;
  assign y = {reg1453,
                 reg1452,
                 reg1451,
                 reg1450,
                 reg1449,
                 forvar1448,
                 reg1447,
                 reg1446,
                 reg1445,
                 forvar1444,
                 reg1443,
                 reg1442,
                 reg1441,
                 reg1440,
                 reg1439,
                 forvar1438,
                 reg1437,
                 reg1436,
                 reg1435,
                 forvar1434,
                 reg1433,
                 forvar1432,
                 reg1431,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1427,
                 reg1426,
                 reg1425,
                 reg1424,
                 reg1423,
                 reg1422,
                 reg1421,
                 forvar1420,
                 forvar1419,
                 reg1418,
                 wire1417,
                 wire1346,
                 wire1320,
                 reg1348,
                 reg1349,
                 forvar1350,
                 forvar1351,
                 reg1352,
                 reg1353,
                 reg1354,
                 reg1355,
                 reg1356,
                 reg1357,
                 forvar1358,
                 reg1359,
                 reg1360,
                 reg1361,
                 reg1362,
                 reg1363,
                 reg1364,
                 reg1365,
                 reg1366,
                 reg1367,
                 reg1368,
                 reg1369,
                 reg1370,
                 reg1371,
                 reg1372,
                 wire1415,
                 (1'h0)};
  assign wire1320 = $unsigned($unsigned(wire1317));
  module1321 modinst1347 (.wire1323(wire1319), .wire1322(wire1317), .wire1325(wire1320), .y(wire1346), .wire1324(wire1316), .wire1326(wire1318), .clk(clk));
  always
    @(posedge clk) begin
      reg1348 <= $unsigned($unsigned(wire1319));
      reg1349 <= $unsigned(($signed(({wire1346,
          wire1316} ^ $signed(wire1319))) ^ (((wire1320 ? wire1318 : wire1317) ?
              $unsigned(wire1317) : wire1316) ?
          (~^$signed((7'h40))) : wire1318[(3'h4):(2'h2)])));
      for (forvar1350 = (1'h0); (forvar1350 < (1'h0)); forvar1350 = (forvar1350 + (1'h1)))
        begin
          for (forvar1351 = (1'h0); (forvar1351 < (2'h3)); forvar1351 = (forvar1351 + (1'h1)))
            begin
              reg1352 <= (((~|wire1346[(4'he):(1'h0)]) ^~ wire1316) ?
                  $signed($unsigned($signed((+wire1320)))) : $unsigned((((!reg1348) == forvar1350[(2'h2):(1'h1)]) >= $signed({wire1346}))));
            end
          reg1353 <= (+(8'had));
          reg1354 <= $signed($unsigned((!(~|reg1349))));
          reg1355 <= $signed(wire1316);
          reg1356 = forvar1350[(4'hf):(1'h1)];
        end
      reg1357 = $signed(((wire1320 ? wire1318 : (~$unsigned(wire1320))) ?
          reg1348[(1'h0):(1'h0)] : $signed(reg1355)));
      for (forvar1358 = (1'h0); (forvar1358 < (1'h0)); forvar1358 = (forvar1358 + (1'h1)))
        begin
          reg1359 <= $signed((8'haf));
          reg1360 <= {$signed($unsigned($unsigned((&(8'haf)))))};
          reg1361 <= wire1317;
        end
    end
  always
    @(posedge clk) begin
      reg1362 = (|wire1319);
      reg1363 <= ($signed(($unsigned((reg1355 <<< forvar1350)) ?
              $unsigned($signed((8'hb7))) : $unsigned(((7'h40) ?
                  reg1354 : reg1354)))) ?
          {{(~&{(8'hb9)}), wire1346},
              ($signed({reg1360, reg1349}) ?
                  forvar1350[(4'h9):(1'h1)] : reg1355)} : (&wire1319));
    end
  always
    @(posedge clk) begin
      reg1364 <= (forvar1358[(4'hd):(4'h8)] > ((reg1349 < (~^forvar1350)) ?
          $unsigned(((~|reg1348) ?
              $signed(reg1353) : reg1356)) : ({$unsigned(reg1352),
              (reg1363 << reg1352)} * (~|$signed(wire1346)))));
      reg1365 = ((reg1354 << reg1352[(3'h7):(1'h0)]) ?
          {((8'hb1) ? wire1320[(3'h7):(3'h4)] : $unsigned($signed(reg1354))),
              $signed(((wire1318 ?
                  reg1354 : reg1360) * $signed(wire1346)))} : ((8'hb2) <= $signed({$unsigned(wire1319),
              (forvar1350 < reg1352)})));
      reg1366 <= $unsigned($unsigned((forvar1350 | reg1355)));
    end
  always
    @(posedge clk) begin
      reg1367 <= (~|reg1360);
      reg1368 <= reg1360[(2'h2):(1'h0)];
      reg1369 <= (({(8'hac)} ?
              (!$signed(reg1366[(3'h5):(1'h0)])) : {$unsigned($unsigned(reg1361))}) ?
          ((wire1319 >= reg1349[(2'h3):(1'h1)]) ?
              (~^reg1361) : {$unsigned((~&wire1346))}) : $signed(((+{reg1362,
                  wire1346}) ?
              wire1316 : $unsigned((wire1317 ? wire1317 : reg1364)))));
    end
  always
    @(posedge clk) begin
      reg1370 <= (reg1353[(4'h9):(3'h5)] ^ wire1316);
      reg1371 <= (8'had);
      reg1372 <= (reg1349 ?
          (~^(((~reg1361) ?
              {reg1349, reg1355} : (~|reg1363)) & (reg1356[(5'h15):(4'hd)] ?
              {reg1352} : forvar1358))) : (($signed((reg1356 ?
                      reg1371 : wire1318)) ?
                  $unsigned($signed(forvar1350)) : ({forvar1350} ?
                      {wire1317} : ((8'haf) || reg1367))) ?
              {reg1371} : (reg1365[(4'h8):(1'h1)] <= (~&reg1359))));
    end
  module1373 modinst1416 (wire1415, clk, wire1319, reg1364, reg1353, reg1348, reg1354);
  assign wire1417 = $signed((~($unsigned((reg1371 ?
                        (7'h43) : wire1346)) ^~ reg1348[(2'h2):(1'h0)])));
  always
    @(posedge clk) begin
      reg1418 = (({(^~(!(8'hb9))),
              (!(forvar1358 ? forvar1358 : reg1371))} > reg1369) ?
          $unsigned((($signed(reg1366) ?
              $signed(reg1370) : (reg1348 <<< wire1319)) >= forvar1351)) : (($unsigned(reg1348[(4'ha):(3'h4)]) != (8'hbd)) ?
              reg1365 : ($signed($signed((7'h40))) != {(reg1371 << forvar1350)})));
      for (forvar1419 = (1'h0); (forvar1419 < (1'h0)); forvar1419 = (forvar1419 + (1'h1)))
        begin
          for (forvar1420 = (1'h0); (forvar1420 < (1'h0)); forvar1420 = (forvar1420 + (1'h1)))
            begin
              reg1421 <= wire1417[(3'h4):(3'h4)];
              reg1422 <= $unsigned((^$unsigned($unsigned($unsigned(wire1415)))));
              reg1423 <= (($unsigned(reg1359) ?
                  {(-(wire1417 ^~ reg1418)),
                      reg1367[(1'h1):(1'h0)]} : $signed(($unsigned((8'hb2)) ?
                      $unsigned(reg1356) : $signed(wire1316)))) > (($unsigned((^reg1362)) <= ($signed(reg1422) ?
                  $unsigned(forvar1351) : reg1354[(5'h11):(4'ha)])) >= $signed(($unsigned(reg1370) ?
                  {reg1353} : (~reg1357)))));
              reg1424 <= $unsigned(forvar1420);
              reg1425 <= (^reg1423[(4'hb):(4'h8)]);
            end
          reg1426 = $unsigned($signed(reg1369));
          reg1427 <= ((+$unsigned(reg1369)) ?
              reg1357 : ((reg1354[(2'h3):(2'h2)] <= (~^(reg1359 || reg1356))) ?
                  (8'hb7) : {wire1415[(1'h1):(1'h1)], reg1425[(1'h1):(1'h1)]}));
        end
      reg1428 = $unsigned((forvar1350[(5'h15):(5'h11)] ?
          $unsigned(((reg1418 ~^ (7'h44)) ?
              (reg1364 || reg1349) : reg1360)) : reg1426[(2'h2):(1'h1)]));
    end
  always
    @(posedge clk) begin
      reg1429 <= ($signed((($signed(wire1346) ?
              $unsigned(reg1426) : {wire1320,
                  forvar1358}) > (~&$signed(reg1355)))) ?
          {(reg1368[(5'h13):(4'h8)] ?
                  (reg1428[(3'h6):(3'h4)] >>> (reg1353 == reg1363)) : {(reg1366 | reg1370),
                      reg1370}),
              (|(reg1421 ?
                  $signed(reg1360) : (reg1357 && reg1352)))} : reg1360);
      reg1430 <= (wire1317 && (~forvar1419[(1'h0):(1'h0)]));
      reg1431 <= ((($unsigned((reg1365 ?
              wire1320 : (8'hb2))) <<< (!(reg1352 << reg1354))) ?
          ((~{reg1426}) ?
              wire1316[(4'h8):(1'h1)] : (reg1362[(1'h1):(1'h0)] || (reg1425 ?
                  reg1349 : (8'ha3)))) : wire1316[(4'hd):(4'ha)]) == {reg1424[(1'h0):(1'h0)],
          ((~|$unsigned((8'hb3))) ?
              $signed((!reg1427)) : $unsigned((forvar1420 ?
                  reg1368 : reg1372)))});
      for (forvar1432 = (1'h0); (forvar1432 < (2'h3)); forvar1432 = (forvar1432 + (1'h1)))
        begin
          reg1433 <= $signed(($unsigned(reg1430[(1'h0):(1'h0)]) < {($unsigned(reg1356) ?
                  reg1369[(1'h1):(1'h0)] : (wire1317 ? reg1357 : reg1362)),
              reg1430}));
          for (forvar1434 = (1'h0); (forvar1434 < (3'h4)); forvar1434 = (forvar1434 + (1'h1)))
            begin
              reg1435 <= reg1421;
              reg1436 = (reg1349 ?
                  $signed((~reg1430[(4'h9):(2'h3)])) : (reg1362 ?
                      ({$signed((8'hbe)), (reg1428 ? reg1431 : wire1316)} ?
                          (~|(reg1364 ?
                              (7'h41) : forvar1419)) : reg1369) : reg1364[(4'hd):(4'h8)]));
              reg1437 = $signed($unsigned($unsigned(({reg1359} < ((8'hbc) ?
                  wire1417 : wire1318)))));
            end
          for (forvar1438 = (1'h0); (forvar1438 < (2'h2)); forvar1438 = (forvar1438 + (1'h1)))
            begin
              reg1439 = reg1427[(1'h1):(1'h0)];
              reg1440 = reg1437[(3'h6):(1'h0)];
              reg1441 = (&($unsigned((((7'h40) ?
                  reg1360 : reg1431) ^ $signed(wire1415))) - reg1424));
              reg1442 <= ($signed($signed(wire1415[(1'h0):(1'h0)])) ?
                  $signed(($signed((~^(8'hb5))) ?
                      (reg1437 ?
                          $signed((8'had)) : (reg1367 || reg1371)) : forvar1350[(1'h1):(1'h1)])) : reg1356);
            end
        end
      if (((((~|(reg1422 < reg1359)) ?
          $signed($unsigned(reg1440)) : reg1348[(1'h0):(1'h0)]) ^ $unsigned({(reg1370 < reg1361),
          (reg1425 ? reg1440 : reg1356)})) + reg1366[(2'h2):(1'h1)]))
        begin
          reg1443 <= (!(-{(reg1423 | $signed(reg1441))}));
        end
      else
        begin
          reg1443 = $unsigned(reg1436[(2'h3):(2'h2)]);
          for (forvar1444 = (1'h0); (forvar1444 < (3'h4)); forvar1444 = (forvar1444 + (1'h1)))
            begin
              reg1445 <= (~forvar1351[(4'he):(4'hd)]);
              reg1446 <= (|((($signed(wire1415) ?
                          (reg1435 ? reg1427 : forvar1420) : (reg1422 ?
                              reg1353 : reg1372)) ?
                      reg1431 : reg1360) ?
                  (-(~(8'hb8))) : $unsigned((~$unsigned((8'hbd))))));
              reg1447 = $unsigned({reg1418[(3'h5):(3'h5)],
                  (((+reg1429) >> reg1369) != (+forvar1438))});
            end
          for (forvar1448 = (1'h0); (forvar1448 < (1'h1)); forvar1448 = (forvar1448 + (1'h1)))
            begin
              reg1449 <= $signed($signed($unsigned(((!reg1366) ?
                  (+forvar1448) : wire1317))));
              reg1450 <= $signed($signed(((~^$signed(forvar1350)) ?
                  ((reg1372 << reg1352) * $unsigned(reg1366)) : (forvar1448[(1'h0):(1'h0)] << (wire1318 ?
                      reg1371 : reg1364)))));
              reg1451 <= (((-(~|{reg1363,
                      reg1427})) - (wire1319[(5'h11):(4'ha)] ?
                      $signed(forvar1351[(3'h6):(3'h5)]) : forvar1358[(4'he):(2'h2)])) ?
                  ((^~(!reg1437)) ?
                      $unsigned(((reg1430 | reg1437) ?
                          (wire1320 ? reg1441 : forvar1358) : (reg1449 ?
                              forvar1438 : reg1371))) : $unsigned(reg1424)) : wire1415[(4'hd):(2'h3)]);
              reg1452 = reg1349;
            end
          reg1453 <= reg1368[(3'h7):(1'h1)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1208
#( parameter param1312 = (+((((~(8'haa)) >> (!(8'hb2))) ? (((8'haf) ^ (8'h9f)) == ((8'hbe) >> (7'h43))) : (((7'h44) ? (8'hb5) : (8'hb8)) ? {(8'hb0)} : ((7'h43) <= (8'ha2)))) | (((+(8'hb5)) < ((8'ha8) ? (8'h9c) : (8'hba))) || (|(+(8'hb6)))))) )
(y, clk, wire1213, wire1212, wire1211, wire1210, wire1209);
  output wire [(32'h228):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire1213;
  input wire signed [(3'h4):(1'h0)] wire1212;
  input wire [(2'h3):(1'h0)] wire1211;
  input wire [(5'h12):(1'h0)] wire1210;
  input wire [(4'hb):(1'h0)] wire1209;
  reg signed [(5'h12):(1'h0)] reg1311 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1310 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1309 = (1'h0);
  wire [(3'h4):(1'h0)] wire1308;
  wire signed [(5'h10):(1'h0)] wire1307;
  wire signed [(3'h5):(1'h0)] wire1305;
  reg [(5'h14):(1'h0)] reg1255 = (1'h0);
  reg [(5'h10):(1'h0)] reg1254 = (1'h0);
  reg [(5'h14):(1'h0)] reg1253 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1252 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1251 = (1'h0);
  reg [(2'h2):(1'h0)] reg1250 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1249 = (1'h0);
  wire [(4'hd):(1'h0)] wire1248;
  wire [(5'h11):(1'h0)] wire1247;
  reg [(5'h14):(1'h0)] reg1246 = (1'h0);
  reg [(2'h3):(1'h0)] reg1245 = (1'h0);
  reg [(5'h12):(1'h0)] reg1244 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1243 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire1242;
  wire [(4'he):(1'h0)] wire1241;
  reg [(5'h11):(1'h0)] reg1240 = (1'h0);
  reg [(4'hd):(1'h0)] reg1239 = (1'h0);
  reg [(5'h13):(1'h0)] reg1238 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1237 = (1'h0);
  reg [(5'h12):(1'h0)] reg1236 = (1'h0);
  reg [(3'h6):(1'h0)] reg1235 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1234 = (1'h0);
  reg [(4'he):(1'h0)] reg1233 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1232 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1231 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1230 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1229 = (1'h0);
  reg [(2'h2):(1'h0)] reg1228 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1227 = (1'h0);
  reg [(3'h5):(1'h0)] reg1226 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1225 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1224 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1223 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1222 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1221 = (1'h0);
  reg [(5'h10):(1'h0)] reg1220 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1219 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1218 = (1'h0);
  reg [(4'hf):(1'h0)] reg1217 = (1'h0);
  reg [(4'hd):(1'h0)] reg1216 = (1'h0);
  wire [(3'h7):(1'h0)] wire1215;
  wire signed [(3'h6):(1'h0)] wire1214;
  assign y = {reg1311,
                 reg1310,
                 reg1309,
                 wire1308,
                 wire1307,
                 wire1305,
                 reg1255,
                 reg1254,
                 reg1253,
                 forvar1252,
                 forvar1251,
                 reg1250,
                 reg1249,
                 wire1248,
                 wire1247,
                 reg1246,
                 reg1245,
                 reg1244,
                 reg1243,
                 wire1242,
                 wire1241,
                 reg1240,
                 reg1239,
                 reg1238,
                 reg1237,
                 reg1236,
                 reg1235,
                 reg1234,
                 reg1233,
                 reg1232,
                 forvar1231,
                 forvar1230,
                 reg1229,
                 reg1228,
                 reg1227,
                 reg1226,
                 reg1225,
                 reg1224,
                 forvar1223,
                 forvar1222,
                 reg1221,
                 reg1220,
                 reg1219,
                 reg1218,
                 reg1217,
                 reg1216,
                 wire1215,
                 wire1214,
                 (1'h0)};
  assign wire1214 = wire1211;
  assign wire1215 = ($unsigned($unsigned($unsigned($signed(wire1214)))) || (wire1210[(5'h11):(3'h5)] ?
                        (wire1212 ?
                            wire1212 : wire1214) : $unsigned(($unsigned(wire1211) ?
                            (+wire1212) : $unsigned(wire1211)))));
  always
    @(posedge clk) begin
      reg1216 <= $signed(((8'hbc) ?
          {$signed(wire1211[(1'h0):(1'h0)]),
              (wire1209[(2'h3):(1'h1)] - $unsigned((8'ha8)))} : (8'hbe)));
      reg1217 <= ((wire1215 ? $signed(wire1209) : wire1212[(1'h0):(1'h0)]) ?
          ($signed(({wire1214, wire1211} - wire1213[(2'h2):(1'h0)])) ?
              $unsigned($unsigned((^~wire1213))) : ($unsigned(wire1213) < wire1215)) : $unsigned(wire1213[(3'h4):(2'h2)]));
    end
  always
    @(posedge clk) begin
      reg1218 <= {reg1216[(2'h2):(1'h1)], (^wire1214)};
      reg1219 <= {$unsigned(wire1212[(1'h0):(1'h0)]),
          $signed((reg1217[(3'h7):(1'h1)] ?
              (wire1210[(3'h4):(1'h1)] ?
                  (wire1213 ?
                      wire1215 : wire1215) : (|wire1214)) : ($signed(wire1214) ?
                  $signed(wire1209) : wire1214)))};
    end
  always
    @(posedge clk) begin
      reg1220 <= {((^reg1217[(4'he):(3'h5)]) || $signed(wire1210)), wire1213};
      reg1221 <= ((8'hbe) ? wire1211 : reg1219[(3'h6):(3'h4)]);
      for (forvar1222 = (1'h0); (forvar1222 < (1'h0)); forvar1222 = (forvar1222 + (1'h1)))
        begin
          for (forvar1223 = (1'h0); (forvar1223 < (1'h0)); forvar1223 = (forvar1223 + (1'h1)))
            begin
              reg1224 <= $signed(forvar1223[(1'h0):(1'h0)]);
              reg1225 <= {($unsigned($unsigned((8'ha6))) ?
                      $unsigned((reg1217 >>> $unsigned(wire1213))) : wire1209)};
              reg1226 <= $signed(wire1213[(1'h0):(1'h0)]);
              reg1227 <= ({(|(^$unsigned(reg1220))),
                  $unsigned($signed($unsigned(wire1215)))} >= reg1220);
            end
          reg1228 <= (forvar1222[(3'h4):(1'h1)] ^~ ($unsigned($signed(wire1212[(1'h0):(1'h0)])) ?
              {$unsigned((reg1220 >>> reg1224)),
                  ((~wire1214) ?
                      wire1215 : $signed(reg1219))} : $signed((~^reg1220))));
          reg1229 <= wire1210[(3'h6):(1'h0)];
        end
      for (forvar1230 = (1'h0); (forvar1230 < (2'h3)); forvar1230 = (forvar1230 + (1'h1)))
        begin
          for (forvar1231 = (1'h0); (forvar1231 < (2'h2)); forvar1231 = (forvar1231 + (1'h1)))
            begin
              reg1232 = (8'ha8);
            end
          reg1233 <= (!((reg1226 ?
              ($signed(reg1228) ?
                  $unsigned(reg1227) : ((8'ha7) || reg1229)) : {(reg1220 ?
                      forvar1223 : (8'hac))}) * (reg1216 ?
              {$signed(reg1224), forvar1230} : {(~|(8'hbf)),
                  (wire1213 ^~ wire1211)})));
          if (reg1226[(1'h1):(1'h0)])
            begin
              reg1234 <= reg1220[(4'hb):(2'h2)];
              reg1235 <= ($unsigned(($unsigned(wire1210[(3'h5):(3'h4)]) ?
                  (~|reg1216[(2'h2):(1'h0)]) : $signed((reg1228 ?
                      reg1233 : (8'ha7))))) + reg1228[(1'h1):(1'h1)]);
              reg1236 <= {(wire1209 | (reg1235[(3'h6):(2'h2)] <<< (~^{(8'h9f),
                      reg1228})))};
              reg1237 <= (-reg1227[(3'h4):(2'h3)]);
            end
          else
            begin
              reg1234 = reg1232;
            end
          reg1238 = ((!wire1209[(4'ha):(1'h1)]) ?
              (&(~|$signed((reg1220 ?
                  wire1211 : reg1221)))) : $unsigned((|(+((8'ha6) | (8'ha7))))));
          reg1239 = forvar1222[(2'h2):(2'h2)];
        end
    end
  always
    @(posedge clk) begin
      reg1240 <= {wire1210[(2'h3):(2'h2)]};
    end
  assign wire1241 = ($signed($unsigned({(reg1237 ?
                            wire1214 : reg1237)})) != (~&($signed((7'h42)) - ($signed(wire1213) ?
                        (reg1227 ? forvar1223 : reg1227) : {reg1220}))));
  assign wire1242 = {(reg1238[(3'h4):(1'h1)] - $unsigned((((8'hb9) - reg1234) << $signed(reg1220))))};
  always
    @(posedge clk) begin
      reg1243 <= reg1226;
      reg1244 <= $signed(reg1218[(4'hb):(3'h6)]);
      reg1245 <= ((wire1209[(1'h1):(1'h1)] ?
              wire1212[(2'h2):(1'h0)] : reg1225) ?
          reg1244 : (reg1224[(2'h2):(2'h2)] ?
              wire1211 : $signed($signed(forvar1231[(1'h1):(1'h1)]))));
    end
  always
    @(posedge clk) begin
      reg1246 <= reg1243;
    end
  assign wire1247 = ($unsigned($signed(reg1227[(1'h1):(1'h1)])) ?
                        reg1239[(4'h8):(3'h4)] : $signed($unsigned((((7'h42) ?
                                reg1234 : wire1212) ?
                            (wire1210 ?
                                wire1212 : wire1210) : wire1214[(2'h2):(1'h1)]))));
  assign wire1248 = (((!$signed((-(7'h40)))) <<< ((reg1244 ^ $unsigned(forvar1223)) ^~ ({reg1237,
                            (7'h40)} || $unsigned(forvar1231)))) ?
                        $unsigned($unsigned(reg1233)) : ({(~|(reg1218 ?
                                forvar1223 : wire1215)),
                            wire1213} && reg1232));
  always
    @(posedge clk) begin
      reg1249 <= (($unsigned(reg1221) ^~ wire1209) - ($signed($signed((wire1211 ?
          (8'h9d) : reg1220))) <= $signed(wire1215[(1'h1):(1'h0)])));
      reg1250 <= forvar1222;
      for (forvar1251 = (1'h0); (forvar1251 < (1'h0)); forvar1251 = (forvar1251 + (1'h1)))
        begin
          for (forvar1252 = (1'h0); (forvar1252 < (1'h1)); forvar1252 = (forvar1252 + (1'h1)))
            begin
              reg1253 = reg1234[(4'hc):(2'h3)];
            end
        end
      reg1254 = ((8'hb3) ?
          (~wire1247[(3'h4):(1'h1)]) : (reg1227 != ($unsigned((~|wire1248)) != ($unsigned(wire1214) ?
              $unsigned(reg1234) : reg1217[(4'hd):(1'h1)]))));
      reg1255 <= $signed($unsigned({wire1242,
          ((reg1227 >= forvar1251) + reg1225)}));
    end
  module1256 modinst1306 (wire1305, clk, reg1220, forvar1231, wire1210, reg1246);
  assign wire1307 = {$unsigned({$signed($signed(forvar1222))}),
                        (wire1209 ?
                            (~^reg1240[(2'h2):(1'h1)]) : ($signed(wire1215[(3'h7):(2'h3)]) == $signed(reg1233)))};
  assign wire1308 = (8'ha8);
  always
    @(posedge clk) begin
      reg1309 = $signed((~(8'ha4)));
      reg1310 <= $unsigned($signed($unsigned($signed(wire1241[(2'h2):(1'h0)]))));
      reg1311 <= wire1305;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1256
#( parameter param1304 = ((~|(~|{((8'hb5) ^~ (8'ha4)), ((8'hb5) ? (8'ha0) : (8'haf))})) ~^ (((8'hb0) || ({(8'hb3), (8'hb1)} != ((8'hbf) & (8'ha2)))) <= (~&(8'hbb)))) )
(y, clk, wire1260, wire1259, wire1258, wire1257);
  output wire [(32'h1dd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire1260;
  input wire [(5'h12):(1'h0)] wire1259;
  input wire signed [(5'h10):(1'h0)] wire1258;
  input wire [(5'h14):(1'h0)] wire1257;
  wire signed [(5'h10):(1'h0)] wire1303;
  wire signed [(5'h12):(1'h0)] wire1302;
  wire signed [(4'h8):(1'h0)] wire1301;
  wire [(4'hd):(1'h0)] wire1300;
  reg [(5'h13):(1'h0)] reg1299 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1298 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1297 = (1'h0);
  reg [(4'hf):(1'h0)] reg1296 = (1'h0);
  reg [(5'h13):(1'h0)] reg1295 = (1'h0);
  reg [(2'h2):(1'h0)] reg1294 = (1'h0);
  reg [(2'h2):(1'h0)] reg1293 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1292 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1291 = (1'h0);
  reg [(3'h4):(1'h0)] reg1290 = (1'h0);
  reg [(5'h13):(1'h0)] reg1289 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1288 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1287 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1286 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire1285;
  wire [(5'h14):(1'h0)] wire1284;
  wire signed [(5'h14):(1'h0)] wire1283;
  wire signed [(3'h4):(1'h0)] wire1282;
  reg signed [(4'hc):(1'h0)] reg1281 = (1'h0);
  reg [(3'h7):(1'h0)] reg1280 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1279 = (1'h0);
  reg [(3'h6):(1'h0)] reg1278 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1277 = (1'h0);
  reg [(5'h13):(1'h0)] reg1276 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1275 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1274 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1273 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1272 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1271 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1270 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1269 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1268 = (1'h0);
  reg [(2'h3):(1'h0)] reg1267 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1266 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1265 = (1'h0);
  reg [(4'h9):(1'h0)] reg1264 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1263 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire1262;
  wire [(3'h7):(1'h0)] wire1261;
  assign y = {wire1303,
                 wire1302,
                 wire1301,
                 wire1300,
                 reg1299,
                 forvar1298,
                 reg1297,
                 reg1296,
                 reg1295,
                 reg1294,
                 reg1293,
                 reg1292,
                 reg1291,
                 reg1290,
                 reg1289,
                 reg1288,
                 forvar1287,
                 forvar1286,
                 wire1285,
                 wire1284,
                 wire1283,
                 wire1282,
                 reg1281,
                 reg1280,
                 forvar1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 forvar1275,
                 reg1274,
                 reg1273,
                 reg1272,
                 reg1271,
                 forvar1270,
                 reg1269,
                 reg1268,
                 reg1267,
                 reg1266,
                 reg1265,
                 reg1264,
                 reg1263,
                 wire1262,
                 wire1261,
                 (1'h0)};
  assign wire1261 = ($unsigned($signed((wire1257 ?
                        wire1258 : (|wire1260)))) & $unsigned((((8'hbf) >>> (wire1258 ?
                            wire1259 : wire1257)) ?
                        $unsigned($unsigned(wire1260)) : (~&$signed(wire1260)))));
  assign wire1262 = (~((8'hb8) ?
                        (^~wire1258) : (wire1257[(4'h8):(3'h6)] & (-(wire1258 ?
                            wire1259 : wire1258)))));
  always
    @(posedge clk) begin
      reg1263 <= wire1257;
      reg1264 = $unsigned(($unsigned($unsigned(wire1260[(3'h7):(3'h5)])) < (wire1257[(2'h3):(2'h2)] ?
          (wire1260[(3'h6):(3'h6)] ?
              (wire1262 <= wire1262) : {(8'haa)}) : (((8'hbd) | wire1259) * (wire1262 ?
              wire1260 : wire1259)))));
      reg1265 <= ($signed((($signed(wire1258) >> wire1261[(2'h2):(1'h1)]) * {{wire1257},
              (reg1264 & (8'h9f))})) ?
          (((wire1257[(3'h5):(1'h0)] * (reg1264 + wire1262)) != wire1257[(4'h8):(3'h5)]) != (reg1263[(2'h2):(1'h1)] ?
              $signed((wire1258 ?
                  reg1263 : wire1257)) : $unsigned(((8'hb2) - wire1261)))) : (|wire1260[(3'h4):(2'h3)]));
      reg1266 <= ($signed(((~|(wire1260 < wire1261)) & $unsigned($signed(wire1258)))) >>> (wire1259 | (8'hbb)));
      reg1267 = (~|(~&$unsigned($unsigned((wire1261 ? wire1261 : reg1263)))));
    end
  always
    @(posedge clk) begin
      reg1268 = reg1265;
      reg1269 = (wire1258[(4'ha):(3'h6)] ?
          wire1259[(4'hb):(4'hb)] : {$unsigned($unsigned((reg1268 ?
                  wire1261 : reg1268))),
              wire1261[(3'h7):(1'h0)]});
      for (forvar1270 = (1'h0); (forvar1270 < (1'h0)); forvar1270 = (forvar1270 + (1'h1)))
        begin
          reg1271 <= (({reg1264[(4'h8):(3'h6)],
                      {(~&wire1261), $signed(reg1266)}} ?
                  $unsigned((reg1263[(2'h3):(1'h0)] > $unsigned(reg1267))) : (&wire1259)) ?
              wire1259[(1'h0):(1'h0)] : (!($unsigned(reg1263) < $unsigned(wire1257))));
          reg1272 = reg1271[(4'h9):(3'h5)];
          reg1273 <= wire1257;
          reg1274 <= (~|(&($signed({wire1257,
              (8'hb6)}) == {reg1265[(3'h4):(1'h1)], $unsigned(reg1269)})));
        end
      for (forvar1275 = (1'h0); (forvar1275 < (1'h0)); forvar1275 = (forvar1275 + (1'h1)))
        begin
          reg1276 <= ($signed(reg1263) ? reg1272[(4'h8):(4'h8)] : forvar1270);
          reg1277 <= reg1273;
          reg1278 <= ((~|$unsigned($signed(wire1257[(3'h5):(2'h2)]))) <<< ((reg1265[(3'h5):(3'h4)] ?
                  $unsigned(reg1265[(3'h4):(3'h4)]) : ((~&reg1267) ?
                      (reg1264 != wire1260) : reg1265)) ?
              ($unsigned($unsigned((7'h41))) <<< ((reg1272 ?
                  reg1277 : reg1274) != $unsigned(reg1274))) : $unsigned({(reg1267 && reg1264),
                  (!forvar1270)})));
        end
    end
  always
    @(posedge clk) begin
      for (forvar1279 = (1'h0); (forvar1279 < (2'h2)); forvar1279 = (forvar1279 + (1'h1)))
        begin
          reg1280 <= $signed({reg1273[(1'h1):(1'h1)], $unsigned(forvar1279)});
          reg1281 = $signed((reg1272[(2'h2):(1'h0)] ?
              $unsigned((~$signed(reg1264))) : wire1262[(1'h1):(1'h1)]));
        end
    end
  assign wire1282 = {((((reg1276 ? reg1278 : forvar1275) ?
                                    ((8'hab) - reg1271) : wire1262) ?
                                ($signed((8'hac)) || (reg1281 ?
                                    forvar1275 : (8'ha0))) : (wire1259 ?
                                    reg1264[(1'h0):(1'h0)] : wire1262[(1'h1):(1'h1)])) ?
                            $signed($signed(wire1258[(5'h10):(4'ha)])) : ((reg1281[(1'h1):(1'h1)] & (&reg1278)) >>> (wire1258[(4'ha):(4'h8)] + (^(8'ha8)))))};
  assign wire1283 = forvar1270;
  assign wire1284 = $unsigned((-$unsigned((~(~|wire1258)))));
  assign wire1285 = (((~|$unsigned(wire1262[(1'h1):(1'h0)])) ?
                        reg1277 : reg1263[(3'h4):(1'h1)]) >> (~|(8'ha6)));
  always
    @(posedge clk) begin
      for (forvar1286 = (1'h0); (forvar1286 < (1'h0)); forvar1286 = (forvar1286 + (1'h1)))
        begin
          for (forvar1287 = (1'h0); (forvar1287 < (1'h1)); forvar1287 = (forvar1287 + (1'h1)))
            begin
              reg1288 <= wire1283[(5'h13):(3'h7)];
              reg1289 = (~&$signed({(~|reg1266),
                  ($signed(wire1260) ?
                      reg1264[(2'h2):(1'h0)] : $signed(reg1265))}));
              reg1290 <= wire1285[(3'h5):(2'h3)];
              reg1291 <= wire1258;
              reg1292 = ($unsigned(($signed(wire1283) && ((reg1281 ^ (8'hb4)) ?
                  {reg1269} : $signed(reg1291)))) <<< $signed((|{(wire1282 && reg1280),
                  (~^reg1277)})));
            end
          reg1293 <= reg1268;
          reg1294 = $unsigned(((~$signed((!reg1264))) | ((wire1261 & $signed(wire1284)) ?
              (wire1261 > (~reg1276)) : wire1262[(1'h0):(1'h0)])));
          reg1295 <= (8'ha4);
        end
      reg1296 <= (^(~&$signed(((-wire1262) - wire1284))));
      reg1297 <= reg1273[(2'h2):(1'h0)];
      for (forvar1298 = (1'h0); (forvar1298 < (1'h0)); forvar1298 = (forvar1298 + (1'h1)))
        begin
          reg1299 <= (forvar1298[(1'h0):(1'h0)] - (((&(|reg1297)) ?
                  wire1262 : $unsigned($unsigned((8'ha0)))) ?
              ($signed($signed(reg1273)) >>> {reg1295[(3'h6):(3'h5)]}) : reg1271[(1'h1):(1'h0)]));
        end
    end
  assign wire1300 = reg1296;
  assign wire1301 = reg1289;
  assign wire1302 = reg1281;
  assign wire1303 = ($unsigned($signed((7'h41))) ^~ ($unsigned(((reg1271 ?
                                forvar1279 : reg1274) ?
                            reg1293 : reg1267[(2'h3):(1'h0)])) ?
                        $unsigned($signed(forvar1270[(3'h6):(1'h1)])) : (reg1281 ?
                            $unsigned((~&reg1280)) : ((!reg1297) || wire1259))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1373
#( parameter param1414 = (~^(((~{(8'hb4)}) ? (((7'h41) ^~ (8'hb5)) ? ((8'ha0) ? (8'ha1) : (8'hbd)) : {(8'ha3), (7'h40)}) : ((-(8'hb7)) ? ((8'hbe) ? (8'hb9) : (8'ha7)) : ((8'hae) + (8'hbc)))) ? {(~((8'hb0) * (8'ha4)))} : ((-(|(7'h42))) ? (^~((8'h9f) ? (8'hb8) : (8'ha9))) : {((8'h9e) > (8'hb5))}))) )
(y, clk, wire1378, wire1377, wire1376, wire1375, wire1374);
  output wire [(32'h1ab):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire1378;
  input wire signed [(5'h14):(1'h0)] wire1377;
  input wire signed [(4'hc):(1'h0)] wire1376;
  input wire signed [(2'h3):(1'h0)] wire1375;
  input wire [(5'h13):(1'h0)] wire1374;
  wire [(5'h13):(1'h0)] wire1413;
  reg signed [(5'h11):(1'h0)] reg1412 = (1'h0);
  reg [(4'h8):(1'h0)] reg1411 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1410 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1409 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1408 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1407 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1406 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1405 = (1'h0);
  reg [(5'h14):(1'h0)] reg1404 = (1'h0);
  reg [(5'h10):(1'h0)] reg1403 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1402 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1401 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1400 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1399 = (1'h0);
  wire [(3'h6):(1'h0)] wire1398;
  wire [(5'h10):(1'h0)] wire1397;
  reg signed [(2'h3):(1'h0)] reg1396 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1395 = (1'h0);
  reg [(5'h10):(1'h0)] reg1394 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1393 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire1392;
  reg signed [(3'h4):(1'h0)] reg1391 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1390 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1389 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1388 = (1'h0);
  reg [(4'hc):(1'h0)] reg1387 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1386 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1383 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1385 = (1'h0);
  reg [(3'h7):(1'h0)] reg1384 = (1'h0);
  reg [(4'hb):(1'h0)] reg1383 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1382 = (1'h0);
  reg [(5'h12):(1'h0)] reg1381 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1380 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire1379;
  assign y = {wire1413,
                 reg1412,
                 reg1411,
                 forvar1410,
                 forvar1409,
                 reg1408,
                 reg1407,
                 forvar1406,
                 reg1405,
                 reg1404,
                 reg1403,
                 reg1402,
                 reg1401,
                 reg1400,
                 reg1399,
                 wire1398,
                 wire1397,
                 reg1396,
                 reg1395,
                 reg1394,
                 reg1393,
                 wire1392,
                 reg1391,
                 reg1390,
                 reg1389,
                 reg1388,
                 reg1387,
                 reg1386,
                 forvar1383,
                 reg1385,
                 reg1384,
                 reg1383,
                 reg1382,
                 reg1381,
                 reg1380,
                 wire1379,
                 (1'h0)};
  assign wire1379 = ($signed((wire1376 << wire1374[(4'hd):(4'h9)])) > (wire1375[(2'h3):(2'h3)] ~^ ({wire1378,
                            (8'ha3)} ?
                        wire1376 : (^~$unsigned(wire1375)))));
  always
    @(posedge clk) begin
      reg1380 <= ((wire1374[(4'hd):(4'h8)] >= ((&wire1375[(1'h1):(1'h1)]) ?
              (+((8'haf) ? wire1378 : wire1376)) : (wire1374[(4'h9):(3'h5)] ?
                  wire1375 : wire1378[(3'h6):(3'h6)]))) ?
          $unsigned(wire1374) : ((~wire1375) ?
              {(wire1376[(2'h2):(2'h2)] ?
                      {wire1378} : ((8'haa) ?
                          wire1379 : wire1376))} : wire1378));
      reg1381 <= ($signed((-$unsigned(((8'ha1) != wire1376)))) * {$unsigned($unsigned($unsigned(reg1380)))});
      reg1382 <= $unsigned((wire1376 ?
          $signed($unsigned((wire1376 | (8'ha6)))) : $unsigned((-reg1381))));
      if ((wire1376 ?
          reg1382 : {(wire1374[(5'h12):(4'ha)] ?
                  wire1379 : wire1377[(4'ha):(3'h4)]),
              reg1382[(3'h5):(1'h1)]}))
        begin
          reg1383 <= $signed($unsigned((((wire1379 <<< wire1377) ?
              reg1381 : wire1374) <<< ((&wire1376) & (wire1378 ~^ wire1377)))));
          reg1384 <= ($unsigned($unsigned(wire1376[(2'h3):(1'h0)])) ?
              (+wire1376) : wire1378[(2'h3):(2'h2)]);
          reg1385 = ((8'ha3) | wire1374[(3'h4):(2'h2)]);
        end
      else
        begin
          for (forvar1383 = (1'h0); (forvar1383 < (1'h0)); forvar1383 = (forvar1383 + (1'h1)))
            begin
              reg1384 <= reg1382;
              reg1385 <= $unsigned(forvar1383[(2'h3):(1'h0)]);
            end
          reg1386 <= wire1377[(4'h9):(3'h4)];
          reg1387 = $unsigned($unsigned($signed(reg1383)));
          reg1388 <= wire1376;
          reg1389 = $unsigned((8'hbf));
        end
      reg1390 <= ($unsigned(reg1385[(4'hf):(4'he)]) ?
          $signed($unsigned((~(wire1379 ?
              (7'h44) : reg1383)))) : {wire1379[(3'h6):(2'h2)]});
    end
  always
    @(posedge clk) begin
      reg1391 <= $unsigned($unsigned(reg1385));
    end
  assign wire1392 = reg1386[(3'h6):(2'h2)];
  always
    @(posedge clk) begin
      reg1393 = $unsigned(wire1376);
      reg1394 <= wire1379[(2'h3):(2'h3)];
      reg1395 <= (~$unsigned($unsigned({$unsigned(reg1390),
          $signed(reg1382)})));
      reg1396 = reg1387[(3'h5):(1'h1)];
    end
  assign wire1397 = reg1384[(3'h4):(2'h2)];
  assign wire1398 = $unsigned(((($signed(wire1397) > $unsigned(wire1379)) ^ (~$unsigned(reg1389))) ?
                        wire1397 : $unsigned(wire1377)));
  always
    @(posedge clk) begin
      reg1399 <= reg1389;
    end
  always
    @(posedge clk) begin
      reg1400 <= $signed(reg1385[(5'h11):(5'h11)]);
      reg1401 <= ($unsigned(wire1374[(4'h9):(3'h4)]) <= ($signed($signed(reg1396[(1'h0):(1'h0)])) ?
          (~|{{reg1388}, $unsigned((8'ha7))}) : $signed((+reg1385))));
      reg1402 <= {(($unsigned((-wire1398)) ?
              $signed($signed(reg1381)) : (-(reg1394 ?
                  reg1391 : reg1399))) + $signed($unsigned((wire1374 ?
              reg1401 : reg1380)))),
          $unsigned(((~$signed((7'h40))) >>> ($signed(reg1396) || (~reg1388))))};
      reg1403 <= wire1375[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg1404 <= ($signed((($unsigned(reg1391) ?
          wire1374[(2'h2):(1'h1)] : $signed(reg1391)) >> reg1389[(1'h0):(1'h0)])) >= ((reg1389[(4'ha):(3'h4)] >> wire1378[(4'he):(2'h2)]) ?
          reg1384 : reg1393[(4'ha):(1'h0)]));
      reg1405 <= ($unsigned(wire1379) ?
          ((~&reg1380) ?
              ($unsigned(reg1403) >= $unsigned(reg1386[(1'h1):(1'h0)])) : reg1393[(4'hf):(3'h5)]) : (8'haf));
      for (forvar1406 = (1'h0); (forvar1406 < (1'h1)); forvar1406 = (forvar1406 + (1'h1)))
        begin
          reg1407 <= $signed((reg1393 * (((-reg1401) << $signed(reg1395)) ?
              ((^(8'ha7)) ?
                  (&wire1379) : reg1400[(3'h5):(1'h1)]) : ((reg1400 >> reg1386) && ((8'h9f) ?
                  reg1401 : reg1389)))));
          reg1408 = reg1405;
        end
      for (forvar1409 = (1'h0); (forvar1409 < (1'h1)); forvar1409 = (forvar1409 + (1'h1)))
        begin
          for (forvar1410 = (1'h0); (forvar1410 < (1'h1)); forvar1410 = (forvar1410 + (1'h1)))
            begin
              reg1411 <= (~&((!{$signed(reg1386),
                  ((8'ha9) ?
                      reg1405 : (8'hbb))}) <= $unsigned($signed((~&reg1395)))));
            end
          reg1412 <= (^(reg1396 ?
              (8'h9c) : (($unsigned(reg1386) ^ $unsigned(reg1383)) - (8'ha4))));
        end
    end
  assign wire1413 = reg1393;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1321
#( parameter param1345 = {((&(((8'h9e) ? (8'ha7) : (8'haf)) ? ((8'ha6) ? (8'ha3) : (8'hbd)) : ((8'hbd) >>> (8'hbe)))) >= ((8'hb0) <= {(-(8'hbc)), ((8'hb0) ? (7'h44) : (8'h9e))})), (((^{(8'hbc)}) ? {(|(8'ha3))} : ((7'h40) ^~ ((8'hb3) ? (8'hbe) : (8'hab)))) && (~|(!((8'hae) << (8'hb5)))))} )
(y, clk, wire1326, wire1325, wire1324, wire1323, wire1322);
  output wire [(32'hd7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire1326;
  input wire signed [(2'h2):(1'h0)] wire1325;
  input wire signed [(4'hf):(1'h0)] wire1324;
  input wire signed [(3'h6):(1'h0)] wire1323;
  input wire signed [(4'h8):(1'h0)] wire1322;
  reg [(3'h7):(1'h0)] forvar1341 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1338 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1337 = (1'h0);
  reg [(4'h8):(1'h0)] reg1344 = (1'h0);
  reg [(4'h9):(1'h0)] reg1343 = (1'h0);
  reg [(4'hf):(1'h0)] reg1342 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1341 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1340 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1339 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1338 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1337 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire1336;
  wire signed [(4'h8):(1'h0)] wire1335;
  reg signed [(4'hf):(1'h0)] reg1334 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1333 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire1332;
  reg [(4'he):(1'h0)] reg1331 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1330 = (1'h0);
  reg [(3'h5):(1'h0)] reg1329 = (1'h0);
  wire [(4'ha):(1'h0)] wire1328;
  wire [(4'ha):(1'h0)] wire1327;
  assign y = {forvar1341,
                 reg1338,
                 forvar1337,
                 reg1344,
                 reg1343,
                 reg1342,
                 reg1341,
                 reg1340,
                 reg1339,
                 forvar1338,
                 reg1337,
                 wire1336,
                 wire1335,
                 reg1334,
                 reg1333,
                 wire1332,
                 reg1331,
                 reg1330,
                 reg1329,
                 wire1328,
                 wire1327,
                 (1'h0)};
  assign wire1327 = $unsigned((!(-$unsigned(wire1322[(1'h0):(1'h0)]))));
  assign wire1328 = (-wire1322);
  always
    @(posedge clk) begin
      reg1329 <= $signed(wire1327);
      reg1330 <= ((wire1328 + (($unsigned((8'hbe)) ?
              (|wire1325) : $signed(wire1328)) > (~|$unsigned((8'hbb))))) ?
          $signed((-wire1323[(2'h3):(2'h3)])) : (wire1324[(3'h4):(2'h3)] | wire1328));
      reg1331 <= $signed(reg1329[(2'h2):(1'h0)]);
    end
  assign wire1332 = wire1325[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg1333 <= {(8'hb1), $unsigned({$signed($signed((8'ha7))), wire1327})};
      reg1334 <= {($unsigned($signed($unsigned(wire1328))) < (wire1327[(3'h4):(2'h2)] >> $signed((reg1333 && wire1324))))};
    end
  assign wire1335 = wire1323[(3'h6):(3'h5)];
  assign wire1336 = (reg1329 ?
                        ($unsigned(wire1335[(1'h1):(1'h0)]) ?
                            (reg1331 + $signed($unsigned(reg1333))) : reg1334) : wire1322[(3'h6):(3'h5)]);
  always
    @(posedge clk) begin
      if ($unsigned(($signed(((wire1323 ? wire1328 : reg1331) ?
          $signed(reg1330) : (wire1324 ? reg1333 : wire1324))) - ((8'h9e) ?
          reg1330[(3'h4):(1'h0)] : $signed(reg1333)))))
        begin
          reg1337 <= (reg1329[(2'h3):(1'h0)] <= reg1333);
          for (forvar1338 = (1'h0); (forvar1338 < (2'h2)); forvar1338 = (forvar1338 + (1'h1)))
            begin
              reg1339 = wire1328;
              reg1340 <= $unsigned(($unsigned(($signed(reg1331) & (wire1326 ?
                  (8'had) : (8'haf)))) | ($signed(reg1334[(4'h8):(1'h1)]) ?
                  wire1322 : wire1324[(3'h5):(1'h1)])));
              reg1341 <= wire1324;
            end
          reg1342 <= forvar1338;
          reg1343 <= {(~&$signed($signed((wire1327 ? wire1326 : reg1339)))),
              $signed(wire1326)};
          reg1344 <= wire1323[(3'h4):(2'h2)];
        end
      else
        begin
          for (forvar1337 = (1'h0); (forvar1337 < (2'h2)); forvar1337 = (forvar1337 + (1'h1)))
            begin
              reg1338 <= ({($signed((reg1343 <= reg1330)) != reg1331[(2'h3):(1'h1)]),
                      $signed((wire1322 || {(8'hb4)}))} ?
                  ({(^((8'hb2) && reg1342))} != (~(wire1327 + (wire1326 <<< forvar1338)))) : wire1325);
              reg1339 <= $unsigned((^$unsigned(reg1341)));
              reg1340 = $signed(reg1333);
            end
          for (forvar1341 = (1'h0); (forvar1341 < (3'h4)); forvar1341 = (forvar1341 + (1'h1)))
            begin
              reg1342 = $unsigned(reg1338[(4'h9):(3'h4)]);
              reg1343 <= reg1330;
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1552
#( parameter param1595 = (~(&((^(^~(8'ha6))) ? (((8'ha9) > (8'hba)) ? ((8'ha4) ? (8'ha0) : (8'hb7)) : ((8'h9d) && (8'hac))) : (((8'hab) ? (8'ha7) : (8'haf)) || (~^(8'had)))))) )
(y, clk, wire1556, wire1555, wire1554, wire1553);
  output wire [(32'h17b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire1556;
  input wire signed [(5'h14):(1'h0)] wire1555;
  input wire signed [(5'h14):(1'h0)] wire1554;
  input wire signed [(4'ha):(1'h0)] wire1553;
  reg [(4'hd):(1'h0)] reg1594 = (1'h0);
  wire signed [(4'he):(1'h0)] wire1593;
  wire signed [(5'h12):(1'h0)] wire1592;
  reg [(5'h13):(1'h0)] reg1591 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1590 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1589 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1588 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1587 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1586 = (1'h0);
  reg [(4'hb):(1'h0)] reg1585 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1584 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1583 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1582 = (1'h0);
  reg [(2'h3):(1'h0)] reg1581 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1580 = (1'h0);
  reg [(2'h3):(1'h0)] reg1579 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1578 = (1'h0);
  reg [(3'h4):(1'h0)] reg1577 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1576 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1575 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1574 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1573 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1572 = (1'h0);
  reg [(4'hb):(1'h0)] reg1571 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire1570;
  reg signed [(3'h6):(1'h0)] reg1569 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1568 = (1'h0);
  reg [(4'hf):(1'h0)] reg1567 = (1'h0);
  reg [(4'hd):(1'h0)] reg1566 = (1'h0);
  reg [(4'hd):(1'h0)] reg1565 = (1'h0);
  reg [(5'h13):(1'h0)] reg1564 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1563 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1562 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1561 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1560 = (1'h0);
  reg [(3'h4):(1'h0)] reg1559 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1558 = (1'h0);
  reg [(4'hd):(1'h0)] reg1557 = (1'h0);
  assign y = {reg1594,
                 wire1593,
                 wire1592,
                 reg1591,
                 reg1590,
                 reg1589,
                 reg1588,
                 reg1587,
                 reg1586,
                 reg1585,
                 reg1584,
                 reg1583,
                 reg1582,
                 reg1581,
                 forvar1580,
                 reg1579,
                 reg1578,
                 reg1577,
                 reg1576,
                 reg1575,
                 forvar1574,
                 reg1573,
                 forvar1572,
                 reg1571,
                 wire1570,
                 reg1569,
                 reg1568,
                 reg1567,
                 reg1566,
                 reg1565,
                 reg1564,
                 reg1563,
                 reg1562,
                 reg1561,
                 forvar1560,
                 reg1559,
                 forvar1558,
                 reg1557,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1557 = wire1553;
      for (forvar1558 = (1'h0); (forvar1558 < (1'h0)); forvar1558 = (forvar1558 + (1'h1)))
        begin
          reg1559 <= wire1553;
          for (forvar1560 = (1'h0); (forvar1560 < (3'h4)); forvar1560 = (forvar1560 + (1'h1)))
            begin
              reg1561 <= $signed((!$signed({wire1555[(5'h13):(1'h0)]})));
              reg1562 <= $signed(forvar1558[(3'h7):(3'h4)]);
              reg1563 <= (((!reg1562) + ($unsigned($unsigned(wire1553)) << reg1559)) ?
                  {$signed(wire1555)} : wire1553[(2'h2):(1'h0)]);
              reg1564 <= {$unsigned(reg1563[(2'h2):(1'h0)])};
              reg1565 <= ($unsigned((($unsigned(reg1557) || $signed(reg1562)) ?
                      {forvar1558} : $unsigned(reg1561))) ?
                  (~{({wire1555} ~^ wire1556[(4'hc):(4'h8)])}) : $unsigned((($unsigned(reg1562) & (reg1559 | reg1563)) ?
                      (forvar1558 ^~ {wire1553}) : (!wire1553[(3'h5):(2'h2)]))));
            end
          reg1566 <= ((7'h41) ?
              reg1563[(1'h1):(1'h1)] : (($signed(reg1562[(1'h1):(1'h1)]) ?
                  wire1554[(5'h13):(2'h3)] : (8'hab)) > ($signed(reg1563[(2'h2):(1'h0)]) && $signed(reg1563))));
        end
      reg1567 = {(wire1555[(4'hc):(3'h6)] ?
              (((~&reg1561) ? $unsigned(wire1555) : (-wire1555)) ?
                  (^~$signed(wire1555)) : reg1561) : (^~reg1563[(3'h4):(3'h4)]))};
      reg1568 = $signed($unsigned($signed(({reg1561,
          reg1562} ^ $unsigned(reg1566)))));
      reg1569 = $unsigned(((~wire1554[(2'h3):(1'h0)]) < wire1553));
    end
  assign wire1570 = reg1559;
  always
    @(posedge clk) begin
      reg1571 <= (+$signed((~(~^$unsigned(wire1556)))));
      for (forvar1572 = (1'h0); (forvar1572 < (2'h2)); forvar1572 = (forvar1572 + (1'h1)))
        begin
          reg1573 <= $unsigned($unsigned({{$signed((8'ha7))},
              {(reg1561 + (8'hb8)), (^~reg1568)}}));
          for (forvar1574 = (1'h0); (forvar1574 < (2'h3)); forvar1574 = (forvar1574 + (1'h1)))
            begin
              reg1575 <= reg1565[(3'h6):(1'h0)];
              reg1576 <= ($unsigned((~^((+reg1561) ?
                  reg1564[(4'hd):(4'hd)] : reg1565))) | reg1575);
              reg1577 <= reg1569[(3'h5):(3'h4)];
            end
          reg1578 = (-$signed((+{$signed(reg1568)})));
        end
    end
  always
    @(posedge clk) begin
      reg1579 <= $unsigned(reg1563);
      for (forvar1580 = (1'h0); (forvar1580 < (3'h4)); forvar1580 = (forvar1580 + (1'h1)))
        begin
          reg1581 = $signed((7'h40));
          reg1582 <= (~&((({reg1566, reg1569} ?
                  (|forvar1558) : $signed(forvar1580)) ?
              forvar1560[(4'hb):(3'h5)] : forvar1558[(4'ha):(1'h0)]) * (!forvar1574[(2'h3):(1'h0)])));
          reg1583 <= $unsigned($signed(($signed($unsigned(wire1554)) ~^ reg1565[(4'ha):(4'h8)])));
        end
      reg1584 <= (forvar1572 ? forvar1558 : (|forvar1574));
    end
  always
    @(posedge clk) begin
      reg1585 <= $signed($unsigned((wire1555[(1'h1):(1'h0)] > (~reg1569[(1'h0):(1'h0)]))));
      reg1586 = (8'had);
    end
  always
    @(posedge clk) begin
      reg1587 <= reg1578;
      reg1588 <= $signed($signed({((reg1577 <<< reg1569) | reg1563)}));
      reg1589 <= $signed({$unsigned(reg1576), reg1569[(1'h1):(1'h0)]});
    end
  always
    @(posedge clk) begin
      reg1590 <= ((forvar1560 ~^ $signed((wire1554 < $unsigned(forvar1580)))) ?
          (!$signed($signed($unsigned(forvar1572)))) : $signed(({(reg1565 ?
                  forvar1574 : reg1583),
              $unsigned(reg1587)} || reg1582)));
      reg1591 <= $unsigned(reg1583);
    end
  assign wire1592 = (!$signed(reg1582[(3'h4):(2'h3)]));
  assign wire1593 = ((^~reg1561[(2'h2):(2'h2)]) ?
                        wire1555[(4'ha):(3'h5)] : reg1561);
  always
    @(posedge clk) begin
      reg1594 = $unsigned(((-reg1582[(3'h4):(3'h4)]) * $unsigned(reg1581)));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1472  (y, clk, wire1476, wire1475, wire1474, wire1473);
  output wire [(32'h170):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire1476;
  input wire signed [(3'h7):(1'h0)] wire1475;
  input wire [(5'h12):(1'h0)] wire1474;
  input wire [(5'h14):(1'h0)] wire1473;
  wire signed [(2'h3):(1'h0)] wire1507;
  reg [(5'h14):(1'h0)] reg1506 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1505 = (1'h0);
  reg [(5'h12):(1'h0)] reg1504 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1503;
  reg [(4'h9):(1'h0)] reg1502 = (1'h0);
  reg [(4'ha):(1'h0)] reg1501 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1500 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1499 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1498 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1497 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1496 = (1'h0);
  reg [(4'hb):(1'h0)] reg1495 = (1'h0);
  reg [(5'h12):(1'h0)] reg1494 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1493 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1492 = (1'h0);
  reg [(3'h5):(1'h0)] reg1491 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1490 = (1'h0);
  reg [(4'hc):(1'h0)] reg1489 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire1488;
  wire signed [(4'h8):(1'h0)] wire1487;
  reg [(4'he):(1'h0)] reg1486 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire1485;
  reg signed [(3'h7):(1'h0)] reg1484 = (1'h0);
  reg [(2'h3):(1'h0)] reg1483 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire1482;
  wire [(4'h8):(1'h0)] wire1481;
  reg signed [(4'hc):(1'h0)] reg1480 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1479 = (1'h0);
  reg [(5'h13):(1'h0)] reg1478 = (1'h0);
  reg [(5'h12):(1'h0)] reg1477 = (1'h0);
  assign y = {wire1507,
                 reg1506,
                 reg1505,
                 reg1504,
                 wire1503,
                 reg1502,
                 reg1501,
                 reg1500,
                 reg1499,
                 reg1498,
                 reg1497,
                 forvar1496,
                 reg1495,
                 reg1494,
                 reg1493,
                 forvar1492,
                 reg1491,
                 forvar1490,
                 reg1489,
                 wire1488,
                 wire1487,
                 reg1486,
                 wire1485,
                 reg1484,
                 reg1483,
                 wire1482,
                 wire1481,
                 reg1480,
                 reg1479,
                 reg1478,
                 reg1477,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1477 <= wire1474;
      reg1478 <= ($signed(wire1475[(1'h1):(1'h0)]) ?
          (wire1474 <<< (wire1474 ?
              ((wire1475 > (7'h42)) || $unsigned(wire1474)) : $unsigned((wire1473 >>> wire1474)))) : ({{(^wire1474),
                  (wire1476 ^~ reg1477)},
              ((wire1475 ? wire1475 : wire1475) ?
                  wire1473 : (wire1474 ? reg1477 : wire1475))} > {(8'ha4)}));
      reg1479 <= $unsigned(reg1477[(2'h2):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg1480 <= $unsigned((wire1476 == (~&(^~(reg1479 ?
          reg1478 : wire1476)))));
    end
  assign wire1481 = ((^~(!(|$unsigned(reg1477)))) ?
                        (^~$unsigned(($signed(reg1477) ?
                            (reg1480 ?
                                reg1479 : reg1478) : $signed(wire1474)))) : (($unsigned(wire1473) ^ ($signed(wire1473) <= {wire1473})) ?
                            $unsigned((reg1478[(4'hc):(3'h6)] ?
                                reg1478[(4'ha):(2'h3)] : wire1473[(4'hf):(4'hf)])) : {(^reg1478)}));
  assign wire1482 = $signed(wire1476);
  always
    @(posedge clk) begin
      reg1483 <= (reg1478 ? $unsigned($signed(wire1473)) : reg1477);
      reg1484 <= $unsigned($signed(reg1480[(4'hb):(4'ha)]));
    end
  assign wire1485 = (^~(~|reg1480[(3'h5):(1'h0)]));
  always
    @(posedge clk) begin
      reg1486 = wire1476;
    end
  assign wire1487 = {reg1478[(1'h0):(1'h0)]};
  assign wire1488 = $signed((($unsigned(wire1473) ?
                        ((&reg1478) || reg1483[(1'h1):(1'h0)]) : $unsigned(reg1486[(4'hc):(3'h6)])) && {($signed(reg1480) > (wire1487 && wire1475))}));
  always
    @(posedge clk) begin
      reg1489 <= $signed(wire1481[(3'h7):(2'h2)]);
      for (forvar1490 = (1'h0); (forvar1490 < (3'h4)); forvar1490 = (forvar1490 + (1'h1)))
        begin
          reg1491 = ($signed((~^{$signed((8'hb1)), reg1483})) || reg1486);
          for (forvar1492 = (1'h0); (forvar1492 < (2'h3)); forvar1492 = (forvar1492 + (1'h1)))
            begin
              reg1493 <= {(forvar1490[(3'h5):(3'h4)] >> $unsigned(reg1486)),
                  reg1477};
              reg1494 = $unsigned(({{(^~reg1493), $unsigned(wire1475)},
                      {{reg1477}, reg1486}} ?
                  wire1475[(2'h2):(2'h2)] : wire1476[(2'h2):(1'h1)]));
            end
          reg1495 <= wire1473[(5'h13):(4'ha)];
        end
      for (forvar1496 = (1'h0); (forvar1496 < (2'h3)); forvar1496 = (forvar1496 + (1'h1)))
        begin
          reg1497 <= $signed((&(8'h9f)));
          reg1498 <= ((wire1481[(3'h4):(1'h1)] ?
              ((-(forvar1490 < wire1485)) <<< $unsigned(reg1478[(5'h11):(3'h4)])) : wire1488[(2'h2):(2'h2)]) != reg1495[(2'h3):(1'h1)]);
          reg1499 <= $unsigned(reg1493);
          reg1500 = $signed((forvar1496 ?
              $unsigned($signed($signed((8'haf)))) : {(^((8'hb6) <<< forvar1492))}));
          reg1501 <= $unsigned(wire1475[(3'h6):(3'h5)]);
        end
    end
  always
    @(posedge clk) begin
      reg1502 <= wire1473;
    end
  assign wire1503 = $unsigned($unsigned((|(reg1497[(3'h4):(1'h1)] ?
                        {wire1487} : $signed(reg1478)))));
  always
    @(posedge clk) begin
      reg1504 <= $signed($signed($unsigned({reg1479, $unsigned(reg1494)})));
      reg1505 <= (~$unsigned((~|((forvar1490 | (8'haf)) ?
          (reg1493 > wire1488) : (reg1483 <<< (8'hb2))))));
      reg1506 = (((|reg1495) ?
          (!(8'hb2)) : $signed(reg1505[(3'h5):(2'h2)])) & wire1476);
    end
  assign wire1507 = $unsigned({$unsigned(({reg1502, wire1474} ?
                            (~&wire1482) : $unsigned(reg1498)))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1718
#( parameter param1884 = ((((((7'h43) ? (8'hb7) : (8'had)) ~^ {(8'ha0), (8'hb9)}) ? (((8'hbd) >>> (8'hab)) ? ((8'hb8) && (8'ha3)) : ((8'had) ? (8'ha0) : (8'hb1))) : (^(~^(8'ha9)))) ? (({(8'ha9), (8'hb8)} ^ ((8'ha1) <= (8'ha8))) ? (((8'hbe) < (8'ha4)) && ((8'haf) > (8'hb8))) : {(!(8'hb3)), ((8'hb9) && (8'hac))}) : (|(((8'ha5) ? (8'ha4) : (8'ha6)) ^ (7'h42)))) ^ {(-(((8'hb4) ? (8'hbe) : (8'h9f)) || (-(8'hb0))))}) )
(y, clk, wire1723, wire1722, wire1721, wire1720, wire1719);
  output wire [(32'h130):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire1723;
  input wire [(4'hf):(1'h0)] wire1722;
  input wire [(5'h12):(1'h0)] wire1721;
  input wire signed [(5'h15):(1'h0)] wire1720;
  input wire [(4'h8):(1'h0)] wire1719;
  wire signed [(5'h10):(1'h0)] wire1883;
  wire [(2'h2):(1'h0)] wire1757;
  wire signed [(4'h8):(1'h0)] wire1759;
  reg signed [(4'ha):(1'h0)] forvar1760 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1761 = (1'h0);
  reg [(4'hc):(1'h0)] reg1762 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1763 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1764 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1765 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1766 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1767 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1768 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1769 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1770 = (1'h0);
  reg [(3'h7):(1'h0)] reg1771 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1772 = (1'h0);
  reg [(5'h15):(1'h0)] reg1773 = (1'h0);
  reg [(4'ha):(1'h0)] reg1774 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1775 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1776 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1777 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1778 = (1'h0);
  wire [(4'ha):(1'h0)] wire1779;
  wire [(5'h13):(1'h0)] wire1780;
  wire [(4'hb):(1'h0)] wire1881;
  assign y = {wire1883,
                 wire1757,
                 wire1759,
                 forvar1760,
                 reg1761,
                 reg1762,
                 reg1763,
                 reg1764,
                 reg1765,
                 reg1766,
                 reg1767,
                 forvar1768,
                 reg1769,
                 forvar1770,
                 reg1771,
                 reg1772,
                 reg1773,
                 reg1774,
                 reg1775,
                 reg1776,
                 reg1777,
                 reg1778,
                 wire1779,
                 wire1780,
                 wire1881,
                 (1'h0)};
  module1724 modinst1758 (wire1757, clk, wire1721, wire1723, wire1720, wire1722, wire1719);
  assign wire1759 = $signed((((((8'hb4) * wire1722) ?
                            (wire1721 != wire1721) : wire1723[(4'h8):(2'h2)]) * wire1723) ?
                        ($unsigned((~^wire1757)) ?
                            wire1722 : $signed(wire1757[(1'h0):(1'h0)])) : wire1719[(1'h1):(1'h1)]));
  always
    @(posedge clk) begin
      for (forvar1760 = (1'h0); (forvar1760 < (3'h4)); forvar1760 = (forvar1760 + (1'h1)))
        begin
          reg1761 <= wire1722;
          reg1762 <= {(({(~|(7'h44)), $signed(reg1761)} + (+(wire1719 ?
                  wire1719 : wire1721))) ^ wire1720),
              $signed(wire1721[(4'hd):(3'h6)])};
        end
      reg1763 <= (($signed(wire1757) ?
          ((~&{(8'hbe), wire1759}) ?
              (wire1722[(4'ha):(4'h8)] ?
                  $unsigned((8'hb9)) : $signed(wire1722)) : reg1761[(2'h2):(1'h1)]) : wire1723[(4'hf):(4'h8)]) == (+wire1723[(3'h4):(2'h3)]));
      reg1764 <= $unsigned(forvar1760[(2'h3):(1'h0)]);
      reg1765 <= reg1764[(2'h2):(2'h2)];
    end
  always
    @(posedge clk) begin
      reg1766 <= wire1721;
    end
  always
    @(posedge clk) begin
      reg1767 = (!$unsigned(forvar1760[(4'h9):(2'h2)]));
      for (forvar1768 = (1'h0); (forvar1768 < (2'h3)); forvar1768 = (forvar1768 + (1'h1)))
        begin
          reg1769 <= wire1721[(2'h3):(2'h2)];
          for (forvar1770 = (1'h0); (forvar1770 < (3'h4)); forvar1770 = (forvar1770 + (1'h1)))
            begin
              reg1771 <= wire1720[(2'h3):(2'h3)];
              reg1772 <= ($signed($unsigned(((+reg1762) ?
                  reg1762 : (wire1723 <= wire1720)))) + {wire1721});
              reg1773 <= (($unsigned((reg1769[(2'h2):(1'h1)] ?
                  $signed(reg1771) : $unsigned(forvar1760))) > (&((wire1759 ?
                  forvar1760 : wire1723) || reg1772))) >>> $signed({reg1761}));
              reg1774 = reg1762[(4'hc):(1'h1)];
            end
          reg1775 <= $signed({$unsigned(reg1769[(3'h5):(1'h1)])});
        end
      reg1776 <= forvar1770;
      reg1777 = wire1759[(2'h2):(1'h1)];
      reg1778 = ({reg1761[(4'h9):(3'h6)], reg1762[(4'h9):(3'h6)]} ?
          (reg1761 ?
              $unsigned($unsigned($unsigned(wire1722))) : $signed($signed(reg1775))) : reg1765[(3'h6):(2'h2)]);
    end
  assign wire1779 = (forvar1760 ?
                        ({$signed(((8'h9e) ? reg1773 : reg1762)),
                                reg1765[(3'h5):(2'h2)]} ?
                            wire1719[(3'h7):(2'h3)] : (!$unsigned((reg1771 ?
                                wire1722 : (8'hb5))))) : wire1723);
  assign wire1780 = $unsigned(((8'hb5) >>> reg1772[(4'hc):(2'h3)]));
  module1781 modinst1882 (.wire1782(reg1767), .wire1784(wire1780), .wire1785(wire1720), .wire1783(wire1722), .wire1786(reg1772), .y(wire1881), .clk(clk));
  assign wire1883 = (8'had);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1781
#( parameter param1880 = ((((7'h44) <= ((^(8'hb0)) ? (-(8'hbe)) : ((8'hb1) ? (8'hbf) : (8'ha4)))) == ((((7'h44) == (8'h9d)) ? (8'hbe) : (-(7'h42))) ? (((8'hbb) ? (8'hbc) : (8'hac)) | {(8'hb9), (8'hac)}) : (~^{(8'hbc)}))) ? {((((8'h9e) ? (8'hb3) : (8'hb3)) ? (~&(8'ha9)) : {(8'ha2)}) >> (+((8'ha1) ? (8'ha0) : (8'hb3))))} : {(8'hae), (~(((8'ha3) > (8'hab)) | {(8'hba), (8'hb5)}))}) )
(y, clk, wire1786, wire1785, wire1784, wire1783, wire1782);
  output wire [(32'h43e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire1786;
  input wire signed [(2'h2):(1'h0)] wire1785;
  input wire [(5'h13):(1'h0)] wire1784;
  input wire [(4'hf):(1'h0)] wire1783;
  input wire [(3'h7):(1'h0)] wire1782;
  wire [(4'hd):(1'h0)] wire1879;
  reg [(4'h8):(1'h0)] reg1878 = (1'h0);
  reg [(4'hb):(1'h0)] reg1877 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1876 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1875 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1874 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1873 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1872 = (1'h0);
  reg [(2'h3):(1'h0)] reg1871 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1868 = (1'h0);
  reg [(5'h10):(1'h0)] reg1870 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1869 = (1'h0);
  reg [(3'h5):(1'h0)] reg1868 = (1'h0);
  reg [(3'h5):(1'h0)] reg1867 = (1'h0);
  wire [(5'h13):(1'h0)] wire1866;
  wire signed [(4'ha):(1'h0)] wire1865;
  wire [(3'h6):(1'h0)] wire1864;
  reg signed [(4'he):(1'h0)] reg1863 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1862 = (1'h0);
  reg [(5'h10):(1'h0)] reg1861 = (1'h0);
  reg [(3'h7):(1'h0)] reg1860 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1859 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1858 = (1'h0);
  reg [(4'hc):(1'h0)] reg1857 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1856 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1855 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1854 = (1'h0);
  reg [(2'h3):(1'h0)] reg1853 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1852 = (1'h0);
  reg [(3'h7):(1'h0)] reg1851 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1850 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1849 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1848 = (1'h0);
  reg [(4'he):(1'h0)] forvar1847 = (1'h0);
  reg [(5'h12):(1'h0)] reg1846 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1845 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1844 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1843 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1842 = (1'h0);
  reg [(2'h3):(1'h0)] reg1841 = (1'h0);
  reg [(2'h3):(1'h0)] reg1840 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1839 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1838 = (1'h0);
  reg [(4'hf):(1'h0)] reg1837 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1836 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1835 = (1'h0);
  wire [(5'h13):(1'h0)] wire1834;
  reg signed [(3'h4):(1'h0)] reg1833 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1832 = (1'h0);
  reg [(3'h6):(1'h0)] reg1831 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire1830;
  reg [(2'h3):(1'h0)] reg1829 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1828 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1827 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1826 = (1'h0);
  reg [(5'h12):(1'h0)] reg1825 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1824 = (1'h0);
  reg [(5'h15):(1'h0)] reg1823 = (1'h0);
  reg [(3'h4):(1'h0)] reg1822 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1821 = (1'h0);
  reg [(4'hf):(1'h0)] reg1820 = (1'h0);
  reg [(4'he):(1'h0)] reg1819 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1818 = (1'h0);
  reg [(4'hc):(1'h0)] reg1817 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1816 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1815 = (1'h0);
  reg [(5'h14):(1'h0)] reg1814 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1813 = (1'h0);
  wire [(5'h14):(1'h0)] wire1812;
  reg signed [(4'h9):(1'h0)] reg1811 = (1'h0);
  reg [(5'h10):(1'h0)] reg1810 = (1'h0);
  reg [(5'h12):(1'h0)] reg1809 = (1'h0);
  reg [(5'h14):(1'h0)] reg1808 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1807 = (1'h0);
  reg [(5'h12):(1'h0)] reg1806 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1805 = (1'h0);
  reg [(5'h15):(1'h0)] reg1804 = (1'h0);
  reg [(5'h11):(1'h0)] reg1803 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1802 = (1'h0);
  reg [(2'h3):(1'h0)] reg1801 = (1'h0);
  reg [(5'h13):(1'h0)] reg1800 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1799 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1798 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1797 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1796 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1795 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire1794;
  reg [(3'h6):(1'h0)] reg1793 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1792 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1791 = (1'h0);
  reg [(2'h2):(1'h0)] reg1790 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1789 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1788 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1787 = (1'h0);
  assign y = {wire1879,
                 reg1878,
                 reg1877,
                 reg1876,
                 reg1875,
                 forvar1874,
                 reg1873,
                 reg1872,
                 reg1871,
                 forvar1868,
                 reg1870,
                 reg1869,
                 reg1868,
                 reg1867,
                 wire1866,
                 wire1865,
                 wire1864,
                 reg1863,
                 reg1862,
                 reg1861,
                 reg1860,
                 reg1859,
                 reg1858,
                 reg1857,
                 reg1856,
                 reg1855,
                 forvar1854,
                 reg1853,
                 reg1852,
                 reg1851,
                 reg1850,
                 reg1849,
                 reg1848,
                 forvar1847,
                 reg1846,
                 reg1845,
                 forvar1844,
                 reg1843,
                 forvar1842,
                 reg1841,
                 reg1840,
                 reg1839,
                 reg1838,
                 reg1837,
                 forvar1836,
                 reg1835,
                 wire1834,
                 reg1833,
                 reg1832,
                 reg1831,
                 wire1830,
                 reg1829,
                 reg1828,
                 reg1827,
                 forvar1826,
                 reg1825,
                 reg1824,
                 reg1823,
                 reg1822,
                 forvar1821,
                 reg1820,
                 reg1819,
                 forvar1818,
                 reg1817,
                 reg1816,
                 forvar1815,
                 reg1814,
                 reg1813,
                 wire1812,
                 reg1811,
                 reg1810,
                 reg1809,
                 reg1808,
                 reg1807,
                 reg1806,
                 forvar1805,
                 reg1804,
                 reg1803,
                 forvar1802,
                 reg1801,
                 reg1800,
                 reg1799,
                 reg1798,
                 forvar1797,
                 reg1796,
                 reg1795,
                 wire1794,
                 reg1793,
                 reg1792,
                 reg1791,
                 reg1790,
                 reg1789,
                 reg1788,
                 forvar1787,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar1787 = (1'h0); (forvar1787 < (1'h1)); forvar1787 = (forvar1787 + (1'h1)))
        begin
          if (wire1782[(3'h6):(1'h0)])
            begin
              reg1788 <= ($unsigned($unsigned(forvar1787[(2'h3):(2'h2)])) + (($unsigned($signed((7'h43))) << (^~(wire1783 ?
                      wire1784 : wire1782))) ?
                  $signed((~&$unsigned(wire1785))) : (wire1782[(1'h1):(1'h1)] | (|(wire1785 != forvar1787)))));
              reg1789 = (+$signed(wire1782[(1'h0):(1'h0)]));
              reg1790 <= (($signed($unsigned(wire1784[(3'h6):(1'h0)])) ?
                  {{(8'hbc)}} : {($signed(reg1789) << (7'h44))}) >= {(reg1789 ?
                      $signed({wire1786, forvar1787}) : (((8'ha1) ?
                          wire1783 : (8'hae)) + (wire1782 > wire1786))),
                  $unsigned((|wire1785))});
            end
          else
            begin
              reg1788 <= $signed(wire1782);
              reg1789 = ((8'hbf) ^ forvar1787);
              reg1790 = $signed(wire1782);
            end
          reg1791 <= (&wire1782);
          reg1792 <= (8'ha2);
          reg1793 <= reg1791;
        end
    end
  assign wire1794 = $signed((|(^~(reg1788 ?
                        (wire1784 ? reg1789 : reg1788) : (reg1792 ?
                            reg1792 : reg1788)))));
  always
    @(posedge clk) begin
      reg1795 <= (|$signed($unsigned(wire1782[(2'h2):(1'h1)])));
      reg1796 = (wire1784[(5'h11):(4'he)] & wire1794[(1'h0):(1'h0)]);
      for (forvar1797 = (1'h0); (forvar1797 < (2'h3)); forvar1797 = (forvar1797 + (1'h1)))
        begin
          reg1798 <= reg1788;
          reg1799 = ($unsigned((&$signed(wire1785[(1'h1):(1'h0)]))) <= (wire1783 ^ reg1791));
          reg1800 <= reg1792[(3'h4):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      reg1801 <= (wire1786 * {$signed(((reg1793 ?
              wire1784 : wire1794) || reg1800[(4'h8):(4'h8)]))});
      for (forvar1802 = (1'h0); (forvar1802 < (2'h2)); forvar1802 = (forvar1802 + (1'h1)))
        begin
          reg1803 = forvar1802;
          reg1804 <= $signed(reg1795);
        end
      for (forvar1805 = (1'h0); (forvar1805 < (3'h4)); forvar1805 = (forvar1805 + (1'h1)))
        begin
          reg1806 <= {$unsigned((^~wire1785[(1'h0):(1'h0)])),
              ($unsigned(reg1803[(4'hc):(2'h3)]) ?
                  reg1793[(1'h0):(1'h0)] : forvar1805)};
          reg1807 <= forvar1805;
          reg1808 <= reg1788;
          reg1809 <= $unsigned({{{$signed(forvar1797), $unsigned(reg1790)}},
              $unsigned(forvar1787)});
        end
      reg1810 = ((wire1794 ?
              {$unsigned(wire1782)} : $unsigned($signed((forvar1805 & reg1798)))) ?
          $unsigned(forvar1787) : (-reg1796));
      reg1811 <= (-$signed((wire1785[(1'h0):(1'h0)] ?
          ($unsigned(wire1794) & (^reg1801)) : {(!reg1806)})));
    end
  assign wire1812 = wire1786;
  always
    @(posedge clk) begin
      reg1813 <= reg1792[(1'h1):(1'h0)];
      reg1814 = $unsigned({{($unsigned(reg1789) ?
                  $signed(wire1786) : reg1793)}});
    end
  always
    @(posedge clk) begin
      for (forvar1815 = (1'h0); (forvar1815 < (1'h1)); forvar1815 = (forvar1815 + (1'h1)))
        begin
          reg1816 <= reg1814;
          reg1817 <= (~|$signed((~reg1795)));
          for (forvar1818 = (1'h0); (forvar1818 < (2'h2)); forvar1818 = (forvar1818 + (1'h1)))
            begin
              reg1819 = $unsigned($unsigned((+$signed((forvar1802 ?
                  reg1796 : (8'ha2))))));
              reg1820 <= $unsigned(wire1794);
            end
          for (forvar1821 = (1'h0); (forvar1821 < (2'h3)); forvar1821 = (forvar1821 + (1'h1)))
            begin
              reg1822 <= reg1804;
            end
          reg1823 = reg1807[(4'hc):(3'h5)];
        end
      reg1824 <= reg1800[(4'hf):(1'h1)];
      reg1825 <= ($unsigned(((-(reg1803 != reg1808)) ?
          {(reg1820 ?
                  (8'hbf) : reg1811)} : wire1794[(2'h2):(2'h2)])) | {(wire1786[(2'h3):(1'h1)] ?
              {$signed(reg1800),
                  ((8'h9d) ? reg1800 : wire1786)} : {reg1792[(1'h1):(1'h1)],
                  (+reg1810)}),
          (((reg1804 ? wire1783 : (8'hb5)) & (|reg1793)) ?
              (wire1794 - $signed(reg1810)) : (reg1810 ^~ forvar1818))});
      for (forvar1826 = (1'h0); (forvar1826 < (2'h3)); forvar1826 = (forvar1826 + (1'h1)))
        begin
          reg1827 <= forvar1797;
          reg1828 <= (~|(reg1809[(5'h12):(3'h5)] ?
              ($signed($signed(reg1820)) - ({reg1801} | (reg1801 < (8'ha0)))) : (forvar1826 ?
                  (~^(!wire1782)) : reg1796[(4'h8):(3'h5)])));
          reg1829 = (8'hb5);
        end
    end
  assign wire1830 = $signed(($signed(reg1793) <= $signed(reg1798)));
  always
    @(posedge clk) begin
      reg1831 = $signed((reg1798[(3'h5):(2'h2)] ?
          {{{(8'hbd)}},
              {$signed((8'hb9)),
                  (forvar1802 ?
                      reg1807 : (8'hbb))}} : {(reg1824 < (!reg1824))}));
      reg1832 = ({$signed($unsigned($unsigned(reg1813)))} ?
          ((reg1792 ?
              $unsigned($signed((8'hb1))) : (~|wire1830[(4'h8):(2'h3)])) >> forvar1797[(4'h9):(3'h7)]) : $unsigned(($unsigned({wire1785}) ?
              $unsigned(reg1817) : {$unsigned(reg1803)})));
      reg1833 <= (reg1820[(4'h8):(4'h8)] < forvar1805);
    end
  assign wire1834 = (^~{forvar1815[(2'h2):(1'h0)], reg1800});
  always
    @(posedge clk) begin
      reg1835 <= (~&reg1799);
      for (forvar1836 = (1'h0); (forvar1836 < (1'h0)); forvar1836 = (forvar1836 + (1'h1)))
        begin
          reg1837 <= $signed($signed($unsigned(($unsigned(reg1825) && $signed(reg1811)))));
          reg1838 <= $unsigned((wire1830 | forvar1787));
          reg1839 <= (($unsigned(wire1812) >>> reg1835) ?
              (~^($unsigned({reg1789,
                  reg1801}) >> reg1817[(4'h8):(4'h8)])) : {(((!forvar1826) != $unsigned(reg1824)) != $unsigned($signed(reg1810))),
                  {$unsigned((reg1793 | wire1786)),
                      {reg1810, $unsigned(reg1822)}}});
        end
      reg1840 <= forvar1787[(3'h6):(2'h2)];
      reg1841 <= reg1796;
      for (forvar1842 = (1'h0); (forvar1842 < (1'h0)); forvar1842 = (forvar1842 + (1'h1)))
        begin
          reg1843 <= $unsigned((!((~&(~&reg1790)) == $signed($signed((8'hac))))));
          for (forvar1844 = (1'h0); (forvar1844 < (2'h2)); forvar1844 = (forvar1844 + (1'h1)))
            begin
              reg1845 = (+reg1811);
              reg1846 <= ((reg1845[(1'h0):(1'h0)] ?
                      (reg1841[(1'h1):(1'h0)] ?
                          $unsigned($unsigned(reg1839)) : ((^reg1807) ?
                              reg1824[(3'h4):(2'h3)] : (8'hb3))) : reg1793) ?
                  {((reg1839[(1'h1):(1'h1)] && (reg1804 | reg1832)) ?
                          $signed((~&reg1800)) : (-(+reg1800))),
                      $signed($signed(forvar1787))} : {(8'hb2),
                      $unsigned(reg1801[(1'h0):(1'h0)])});
            end
          for (forvar1847 = (1'h0); (forvar1847 < (1'h0)); forvar1847 = (forvar1847 + (1'h1)))
            begin
              reg1848 <= {(^~(($signed(reg1819) == reg1788) * (&wire1782)))};
              reg1849 <= $unsigned(($unsigned(wire1782) ?
                  (^~$signed((+reg1816))) : $unsigned(((reg1810 * reg1823) ?
                      $signed(reg1813) : (reg1841 ? reg1792 : wire1812)))));
              reg1850 <= ($unsigned($unsigned((((8'ha8) ?
                      (8'hbf) : forvar1805) ?
                  $signed(wire1830) : (^~wire1784)))) > ({((+reg1809) >>> (reg1840 >>> (8'hae)))} || $unsigned(reg1831[(3'h6):(3'h5)])));
            end
        end
    end
  always
    @(posedge clk) begin
      reg1851 <= $unsigned(reg1789);
      reg1852 <= (|(8'hab));
      reg1853 <= (^forvar1787);
    end
  always
    @(posedge clk) begin
      for (forvar1854 = (1'h0); (forvar1854 < (2'h3)); forvar1854 = (forvar1854 + (1'h1)))
        begin
          reg1855 <= (reg1832 && $unsigned((|$unsigned($signed(reg1819)))));
          reg1856 <= reg1829;
          reg1857 = forvar1844[(5'h12):(4'hd)];
          reg1858 <= (~&forvar1805);
          reg1859 = ((~&{$unsigned({reg1793}),
                  $signed(reg1810[(4'hd):(3'h6)])}) ?
              reg1807[(2'h2):(1'h0)] : forvar1844[(5'h12):(3'h4)]);
        end
      reg1860 <= ($signed(((reg1799[(4'h8):(3'h6)] ?
          (8'hb9) : reg1810[(4'hd):(4'hb)]) | ((~&forvar1815) + reg1807))) < reg1839[(1'h1):(1'h0)]);
      reg1861 = $unsigned((({$signed(reg1827)} > $signed((~|(8'h9e)))) ?
          ($signed($signed(wire1783)) - reg1803) : $unsigned($signed($unsigned(reg1835)))));
      reg1862 <= ($signed($signed($signed((reg1827 & (8'hb6))))) ^ reg1806[(2'h2):(2'h2)]);
      reg1863 <= {(((|(wire1786 << reg1824)) | reg1851[(3'h4):(2'h2)]) | (wire1782 ?
              ($signed(reg1837) ?
                  (reg1790 ?
                      (8'ha6) : (8'hb3)) : reg1811) : $unsigned((reg1833 ?
                  forvar1854 : (8'hbf)))))};
    end
  assign wire1864 = reg1811[(1'h1):(1'h1)];
  assign wire1865 = $signed({{$unsigned({reg1857})}});
  assign wire1866 = {reg1799};
  always
    @(posedge clk) begin
      reg1867 <= reg1829;
    end
  always
    @(posedge clk) begin
      if ($unsigned((-(8'ha1))))
        begin
          reg1868 <= reg1829;
          reg1869 = $unsigned($signed($signed($unsigned((wire1864 <= reg1819)))));
          reg1870 <= reg1823[(4'hd):(3'h5)];
        end
      else
        begin
          for (forvar1868 = (1'h0); (forvar1868 < (3'h4)); forvar1868 = (forvar1868 + (1'h1)))
            begin
              reg1869 <= $unsigned($signed($unsigned((^~reg1840[(1'h1):(1'h0)]))));
              reg1870 <= reg1791[(3'h5):(3'h5)];
              reg1871 = (+reg1799);
              reg1872 = $unsigned(reg1853[(2'h3):(1'h1)]);
              reg1873 = ((~^({forvar1815, (^~(7'h40))} ?
                      $signed((wire1865 != wire1783)) : (reg1789 >>> reg1793[(3'h6):(3'h5)]))) ?
                  reg1870 : $signed($unsigned($signed($unsigned(wire1866)))));
            end
          for (forvar1874 = (1'h0); (forvar1874 < (1'h0)); forvar1874 = (forvar1874 + (1'h1)))
            begin
              reg1875 <= ((reg1840[(2'h3):(2'h3)] ~^ (~|(|reg1838))) && reg1798);
            end
        end
      reg1876 <= (wire1794[(2'h3):(1'h1)] ?
          (+reg1806[(2'h3):(1'h0)]) : ($signed(((^~(8'h9e)) ^~ (^(8'hb4)))) ?
              $signed(({reg1793, reg1800} ?
                  (wire1794 >> reg1808) : $unsigned(reg1840))) : (&$unsigned(forvar1874))));
      reg1877 <= (reg1816 <<< {((8'hb7) ? (8'hbb) : (|reg1875)),
          reg1858[(2'h2):(1'h0)]});
      reg1878 <= reg1846[(3'h5):(2'h2)];
    end
  assign wire1879 = (~|((($unsigned((8'hae)) ?
                            wire1866[(1'h1):(1'h1)] : (reg1876 ?
                                (8'h9d) : reg1799)) && reg1807) ?
                        $signed($signed(reg1788)) : $signed(({forvar1797,
                                reg1832} ?
                            (!reg1790) : (|reg1863)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1724  (y, clk, wire1729, wire1728, wire1727, wire1726, wire1725);
  output wire [(32'h166):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire1729;
  input wire [(4'hf):(1'h0)] wire1728;
  input wire [(5'h14):(1'h0)] wire1727;
  input wire [(2'h3):(1'h0)] wire1726;
  input wire signed [(2'h2):(1'h0)] wire1725;
  reg signed [(5'h10):(1'h0)] reg1756 = (1'h0);
  reg [(5'h15):(1'h0)] reg1755 = (1'h0);
  reg [(5'h14):(1'h0)] reg1754 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1753 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1752 = (1'h0);
  reg [(4'hf):(1'h0)] reg1751 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1750 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1749 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1748 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1747 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1746 = (1'h0);
  reg [(4'hd):(1'h0)] reg1745 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire1744;
  wire [(5'h11):(1'h0)] wire1743;
  reg signed [(4'ha):(1'h0)] reg1742 = (1'h0);
  wire [(4'hd):(1'h0)] wire1741;
  wire signed [(5'h14):(1'h0)] wire1740;
  wire signed [(5'h12):(1'h0)] wire1739;
  wire signed [(5'h10):(1'h0)] wire1738;
  reg [(5'h11):(1'h0)] reg1737 = (1'h0);
  reg [(4'hb):(1'h0)] reg1736 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1735 = (1'h0);
  reg [(5'h13):(1'h0)] reg1734 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1733 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1732 = (1'h0);
  wire [(4'ha):(1'h0)] wire1731;
  wire signed [(2'h2):(1'h0)] wire1730;
  assign y = {reg1756,
                 reg1755,
                 reg1754,
                 reg1753,
                 reg1752,
                 reg1751,
                 reg1750,
                 forvar1749,
                 reg1748,
                 reg1747,
                 forvar1746,
                 reg1745,
                 wire1744,
                 wire1743,
                 reg1742,
                 wire1741,
                 wire1740,
                 wire1739,
                 wire1738,
                 reg1737,
                 reg1736,
                 reg1735,
                 reg1734,
                 reg1733,
                 forvar1732,
                 wire1731,
                 wire1730,
                 (1'h0)};
  assign wire1730 = $signed((~^wire1728[(4'ha):(3'h7)]));
  assign wire1731 = $signed($signed($signed(({wire1726,
                        wire1730} * $signed(wire1727)))));
  always
    @(posedge clk) begin
      for (forvar1732 = (1'h0); (forvar1732 < (3'h4)); forvar1732 = (forvar1732 + (1'h1)))
        begin
          reg1733 <= $unsigned(wire1730);
        end
      reg1734 <= $signed(wire1725[(1'h1):(1'h1)]);
      reg1735 <= {$unsigned((&(wire1726 ? wire1725 : (+wire1726)))),
          $unsigned((&{wire1726[(1'h1):(1'h1)]}))};
      reg1736 <= forvar1732[(1'h1):(1'h0)];
      reg1737 <= (($signed(wire1729[(2'h2):(2'h2)]) + ((|$signed(wire1727)) ?
              $unsigned({wire1729}) : wire1730[(2'h2):(1'h1)])) ?
          wire1728[(1'h1):(1'h1)] : reg1734);
    end
  assign wire1738 = (-wire1729[(5'h12):(4'he)]);
  assign wire1739 = $unsigned($unsigned($unsigned(((|(8'ha2)) <= (~&wire1727)))));
  assign wire1740 = reg1737;
  assign wire1741 = (wire1740 ?
                        wire1729[(5'h12):(1'h0)] : (reg1734[(4'hf):(4'ha)] ^ ($unsigned($signed(wire1738)) ?
                            (~&((8'ha8) < (8'hbf))) : wire1729[(5'h12):(4'he)])));
  always
    @(posedge clk) begin
      reg1742 <= reg1737;
    end
  assign wire1743 = ({reg1733, wire1739[(4'ha):(4'ha)]} <<< {wire1728,
                        wire1738});
  assign wire1744 = (reg1735 & $signed((&(wire1740[(5'h12):(4'h8)] >> (wire1740 ?
                        reg1737 : reg1736)))));
  always
    @(posedge clk) begin
      reg1745 <= $unsigned((~$signed(((wire1739 ? wire1741 : (8'hae)) ?
          {wire1739} : $unsigned(wire1740)))));
      for (forvar1746 = (1'h0); (forvar1746 < (2'h2)); forvar1746 = (forvar1746 + (1'h1)))
        begin
          reg1747 <= $signed(wire1739);
          reg1748 <= wire1739;
          for (forvar1749 = (1'h0); (forvar1749 < (1'h0)); forvar1749 = (forvar1749 + (1'h1)))
            begin
              reg1750 <= $signed((&{$signed($unsigned(wire1744))}));
            end
          reg1751 <= ($unsigned((($signed(forvar1732) ?
                  wire1731[(1'h0):(1'h0)] : $unsigned((8'ha4))) ?
              wire1727[(5'h10):(1'h1)] : (^{wire1741,
                  wire1740}))) + {($signed((wire1729 * forvar1732)) << (~&wire1743)),
              ($signed($unsigned(wire1740)) ?
                  $unsigned(((8'hae) < wire1728)) : wire1739)});
        end
      reg1752 <= (^$signed((-(~$unsigned(wire1738)))));
      if ($signed((reg1734[(2'h2):(1'h0)] >>> $signed((wire1739[(4'he):(4'he)] < wire1729)))))
        begin
          reg1753 <= (reg1751 ?
              wire1740[(5'h11):(3'h6)] : reg1752[(3'h5):(2'h2)]);
        end
      else
        begin
          reg1753 = ({(~|(reg1737[(3'h5):(2'h3)] ^~ (wire1739 ?
                  reg1751 : wire1730)))} | {($signed({wire1725,
                  wire1725}) * (((8'ha5) >> wire1738) + (8'h9c)))});
          reg1754 <= (((^$unsigned((+reg1747))) ?
                  (($signed(reg1753) & (wire1731 ? wire1738 : forvar1746)) ?
                      $unsigned(wire1739) : $signed(forvar1749[(4'h8):(3'h7)])) : (~wire1738[(3'h5):(3'h5)])) ?
              $unsigned(reg1747[(2'h3):(1'h1)]) : reg1752);
          reg1755 <= $signed((-((7'h40) < (~^$signed(reg1747)))));
          reg1756 = wire1744[(3'h4):(2'h3)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2173
#(parameter param2626 = {(7'h40)}, parameter param2627 = (8'hbf))
(y, clk, wire2178, wire2177, wire2176, wire2175, wire2174);
  output wire [(32'h2f3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire2178;
  input wire [(3'h6):(1'h0)] wire2177;
  input wire [(3'h7):(1'h0)] wire2176;
  input wire [(5'h13):(1'h0)] wire2175;
  input wire [(4'hd):(1'h0)] wire2174;
  reg signed [(4'hd):(1'h0)] reg2625 = (1'h0);
  reg [(3'h4):(1'h0)] reg2624 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2623 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2622 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2621 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2620 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2619 = (1'h0);
  reg [(4'he):(1'h0)] reg2618 = (1'h0);
  reg [(4'hf):(1'h0)] reg2617 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2616 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2615 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2614 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2613 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2612 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2611 = (1'h0);
  reg [(4'hb):(1'h0)] reg2610 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2609 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2608 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2607 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire2555;
  wire signed [(3'h5):(1'h0)] wire2393;
  reg [(4'hf):(1'h0)] reg2374 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2369 = (1'h0);
  reg [(4'h8):(1'h0)] reg2367 = (1'h0);
  reg [(4'hc):(1'h0)] reg2373 = (1'h0);
  reg [(5'h15):(1'h0)] reg2372 = (1'h0);
  reg [(3'h7):(1'h0)] reg2371 = (1'h0);
  reg [(4'hb):(1'h0)] reg2370 = (1'h0);
  reg [(5'h13):(1'h0)] reg2369 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2368 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2367 = (1'h0);
  reg [(4'he):(1'h0)] reg2366 = (1'h0);
  wire [(4'hc):(1'h0)] wire2307;
  wire [(4'ha):(1'h0)] wire2252;
  wire signed [(4'hc):(1'h0)] wire2227;
  wire [(5'h13):(1'h0)] wire2185;
  wire signed [(5'h14):(1'h0)] wire2184;
  reg [(5'h12):(1'h0)] reg2183 = (1'h0);
  reg [(5'h14):(1'h0)] reg2182 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire2181;
  wire [(2'h2):(1'h0)] wire2180;
  reg [(4'h9):(1'h0)] reg2179 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2309 = (1'h0);
  reg [(5'h13):(1'h0)] reg2310 = (1'h0);
  reg [(4'hc):(1'h0)] reg2311 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2312 = (1'h0);
  reg [(2'h2):(1'h0)] reg2313 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire2364;
  wire signed [(2'h3):(1'h0)] wire2395;
  reg signed [(4'hf):(1'h0)] reg2396 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2397 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2398 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2399 = (1'h0);
  reg [(5'h14):(1'h0)] reg2400 = (1'h0);
  wire [(5'h12):(1'h0)] wire2401;
  wire [(4'ha):(1'h0)] wire2489;
  wire [(4'hb):(1'h0)] wire2557;
  wire [(5'h15):(1'h0)] wire2605;
  assign y = {reg2625,
                 reg2624,
                 reg2623,
                 reg2622,
                 reg2621,
                 reg2620,
                 reg2619,
                 reg2618,
                 reg2617,
                 reg2616,
                 reg2615,
                 reg2614,
                 reg2613,
                 forvar2612,
                 forvar2611,
                 reg2610,
                 reg2609,
                 reg2608,
                 reg2607,
                 wire2555,
                 wire2393,
                 reg2374,
                 forvar2369,
                 reg2367,
                 reg2373,
                 reg2372,
                 reg2371,
                 reg2370,
                 reg2369,
                 reg2368,
                 forvar2367,
                 reg2366,
                 wire2307,
                 wire2252,
                 wire2227,
                 wire2185,
                 wire2184,
                 reg2183,
                 reg2182,
                 wire2181,
                 wire2180,
                 reg2179,
                 reg2309,
                 reg2310,
                 reg2311,
                 reg2312,
                 reg2313,
                 wire2364,
                 wire2395,
                 reg2396,
                 reg2397,
                 reg2398,
                 reg2399,
                 reg2400,
                 wire2401,
                 wire2489,
                 wire2557,
                 wire2605,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg2179 <= ($signed($unsigned((+wire2176))) ?
          (($unsigned($unsigned(wire2176)) ?
                  $signed((wire2178 ? wire2178 : wire2177)) : wire2176) ?
              ({(wire2178 ? wire2175 : wire2177)} * $signed(((8'ha3) ?
                  wire2176 : wire2177))) : (8'haf)) : (wire2175 ?
              ((|(+wire2174)) ^ $unsigned(wire2178)) : (8'hb2)));
    end
  assign wire2180 = $unsigned(wire2177);
  assign wire2181 = ({(-$signed(wire2174[(4'h9):(4'h9)])),
                        $signed(wire2178[(1'h0):(1'h0)])} > (~wire2174));
  always
    @(posedge clk) begin
      reg2182 = wire2174;
      reg2183 <= (&wire2177);
    end
  assign wire2184 = reg2179;
  assign wire2185 = ((-$signed((^~(~^wire2174)))) ?
                        $unsigned($signed(({wire2175} <= $signed(wire2181)))) : ($unsigned(({reg2179,
                                wire2178} != $signed(wire2174))) ?
                            {(|$signed(wire2180)),
                                wire2178[(3'h6):(3'h4)]} : $signed($signed((wire2180 != wire2184)))));
  module2186 modinst2228 (wire2227, clk, wire2176, wire2178, wire2177, wire2184);
  module2229 modinst2253 (wire2252, clk, wire2184, wire2175, wire2174, wire2181);
  module2254 modinst2308 (.wire2259(wire2184), .clk(clk), .wire2255(wire2177), .wire2256(wire2185), .wire2258(wire2252), .y(wire2307), .wire2257(wire2175));
  always
    @(posedge clk) begin
      reg2309 <= wire2177[(3'h6):(3'h6)];
      reg2310 <= {({(~&reg2182[(3'h5):(3'h5)]),
              $signed($unsigned(wire2176))} >> ((&(~reg2179)) || {$signed(wire2307),
              ((8'hbb) ? wire2177 : wire2178)})),
          ((8'haa) <<< $signed($signed(wire2181[(1'h1):(1'h0)])))};
      reg2311 <= ((reg2183[(3'h6):(3'h4)] ?
              $signed($unsigned($signed((8'ha0)))) : $unsigned(((reg2183 && (8'hab)) ?
                  (wire2185 - wire2184) : $unsigned(wire2178)))) ?
          reg2309 : $signed($signed(wire2177[(3'h5):(3'h5)])));
      reg2312 <= ((({{reg2179}} ^ $signed(wire2180[(1'h0):(1'h0)])) * (((reg2309 ?
              reg2311 : (8'ha4)) ?
          (|wire2307) : reg2183) <<< (!wire2252))) <= ((((reg2183 ~^ wire2181) >>> $signed(wire2174)) ^ ($signed(wire2180) ^~ reg2182[(4'hf):(3'h5)])) ?
          ($unsigned((&wire2184)) ?
              {((8'h9d) ? wire2307 : (8'ha9)),
                  (+reg2310)} : (-(~reg2179))) : (((wire2177 ~^ wire2181) ?
              wire2307[(4'h8):(1'h1)] : {(8'hbe), wire2178}) >= {(wire2176 ?
                  (8'hb3) : wire2175),
              ((7'h40) < wire2177)})));
      reg2313 = (($signed($signed(((8'ha5) + (8'hb4)))) ?
          (wire2177[(2'h2):(2'h2)] >= wire2178[(5'h13):(3'h4)]) : ((wire2184 ?
              {(7'h44),
                  reg2183} : (|wire2307)) ^ $unsigned($unsigned(wire2180)))) << wire2177);
    end
  module2314 modinst2365 (.wire2315(wire2181), .clk(clk), .wire2316(wire2184), .y(wire2364), .wire2319(reg2312), .wire2318(reg2311), .wire2317(reg2309));
  always
    @(posedge clk) begin
      reg2366 <= (($unsigned($unsigned((&reg2182))) ~^ reg2313) ?
          ((((reg2313 ?
                  wire2174 : wire2174) >> $signed(wire2180)) >> (~&(reg2311 * (8'ha7)))) ?
              (&((^~reg2312) || (wire2307 ?
                  wire2184 : wire2185))) : ((wire2177[(3'h6):(2'h2)] ?
                      wire2184[(4'he):(1'h1)] : {wire2174}) ?
                  $signed($unsigned(reg2312)) : (&{reg2182,
                      reg2311}))) : (~^reg2310));
      if ($signed((^wire2181[(3'h6):(1'h0)])))
        begin
          for (forvar2367 = (1'h0); (forvar2367 < (2'h2)); forvar2367 = (forvar2367 + (1'h1)))
            begin
              reg2368 <= {(wire2176[(1'h0):(1'h0)] || {wire2184[(1'h1):(1'h1)]})};
              reg2369 <= (-(wire2178 & reg2179));
              reg2370 <= (8'hb9);
              reg2371 = $signed(wire2185[(5'h13):(4'hb)]);
              reg2372 <= (wire2178 + (reg2369[(1'h1):(1'h1)] ^~ $unsigned((~$signed(reg2313)))));
            end
          reg2373 <= wire2176[(3'h5):(2'h3)];
        end
      else
        begin
          reg2367 <= $unsigned((wire2174 ^ wire2181));
          reg2368 = (~|reg2313);
          for (forvar2369 = (1'h0); (forvar2369 < (2'h2)); forvar2369 = (forvar2369 + (1'h1)))
            begin
              reg2370 <= reg2367;
              reg2371 = {$signed({wire2180,
                      (reg2182[(2'h3):(2'h3)] ?
                          $signed(wire2176) : ((8'hbf) ? wire2184 : reg2366))}),
                  $unsigned(wire2185[(5'h12):(3'h6)])};
              reg2372 <= (^~(reg2313 ?
                  $unsigned(reg2371) : $signed((wire2185[(4'hb):(4'h9)] > reg2182[(4'hf):(3'h7)]))));
              reg2373 <= $unsigned($signed((((|(8'ha3)) ?
                  (forvar2369 ?
                      wire2307 : wire2174) : wire2177[(3'h5):(2'h3)]) >= reg2369)));
            end
          reg2374 = ((((8'ha1) || (wire2307[(4'hb):(4'h9)] << $signed(wire2180))) ?
              {(-$unsigned(wire2177)), wire2175} : (wire2252 ?
                  (((8'h9f) ?
                      wire2178 : reg2371) >= (~|reg2183)) : $unsigned(reg2179[(3'h6):(3'h6)]))) | $unsigned((~$signed($unsigned(reg2183)))));
        end
    end
  module2375 modinst2394 (wire2393, clk, reg2367, wire2181, reg2372, wire2184, wire2177);
  assign wire2395 = (!wire2307[(3'h7):(1'h1)]);
  always
    @(posedge clk) begin
      reg2396 <= reg2370[(4'h9):(4'h9)];
      reg2397 <= reg2366[(3'h5):(3'h5)];
      reg2398 <= $unsigned(wire2364);
      reg2399 <= {((+reg2372) ?
              (&wire2181) : (!({wire2175} ?
                  $unsigned(wire2181) : wire2307[(1'h1):(1'h0)]))),
          forvar2369[(3'h5):(2'h3)]};
    end
  always
    @(posedge clk) begin
      reg2400 = $signed($unsigned(($signed(reg2370[(4'h9):(3'h6)]) & wire2177)));
    end
  assign wire2401 = $unsigned(((^$signed($signed(reg2313))) ^~ (reg2397 ?
                        $signed(((7'h44) ?
                            (8'ha5) : reg2309)) : {$signed(reg2368)})));
  module2402 modinst2490 (wire2489, clk, reg2368, wire2227, reg2374, wire2176, reg2373);
  module2491 modinst2556 (wire2555, clk, reg2373, wire2227, reg2310, wire2184, wire2393);
  assign wire2557 = $unsigned(reg2366);
  module2558 modinst2606 (wire2605, clk, reg2309, wire2555, wire2175, reg2182, wire2174);
  always
    @(posedge clk) begin
      reg2607 <= {(reg2179[(2'h2):(1'h1)] ?
              ($unsigned((wire2174 | wire2176)) & forvar2369) : (+(+$signed(reg2396))))};
      reg2608 <= wire2181[(3'h7):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg2609 <= $unsigned(wire2184);
      reg2610 <= $unsigned($unsigned(((&(wire2307 + wire2227)) ?
          $unsigned($signed(wire2227)) : ($unsigned((8'hba)) | (reg2371 ?
              wire2175 : reg2400)))));
      for (forvar2611 = (1'h0); (forvar2611 < (1'h0)); forvar2611 = (forvar2611 + (1'h1)))
        begin
          for (forvar2612 = (1'h0); (forvar2612 < (2'h2)); forvar2612 = (forvar2612 + (1'h1)))
            begin
              reg2613 <= forvar2611[(4'h8):(2'h3)];
              reg2614 <= $signed($signed($signed(forvar2612[(2'h3):(2'h2)])));
              reg2615 <= (^~(((+(^wire2555)) ?
                  $signed($unsigned(wire2177)) : reg2183[(4'ha):(4'h8)]) + wire2181));
              reg2616 <= {(&{(8'hbd), (~|{(8'hb4), reg2609})}),
                  ({{{reg2370, reg2371}},
                      ((reg2367 <= wire2227) ?
                          wire2184[(5'h14):(3'h6)] : wire2184)} * reg2309)};
              reg2617 <= {{wire2181}};
            end
          reg2618 <= wire2178;
          if ($signed($signed((+(reg2313 * reg2618)))))
            begin
              reg2619 = ($signed(((^~(wire2555 && reg2617)) ?
                      wire2227 : $unsigned((wire2401 ? reg2309 : (8'hbe))))) ?
                  (((!(-reg2373)) ^~ $unsigned((&wire2175))) <= $signed(reg2313[(2'h2):(1'h1)])) : $signed(wire2227));
              reg2620 <= $unsigned(reg2373[(4'h9):(4'h8)]);
              reg2621 <= (({$unsigned($signed(reg2311))} ?
                      wire2364[(4'he):(4'h9)] : (wire2605[(3'h5):(2'h3)] >> ($signed(reg2367) ?
                          forvar2369[(1'h1):(1'h0)] : reg2372))) ?
                  ((reg2369[(5'h11):(3'h4)] ?
                          $signed((8'hbc)) : ($signed((8'haf)) << (-reg2619))) ?
                      $signed($signed((forvar2612 != (8'haf)))) : reg2620) : (^~reg2399[(3'h6):(2'h3)]));
              reg2622 = wire2175;
              reg2623 = $signed({(((^wire2489) ?
                      $signed((8'hac)) : ((8'haa) ~^ reg2400)) == (~^(wire2227 ?
                      reg2309 : reg2310)))});
            end
          else
            begin
              reg2619 <= $unsigned(({$unsigned((reg2374 ?
                      reg2367 : wire2181))} > wire2307));
              reg2620 = wire2227[(4'ha):(3'h4)];
            end
          reg2624 = $signed(((~&$signed($unsigned(reg2366))) & $signed(((reg2310 ?
                  wire2175 : forvar2367) ?
              (forvar2611 <<< (8'ha1)) : reg2313[(1'h0):(1'h0)]))));
          reg2625 <= ((~&reg2371) ?
              {$unsigned(forvar2367[(1'h1):(1'h1)])} : (-$unsigned(reg2622[(3'h4):(2'h2)])));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1930
#( parameter param2169 = ((-((((7'h43) ? (8'hb5) : (7'h41)) ? ((8'hb4) ? (8'hb4) : (8'hbe)) : (~|(8'hbc))) ? ((^~(8'haa)) | ((8'hbc) ? (8'hb4) : (8'hb3))) : (((8'hb2) ? (8'hae) : (8'ha3)) && (~^(7'h44))))) < {(((~|(8'hbc)) | ((8'hb7) ? (7'h44) : (8'hbc))) ? (((8'hb0) - (8'ha2)) ? ((8'hb0) << (8'h9e)) : ((8'h9f) >>> (8'hbf))) : ((+(8'hb6)) ? ((8'hbb) <= (8'ha7)) : (^~(8'hae))))}) )
(y, clk, wire1935, wire1934, wire1933, wire1932, wire1931);
  output wire [(32'h39b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire1935;
  input wire [(4'ha):(1'h0)] wire1934;
  input wire [(5'h14):(1'h0)] wire1933;
  input wire [(5'h14):(1'h0)] wire1932;
  input wire [(3'h7):(1'h0)] wire1931;
  reg [(2'h3):(1'h0)] reg2168 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2167 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2166 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2165 = (1'h0);
  reg [(4'ha):(1'h0)] reg2164 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2163 = (1'h0);
  wire [(4'hf):(1'h0)] wire2162;
  wire [(4'h9):(1'h0)] wire2161;
  reg signed [(5'h13):(1'h0)] reg2160 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2159 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2158 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2157 = (1'h0);
  reg [(5'h15):(1'h0)] reg2156 = (1'h0);
  reg [(5'h13):(1'h0)] reg2155 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2154 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire2153;
  reg signed [(5'h12):(1'h0)] reg2152 = (1'h0);
  reg [(3'h4):(1'h0)] reg2151 = (1'h0);
  reg [(4'he):(1'h0)] reg2150 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2149 = (1'h0);
  reg [(3'h6):(1'h0)] reg2148 = (1'h0);
  reg [(4'hb):(1'h0)] reg2147 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2146 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2145 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2144 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2143 = (1'h0);
  reg [(3'h7):(1'h0)] reg2142 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2141 = (1'h0);
  reg [(4'h9):(1'h0)] reg2140 = (1'h0);
  reg [(3'h6):(1'h0)] reg2139 = (1'h0);
  reg [(4'h8):(1'h0)] reg2138 = (1'h0);
  reg [(4'ha):(1'h0)] reg2137 = (1'h0);
  reg [(5'h13):(1'h0)] reg2136 = (1'h0);
  reg [(2'h2):(1'h0)] reg2135 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2134 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2133 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2132 = (1'h0);
  reg [(5'h12):(1'h0)] reg2131 = (1'h0);
  wire [(5'h13):(1'h0)] wire2130;
  wire [(5'h12):(1'h0)] wire2129;
  reg [(4'hb):(1'h0)] reg2128 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire2127;
  reg [(4'ha):(1'h0)] reg2126 = (1'h0);
  reg [(4'ha):(1'h0)] reg2125 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2124 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2123 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2122 = (1'h0);
  reg [(2'h2):(1'h0)] reg2121 = (1'h0);
  reg [(5'h12):(1'h0)] reg2120 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2119 = (1'h0);
  reg [(5'h10):(1'h0)] reg2118 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2117 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2116 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2115 = (1'h0);
  reg [(2'h2):(1'h0)] reg2114 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar2113 = (1'h0);
  reg [(5'h15):(1'h0)] reg2112 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2111 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2110 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2109 = (1'h0);
  reg [(3'h6):(1'h0)] reg2108 = (1'h0);
  reg [(5'h11):(1'h0)] reg2107 = (1'h0);
  reg [(4'he):(1'h0)] reg2106 = (1'h0);
  reg [(4'h9):(1'h0)] reg2105 = (1'h0);
  wire [(5'h15):(1'h0)] wire2104;
  reg signed [(5'h12):(1'h0)] reg2103 = (1'h0);
  reg [(4'hd):(1'h0)] reg2102 = (1'h0);
  reg [(4'h9):(1'h0)] reg2101 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2100 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2099 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2098 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2097 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire2095;
  wire signed [(5'h15):(1'h0)] wire2001;
  wire signed [(5'h12):(1'h0)] wire2000;
  wire [(5'h13):(1'h0)] wire1999;
  wire [(3'h5):(1'h0)] wire1998;
  wire [(4'hd):(1'h0)] wire1996;
  wire [(5'h10):(1'h0)] wire1936;
  assign y = {reg2168,
                 reg2167,
                 reg2166,
                 forvar2165,
                 reg2164,
                 reg2163,
                 wire2162,
                 wire2161,
                 reg2160,
                 reg2159,
                 reg2158,
                 reg2157,
                 reg2156,
                 reg2155,
                 forvar2154,
                 wire2153,
                 reg2152,
                 reg2151,
                 reg2150,
                 reg2149,
                 reg2148,
                 reg2147,
                 forvar2146,
                 reg2145,
                 reg2144,
                 forvar2143,
                 reg2142,
                 reg2141,
                 reg2140,
                 reg2139,
                 reg2138,
                 reg2137,
                 reg2136,
                 reg2135,
                 forvar2134,
                 forvar2133,
                 reg2132,
                 reg2131,
                 wire2130,
                 wire2129,
                 reg2128,
                 wire2127,
                 reg2126,
                 reg2125,
                 reg2124,
                 forvar2123,
                 reg2122,
                 reg2121,
                 reg2120,
                 reg2119,
                 reg2118,
                 reg2117,
                 forvar2116,
                 reg2115,
                 reg2114,
                 forvar2113,
                 reg2112,
                 reg2111,
                 reg2110,
                 forvar2109,
                 reg2108,
                 reg2107,
                 reg2106,
                 reg2105,
                 wire2104,
                 reg2103,
                 reg2102,
                 reg2101,
                 forvar2100,
                 reg2099,
                 forvar2098,
                 reg2097,
                 wire2095,
                 wire2001,
                 wire2000,
                 wire1999,
                 wire1998,
                 wire1996,
                 wire1936,
                 (1'h0)};
  assign wire1936 = (wire1931 ?
                        wire1935[(4'h8):(1'h1)] : {$unsigned((~{wire1935})),
                            $unsigned(((-wire1933) ?
                                (~&wire1934) : (wire1934 >>> wire1933)))});
  module1937 modinst1997 (wire1996, clk, wire1936, wire1932, wire1931, wire1933);
  assign wire1998 = wire1996;
  assign wire1999 = wire1998;
  assign wire2000 = $signed($unsigned((8'ha8)));
  assign wire2001 = wire1936[(1'h1):(1'h0)];
  module2002 modinst2096 (.y(wire2095), .clk(clk), .wire2006(wire1932), .wire2005(wire2001), .wire2003(wire1996), .wire2004(wire2000));
  always
    @(posedge clk) begin
      reg2097 <= (wire1932[(5'h11):(4'hd)] - (~|$signed($unsigned($signed(wire1936)))));
      for (forvar2098 = (1'h0); (forvar2098 < (2'h2)); forvar2098 = (forvar2098 + (1'h1)))
        begin
          reg2099 <= wire1934[(2'h3):(2'h2)];
          for (forvar2100 = (1'h0); (forvar2100 < (1'h0)); forvar2100 = (forvar2100 + (1'h1)))
            begin
              reg2101 <= $unsigned((wire1932[(3'h7):(3'h4)] ?
                  {((wire1999 ? (8'hac) : wire1934) > $signed(reg2099)),
                      $signed(forvar2098)} : (^~$unsigned($signed(wire1932)))));
            end
          reg2102 <= {$unsigned((^(reg2099 || {wire1934, forvar2098}))),
              wire1998[(2'h2):(1'h0)]};
        end
      reg2103 <= $signed(((|$unsigned((wire1932 ~^ wire2000))) ~^ (8'ha2)));
    end
  assign wire2104 = reg2097;
  always
    @(posedge clk) begin
      if ($signed((^~(wire1935 ?
          (^~(forvar2100 ? reg2101 : reg2097)) : wire1934))))
        begin
          reg2105 <= $signed($signed((|((-(8'ha1)) ^ (wire1932 ?
              wire2104 : wire1933)))));
          reg2106 <= $signed($unsigned({($unsigned(reg2097) ?
                  (|forvar2100) : $signed(forvar2098))}));
          reg2107 <= (((^wire1934[(1'h0):(1'h0)]) ?
                  {$signed((wire2095 ? (8'hac) : (8'hbd))),
                      $signed($signed((8'ha5)))} : $signed($unsigned({wire1935,
                      reg2103}))) ?
              (~|(($unsigned(reg2103) == forvar2100) * (8'hac))) : ($unsigned($unsigned($signed(wire1996))) ?
                  (wire1932 ?
                      (~&$unsigned(wire2000)) : $unsigned((~|forvar2098))) : reg2103));
          reg2108 <= (~wire1999);
        end
      else
        begin
          reg2105 = (($signed(($unsigned(reg2101) ?
              (!(7'h42)) : (-wire1931))) != (^(&reg2101[(3'h7):(2'h3)]))) & $unsigned($signed({{wire1935,
                  wire2001},
              forvar2098[(2'h3):(2'h3)]})));
          reg2106 <= forvar2098[(1'h1):(1'h0)];
          reg2107 <= (forvar2100[(2'h2):(2'h2)] ?
              ((reg2108[(2'h2):(1'h0)] ?
                      $signed($unsigned(wire2000)) : $signed({(8'hae),
                          (8'ha0)})) ?
                  $signed((wire1934 ?
                      reg2101[(3'h4):(1'h1)] : (wire1999 ?
                          reg2103 : wire1931))) : (~|$unsigned((^~reg2106)))) : wire2000);
          reg2108 <= ((+(($unsigned(forvar2100) - $signed(wire1935)) + $signed((^wire1932)))) * wire1999);
        end
      for (forvar2109 = (1'h0); (forvar2109 < (3'h4)); forvar2109 = (forvar2109 + (1'h1)))
        begin
          reg2110 <= (~&$signed($unsigned(wire1931)));
          reg2111 <= $unsigned((|($unsigned($unsigned(wire2001)) == (8'hac))));
        end
      reg2112 <= (wire2104 | (|(((reg2106 ?
          wire2095 : wire1998) <<< $unsigned(wire1934)) * $unsigned({wire1999,
          forvar2109}))));
      for (forvar2113 = (1'h0); (forvar2113 < (3'h4)); forvar2113 = (forvar2113 + (1'h1)))
        begin
          reg2114 <= (|(((wire1932[(2'h2):(1'h1)] ?
                  (~^wire1934) : (reg2111 ? wire1996 : reg2105)) ?
              (&reg2112) : ($unsigned(wire2104) > {reg2108,
                  reg2112})) + forvar2109));
          reg2115 <= wire1931[(1'h1):(1'h1)];
          for (forvar2116 = (1'h0); (forvar2116 < (1'h1)); forvar2116 = (forvar2116 + (1'h1)))
            begin
              reg2117 <= (|$unsigned((~&reg2101[(1'h0):(1'h0)])));
              reg2118 <= (8'hb7);
              reg2119 = $signed($unsigned($signed((!(forvar2113 ?
                  (8'ha1) : wire1931)))));
              reg2120 = reg2115;
              reg2121 <= $unsigned(reg2118);
            end
          reg2122 <= (($unsigned(reg2106) ?
              (wire1998 < (reg2105[(3'h4):(2'h2)] + (~|forvar2098))) : $unsigned(wire1996[(3'h4):(2'h2)])) || (&(wire1933 <= (~|((8'hbf) | reg2117)))));
          for (forvar2123 = (1'h0); (forvar2123 < (2'h2)); forvar2123 = (forvar2123 + (1'h1)))
            begin
              reg2124 <= (^~(~reg2101[(2'h3):(1'h1)]));
              reg2125 = (((-wire2095) ?
                  (wire1934[(3'h4):(3'h4)] ?
                      {(+forvar2116),
                          $unsigned((7'h42))} : $unsigned((forvar2113 >= reg2099))) : (^(+$unsigned(wire2095)))) == {(~&((~&wire1936) ?
                      (reg2112 ? reg2105 : forvar2098) : $signed(wire1999)))});
            end
        end
      reg2126 <= reg2110[(3'h5):(1'h1)];
    end
  assign wire2127 = reg2097[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg2128 <= reg2102;
    end
  assign wire2129 = ((~^(($unsigned(forvar2109) ?
                            {(8'hae),
                                forvar2116} : reg2126[(4'h8):(3'h5)]) >>> $unsigned(((8'ha5) ?
                            reg2125 : reg2111)))) ?
                        ($signed((&(wire1998 ^~ reg2101))) ?
                            (+({(8'hba)} ?
                                (reg2114 ?
                                    reg2119 : (8'ha5)) : (8'h9f))) : $unsigned((~&{forvar2116,
                                (8'hb1)}))) : $signed(reg2125[(3'h5):(3'h5)]));
  assign wire2130 = (reg2122[(1'h1):(1'h0)] ?
                        (!(reg2101 ?
                            $signed($signed(reg2102)) : $unsigned((-reg2126)))) : $signed((forvar2123 ?
                            {(reg2099 || forvar2113),
                                (wire2104 >>> forvar2098)} : (~(reg2128 >= reg2112)))));
  always
    @(posedge clk) begin
      reg2131 <= ($signed($unsigned($signed(reg2112[(5'h14):(3'h7)]))) >> (8'ha1));
      reg2132 <= (~|forvar2109);
    end
  always
    @(posedge clk) begin
      for (forvar2133 = (1'h0); (forvar2133 < (1'h1)); forvar2133 = (forvar2133 + (1'h1)))
        begin
          for (forvar2134 = (1'h0); (forvar2134 < (2'h3)); forvar2134 = (forvar2134 + (1'h1)))
            begin
              reg2135 <= $signed((wire1996 ?
                  $unsigned((wire2104 >>> $signed(reg2120))) : (-reg2105[(3'h7):(2'h3)])));
              reg2136 <= (reg2122[(4'h8):(1'h0)] <<< $unsigned(reg2099));
              reg2137 <= wire1999;
              reg2138 <= reg2121[(1'h1):(1'h1)];
            end
          reg2139 <= reg2137[(2'h3):(2'h2)];
          reg2140 <= (forvar2098 ?
              (~^forvar2100[(4'hd):(4'h9)]) : ((~&(8'ha6)) ?
                  reg2105[(4'h9):(3'h4)] : $unsigned({$signed(wire2130),
                      wire2001})));
        end
    end
  always
    @(posedge clk) begin
      reg2141 <= {($unsigned($signed($unsigned((8'ha0)))) ?
              {((8'h9f) ? $unsigned(reg2119) : $unsigned(wire2104)),
                  $signed((reg2107 || reg2097))} : $unsigned($signed({reg2110}))),
          reg2128};
      reg2142 <= (~$signed((({wire1999, wire2001} ?
          (reg2138 <= reg2135) : ((7'h41) ?
              wire2104 : forvar2116)) ~^ reg2136[(3'h6):(1'h1)])));
      for (forvar2143 = (1'h0); (forvar2143 < (2'h2)); forvar2143 = (forvar2143 + (1'h1)))
        begin
          reg2144 <= forvar2100[(4'h9):(4'h8)];
          reg2145 = $signed($unsigned((-{(~^reg2101), {(8'h9c)}})));
          for (forvar2146 = (1'h0); (forvar2146 < (1'h1)); forvar2146 = (forvar2146 + (1'h1)))
            begin
              reg2147 <= (~^({({wire1934, wire1933} ?
                          (-reg2124) : (reg2110 ? wire2001 : reg2140)),
                      reg2099} ?
                  $signed($unsigned(reg2140)) : reg2120));
              reg2148 = (($unsigned($signed($signed(forvar2143))) + wire1999[(1'h1):(1'h0)]) != {(^~((reg2140 ?
                          forvar2116 : reg2136) ?
                      forvar2133 : (^forvar2100)))});
              reg2149 <= (reg2110 + (&$unsigned(reg2119[(2'h2):(1'h0)])));
              reg2150 <= reg2132[(3'h4):(2'h2)];
            end
          reg2151 <= reg2112;
          reg2152 = ($signed((($signed(wire1932) != $unsigned(reg2137)) ^ (wire1934 ?
              $signed(reg2141) : (reg2117 ?
                  (7'h43) : (8'hbf))))) && (^~(~$signed((reg2135 ?
              reg2108 : reg2138)))));
        end
    end
  assign wire2153 = ($signed((($unsigned(reg2142) ?
                            {wire2129,
                                reg2150} : (+(8'hb4))) ^~ $signed((-wire1934)))) ?
                        ($signed(((~^wire2104) ?
                            reg2108[(3'h6):(3'h6)] : $unsigned(reg2144))) * $signed(($signed(wire2129) ?
                            reg2115[(4'hf):(4'ha)] : {wire2130,
                                forvar2146}))) : forvar2146);
  always
    @(posedge clk) begin
      for (forvar2154 = (1'h0); (forvar2154 < (2'h3)); forvar2154 = (forvar2154 + (1'h1)))
        begin
          reg2155 <= ({reg2128[(3'h5):(3'h4)],
                  $unsigned((~reg2103[(4'he):(4'hc)]))} ?
              (($signed((forvar2109 ^~ reg2141)) ^~ reg2147[(4'h8):(1'h1)]) >> $signed(((reg2106 ?
                  forvar2133 : forvar2154) * (reg2124 - reg2144)))) : reg2137[(3'h4):(1'h0)]);
          reg2156 <= ({$unsigned(reg2136[(3'h4):(2'h2)]),
              wire2127} + reg2103[(5'h10):(4'he)]);
        end
      reg2157 = (~^{reg2128[(3'h6):(1'h1)],
          $unsigned(wire1934[(3'h6):(3'h4)])});
      reg2158 = $signed(($signed(((wire1934 ? reg2120 : (7'h40)) ?
          ((8'hb9) << forvar2109) : forvar2133[(3'h7):(3'h6)])) ^ {(8'hb3)}));
      reg2159 <= wire2095;
      reg2160 <= {$unsigned((reg2099[(1'h0):(1'h0)] <<< $signed({reg2152,
              (7'h44)}))),
          reg2119};
    end
  assign wire2161 = {{reg2119, {$unsigned((~&wire1936)), (^forvar2098)}}};
  assign wire2162 = $signed((~^$signed($unsigned((wire2161 ^~ wire1999)))));
  always
    @(posedge clk) begin
      reg2163 <= (8'h9e);
      reg2164 <= $unsigned(reg2126);
      for (forvar2165 = (1'h0); (forvar2165 < (3'h4)); forvar2165 = (forvar2165 + (1'h1)))
        begin
          reg2166 <= ($signed(reg2126[(1'h0):(1'h0)]) ~^ (+(|reg2097)));
          reg2167 = reg2158[(3'h5):(1'h1)];
          reg2168 <= (((($signed(reg2152) ?
                  reg2135[(2'h2):(1'h0)] : $unsigned(reg2118)) << ((!wire1931) != reg2145[(4'hd):(2'h2)])) ?
              reg2103 : $signed(reg2097[(2'h3):(1'h1)])) >= reg2155[(4'hd):(4'h9)]);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2002
#( parameter param2094 = ((8'ha6) >= (~((((8'haf) ? (8'hbd) : (8'ha1)) ? ((8'ha2) ? (7'h43) : (7'h41)) : ((8'hba) ? (8'h9c) : (8'ha0))) == (~&(8'h9c))))) )
(y, clk, wire2006, wire2005, wire2004, wire2003);
  output wire [(32'h41f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire2006;
  input wire signed [(5'h15):(1'h0)] wire2005;
  input wire signed [(5'h12):(1'h0)] wire2004;
  input wire signed [(2'h3):(1'h0)] wire2003;
  wire signed [(5'h10):(1'h0)] wire2093;
  reg [(3'h4):(1'h0)] reg2092 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2091 = (1'h0);
  reg [(2'h3):(1'h0)] reg2090 = (1'h0);
  reg [(5'h11):(1'h0)] reg2089 = (1'h0);
  reg [(4'hd):(1'h0)] reg2088 = (1'h0);
  reg [(2'h3):(1'h0)] reg2087 = (1'h0);
  reg [(4'hd):(1'h0)] reg2086 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2085 = (1'h0);
  reg [(4'ha):(1'h0)] reg2084 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2083 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2082 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2081 = (1'h0);
  reg [(4'hd):(1'h0)] reg2080 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2079 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2078 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2077 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2076 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2075 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2074 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire2073;
  reg [(3'h7):(1'h0)] reg2072 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2071 = (1'h0);
  reg [(3'h5):(1'h0)] reg2070 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2069 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire2068;
  wire signed [(5'h13):(1'h0)] wire2067;
  reg [(4'h9):(1'h0)] reg2066 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2065 = (1'h0);
  reg [(3'h6):(1'h0)] reg2064 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2063 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2062 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2061 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire2060;
  reg [(3'h7):(1'h0)] reg2059 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2058 = (1'h0);
  reg [(3'h5):(1'h0)] reg2057 = (1'h0);
  reg [(5'h13):(1'h0)] reg2056 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2055 = (1'h0);
  reg [(5'h11):(1'h0)] reg2054 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2053 = (1'h0);
  reg [(5'h10):(1'h0)] reg2052 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar2051 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2050 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2049 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2048 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2047 = (1'h0);
  reg [(3'h4):(1'h0)] reg2046 = (1'h0);
  reg [(4'h8):(1'h0)] reg2045 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2044 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2043 = (1'h0);
  reg [(4'hc):(1'h0)] reg2042 = (1'h0);
  reg [(2'h2):(1'h0)] reg2041 = (1'h0);
  reg [(3'h6):(1'h0)] reg2040 = (1'h0);
  reg [(5'h14):(1'h0)] reg2039 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2038 = (1'h0);
  reg [(5'h15):(1'h0)] reg2037 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2036 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2035 = (1'h0);
  reg [(4'hc):(1'h0)] reg2034 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2033 = (1'h0);
  reg [(4'hd):(1'h0)] reg2032 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2031 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2030 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2029 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2028 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2027 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2026 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2025 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2024 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2023 = (1'h0);
  reg [(4'ha):(1'h0)] reg2022 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2021 = (1'h0);
  reg [(4'he):(1'h0)] reg2020 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2019 = (1'h0);
  reg [(4'hb):(1'h0)] reg2018 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2017 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2016 = (1'h0);
  reg [(3'h6):(1'h0)] reg2015 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire2014;
  reg [(4'h8):(1'h0)] reg2013 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2012 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2011 = (1'h0);
  reg [(5'h10):(1'h0)] reg2010 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2009 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2008 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2007 = (1'h0);
  assign y = {wire2093,
                 reg2092,
                 reg2091,
                 reg2090,
                 reg2089,
                 reg2088,
                 reg2087,
                 reg2086,
                 reg2085,
                 reg2084,
                 reg2083,
                 reg2082,
                 reg2081,
                 reg2080,
                 reg2079,
                 reg2078,
                 reg2077,
                 forvar2076,
                 reg2075,
                 forvar2074,
                 wire2073,
                 reg2072,
                 reg2071,
                 reg2070,
                 reg2069,
                 wire2068,
                 wire2067,
                 reg2066,
                 reg2065,
                 reg2064,
                 reg2063,
                 reg2062,
                 forvar2061,
                 wire2060,
                 reg2059,
                 reg2058,
                 reg2057,
                 reg2056,
                 reg2055,
                 reg2054,
                 reg2053,
                 reg2052,
                 forvar2051,
                 reg2050,
                 forvar2049,
                 reg2048,
                 reg2047,
                 reg2046,
                 reg2045,
                 reg2044,
                 reg2043,
                 reg2042,
                 reg2041,
                 reg2040,
                 reg2039,
                 reg2038,
                 reg2037,
                 forvar2036,
                 reg2035,
                 reg2034,
                 reg2033,
                 reg2032,
                 reg2031,
                 forvar2030,
                 reg2029,
                 reg2028,
                 reg2027,
                 reg2026,
                 reg2025,
                 reg2024,
                 forvar2023,
                 reg2022,
                 forvar2021,
                 reg2020,
                 reg2019,
                 reg2018,
                 reg2017,
                 reg2016,
                 reg2015,
                 wire2014,
                 reg2013,
                 forvar2012,
                 reg2011,
                 reg2010,
                 reg2009,
                 forvar2008,
                 reg2007,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg2007 <= $unsigned({wire2003});
    end
  always
    @(posedge clk) begin
      for (forvar2008 = (1'h0); (forvar2008 < (2'h3)); forvar2008 = (forvar2008 + (1'h1)))
        begin
          reg2009 <= wire2005[(4'ha):(4'h9)];
        end
      reg2010 <= wire2004;
      reg2011 <= (($signed(reg2010[(4'hb):(1'h0)]) ^~ {$unsigned($signed((8'h9f))),
              (wire2005[(4'h8):(3'h6)] ? (!forvar2008) : $signed(wire2004))}) ?
          (~(8'ha2)) : wire2003);
      for (forvar2012 = (1'h0); (forvar2012 < (1'h0)); forvar2012 = (forvar2012 + (1'h1)))
        begin
          reg2013 <= $unsigned(reg2010[(4'hb):(3'h6)]);
        end
    end
  assign wire2014 = wire2004[(4'hf):(4'h9)];
  always
    @(posedge clk) begin
      reg2015 <= (^~(~|($unsigned((-reg2013)) || ($unsigned(wire2006) << (reg2013 >= reg2010)))));
      reg2016 = reg2010[(4'h9):(1'h1)];
      reg2017 <= ($unsigned(reg2016[(3'h4):(3'h4)]) ^ reg2009[(3'h6):(2'h3)]);
    end
  always
    @(posedge clk) begin
      reg2018 <= (((reg2011[(4'h9):(3'h7)] ?
                  ((reg2009 <= wire2014) ?
                      reg2011 : {forvar2012}) : $signed({wire2004, (8'hba)})) ?
              ($signed((^forvar2008)) && $unsigned((reg2017 ^ reg2010))) : wire2003) ?
          $unsigned($unsigned($signed((reg2010 < reg2007)))) : reg2010);
    end
  always
    @(posedge clk) begin
      reg2019 <= ((^reg2011[(3'h4):(2'h2)]) ^~ (^~reg2009[(2'h2):(1'h0)]));
      reg2020 <= (reg2019[(4'h9):(1'h1)] < {($unsigned(wire2014[(3'h6):(3'h5)]) ?
              {(+wire2014), (wire2014 < reg2015)} : wire2004),
          $unsigned(forvar2012)});
      for (forvar2021 = (1'h0); (forvar2021 < (3'h4)); forvar2021 = (forvar2021 + (1'h1)))
        begin
          reg2022 = ((({(wire2005 <<< wire2003), reg2019} ?
                  (!(forvar2012 ^~ reg2016)) : (|{reg2010,
                      forvar2012})) - wire2003) ?
              {$unsigned(((~wire2005) ^~ $unsigned(reg2019)))} : reg2009);
          for (forvar2023 = (1'h0); (forvar2023 < (1'h0)); forvar2023 = (forvar2023 + (1'h1)))
            begin
              reg2024 <= (forvar2023 ~^ ((((7'h43) ?
                          $signed(reg2010) : (reg2020 ?
                              forvar2021 : forvar2021)) ?
                      wire2003[(1'h0):(1'h0)] : {(8'h9f),
                          reg2015[(2'h3):(2'h3)]}) ?
                  $unsigned(($unsigned(reg2007) + {reg2015})) : (~^$unsigned(wire2014))));
              reg2025 <= (({(8'h9e),
                          ((forvar2012 >> reg2010) ?
                              $unsigned(reg2007) : (^forvar2008))} ?
                      {(8'hab)} : $signed(($unsigned(forvar2023) | (+reg2010)))) ?
                  ((reg2015 <<< forvar2008[(2'h3):(2'h2)]) ~^ (($unsigned(forvar2021) + (wire2005 ~^ forvar2021)) ^~ ($signed(wire2014) && reg2011))) : reg2018);
              reg2026 = (($unsigned($unsigned((reg2024 ?
                      forvar2021 : wire2006))) >>> $signed(reg2011)) ?
                  $unsigned(reg2024) : $signed($signed({(^~(8'hbf))})));
              reg2027 <= reg2010[(3'h5):(2'h3)];
              reg2028 <= (({((reg2022 ~^ (7'h42)) ?
                          $signed((8'hab)) : (wire2004 + wire2014)),
                      (&$unsigned(reg2007))} + reg2015) ?
                  (^reg2009[(3'h7):(3'h6)]) : ($unsigned(reg2016) ^ reg2025));
            end
          reg2029 <= (reg2015 || reg2013[(2'h3):(2'h2)]);
          for (forvar2030 = (1'h0); (forvar2030 < (3'h4)); forvar2030 = (forvar2030 + (1'h1)))
            begin
              reg2031 <= reg2013;
              reg2032 <= {$signed(reg2028[(4'h9):(2'h3)])};
              reg2033 <= $unsigned(reg2016);
              reg2034 <= ((!((~|(~reg2020)) == {wire2014, wire2004})) ?
                  ((reg2026 ? reg2028 : $unsigned($unsigned((8'hbd)))) ?
                      $unsigned((^$unsigned(reg2011))) : $unsigned(((reg2017 ?
                          forvar2008 : (8'ha5)) | reg2020))) : reg2018[(2'h3):(2'h3)]);
              reg2035 <= $signed(forvar2023[(4'hf):(4'hc)]);
            end
          for (forvar2036 = (1'h0); (forvar2036 < (3'h4)); forvar2036 = (forvar2036 + (1'h1)))
            begin
              reg2037 <= (+$signed($signed(($signed(reg2032) ?
                  (!reg2024) : ((8'hb8) << reg2027)))));
            end
        end
      reg2038 <= ((forvar2008[(3'h6):(2'h2)] ?
          forvar2021 : (~^$unsigned((8'hb5)))) && (8'ha9));
      reg2039 <= forvar2030[(5'h11):(4'hf)];
    end
  always
    @(posedge clk) begin
      reg2040 <= $unsigned($unsigned(($unsigned(reg2024[(3'h6):(1'h1)]) ?
          (~|(^reg2022)) : $unsigned({wire2005, reg2034}))));
      reg2041 = reg2022;
      reg2042 <= ((|forvar2008) ?
          (($signed((&(8'hab))) ?
              {$unsigned(forvar2008),
                  forvar2036} : $signed((^~(8'had)))) | $unsigned(reg2040)) : reg2009[(2'h3):(1'h1)]);
      reg2043 = wire2006;
      reg2044 <= ($signed(forvar2008[(4'hc):(3'h5)]) ?
          $unsigned($unsigned((-$signed(reg2019)))) : $unsigned((+reg2025[(3'h4):(2'h2)])));
    end
  always
    @(posedge clk) begin
      reg2045 <= $unsigned((8'ha7));
      reg2046 <= $unsigned($unsigned((forvar2036 ?
          (~&((8'h9f) > reg2045)) : {(~^reg2028)})));
      reg2047 = ((+($unsigned($signed(reg2037)) ?
          reg2024[(4'h8):(2'h3)] : ((~^reg2035) <<< $unsigned(reg2025)))) ~^ $signed(reg2018[(4'ha):(2'h2)]));
    end
  always
    @(posedge clk) begin
      reg2048 <= reg2039[(1'h0):(1'h0)];
      for (forvar2049 = (1'h0); (forvar2049 < (3'h4)); forvar2049 = (forvar2049 + (1'h1)))
        begin
          reg2050 <= reg2040;
          for (forvar2051 = (1'h0); (forvar2051 < (1'h0)); forvar2051 = (forvar2051 + (1'h1)))
            begin
              reg2052 <= ((({reg2041} == $signed(reg2041[(1'h1):(1'h1)])) ?
                      reg2033 : (wire2004[(3'h7):(2'h3)] < {wire2006,
                          $signed((8'hbc))})) ?
                  ((!(((8'hbf) ?
                      (8'had) : forvar2021) > (~^(8'ha3)))) ^ reg2039[(4'he):(1'h0)]) : (reg2028 ?
                      (8'h9d) : reg2039));
              reg2053 <= reg2016[(3'h4):(1'h1)];
              reg2054 = $signed($signed((|$unsigned((~&reg2018)))));
              reg2055 <= reg2019[(3'h6):(2'h2)];
              reg2056 <= {($signed(reg2028[(4'h8):(3'h6)]) ?
                      $unsigned(($unsigned((7'h44)) ?
                          $signed(reg2010) : $signed((8'hbf)))) : {((reg2042 ?
                                  wire2006 : reg2047) ?
                              $unsigned(reg2053) : $unsigned(reg2016))})};
            end
        end
      reg2057 <= wire2005;
      reg2058 <= (reg2040[(1'h1):(1'h1)] ?
          $signed(reg2041) : reg2042[(4'hc):(4'h8)]);
      reg2059 <= reg2053[(4'ha):(2'h2)];
    end
  assign wire2060 = reg2038[(4'ha):(3'h5)];
  always
    @(posedge clk) begin
      for (forvar2061 = (1'h0); (forvar2061 < (2'h3)); forvar2061 = (forvar2061 + (1'h1)))
        begin
          reg2062 = (reg2019[(4'h8):(2'h3)] ?
              $unsigned((reg2016 ?
                  $unsigned(reg2042) : forvar2023[(4'ha):(1'h0)])) : (+((!$signed(reg2029)) < {wire2060[(2'h3):(2'h2)]})));
          reg2063 <= reg2015[(1'h1):(1'h1)];
          reg2064 <= (+$signed((8'hae)));
        end
      reg2065 = {(((|(8'hb7)) ?
                  (((8'hb3) ?
                      reg2064 : reg2054) * wire2014[(3'h5):(3'h4)]) : $unsigned((reg2064 | reg2038))) ?
              (8'hbb) : ($unsigned(reg2057[(1'h0):(1'h0)]) <= $signed(reg2017))),
          (reg2015[(2'h3):(2'h2)] ? reg2040[(2'h2):(1'h1)] : (8'ha7))};
      reg2066 <= reg2035;
    end
  assign wire2067 = {forvar2036[(1'h0):(1'h0)]};
  assign wire2068 = reg2031[(4'he):(3'h6)];
  always
    @(posedge clk) begin
      reg2069 <= (reg2040 ?
          $signed($signed(({reg2056} ?
              (wire2067 << reg2034) : reg2024[(3'h5):(3'h4)]))) : ($signed($signed((reg2015 >> reg2044))) > (reg2052 ?
              $unsigned(reg2032[(2'h2):(1'h1)]) : $unsigned((+forvar2061)))));
      reg2070 <= $signed(reg2048);
      reg2071 = $unsigned((8'hbf));
      reg2072 <= (reg2054[(4'hd):(4'hd)] ?
          reg2052[(4'hb):(3'h6)] : {(((reg2063 ? reg2046 : reg2026) ?
                      $signed(reg2032) : reg2025) ?
                  (((8'ha1) ?
                      reg2056 : (8'hb5)) >= reg2054) : $signed((wire2068 << reg2053)))});
    end
  assign wire2073 = ($unsigned($unsigned(reg2044[(4'h8):(3'h7)])) ?
                        ((^~($signed(reg2071) ?
                            reg2058 : $unsigned(reg2007))) * (-reg2032)) : $unsigned($unsigned($unsigned({wire2014}))));
  always
    @(posedge clk) begin
      for (forvar2074 = (1'h0); (forvar2074 < (1'h0)); forvar2074 = (forvar2074 + (1'h1)))
        begin
          reg2075 <= ($signed((((+(8'had)) != {wire2006}) ?
              ({(7'h44)} > (!reg2070)) : (reg2043 ?
                  (^reg2009) : reg2066[(4'h8):(3'h4)]))) + $signed((+$unsigned({(8'haf),
              wire2068}))));
          for (forvar2076 = (1'h0); (forvar2076 < (1'h0)); forvar2076 = (forvar2076 + (1'h1)))
            begin
              reg2077 <= {(&(reg2066 ^ {(+reg2047), reg2009[(3'h5):(3'h4)]})),
                  $signed($signed(reg2024[(1'h1):(1'h1)]))};
              reg2078 <= reg2048[(3'h7):(3'h5)];
              reg2079 <= {((forvar2008 ?
                          {$signed(reg2032),
                              reg2077[(3'h5):(2'h2)]} : ($signed(reg2013) == (reg2075 ?
                              (7'h43) : reg2007))) ?
                      $signed(reg2039) : ($unsigned((reg2053 * wire2073)) ?
                          ((reg2078 ?
                              forvar2030 : (8'h9e)) == $unsigned(reg2072)) : (!(8'hb0))))};
            end
          reg2080 <= $signed($signed(wire2068));
          reg2081 = (reg2034[(1'h0):(1'h0)] ?
              $unsigned({(wire2003 ?
                      reg2037[(3'h7):(1'h0)] : wire2067)}) : (&forvar2036));
        end
      reg2082 <= reg2081[(4'hb):(3'h7)];
      reg2083 <= reg2045[(3'h7):(3'h5)];
      reg2084 <= $unsigned(((8'had) ?
          reg2029 : (($unsigned((7'h44)) | reg2071[(4'ha):(4'h8)]) ?
              $unsigned({reg2024}) : reg2053)));
      reg2085 <= ({(($unsigned(reg2057) << $unsigned(reg2070)) ?
                  reg2027[(2'h2):(2'h2)] : {$unsigned(reg2026),
                      $unsigned(reg2024)})} ?
          reg2034 : (-(8'hb9)));
    end
  always
    @(posedge clk) begin
      reg2086 = (8'hb5);
      reg2087 = (($signed($signed((8'hbb))) - {$unsigned(forvar2049),
          ($signed(wire2073) >>> reg2027)}) || {((!(reg2065 <<< reg2069)) - (+reg2007[(4'ha):(2'h2)])),
          $unsigned($signed($signed(reg2026)))});
    end
  always
    @(posedge clk) begin
      reg2088 <= (~|(($signed($unsigned(reg2022)) == {$unsigned((8'ha5))}) ?
          (!reg2054) : {((8'ha7) ?
                  (reg2065 + reg2056) : reg2077[(4'h9):(3'h4)])}));
      reg2089 = (-reg2046[(3'h4):(3'h4)]);
      reg2090 <= $signed(reg2089);
      reg2091 <= reg2066[(3'h5):(3'h4)];
      reg2092 <= $unsigned($signed(($signed(reg2085[(1'h0):(1'h0)]) & $signed((reg2087 > (8'hb9))))));
    end
  assign wire2093 = $signed((^(~$unsigned($unsigned(reg2069)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1937  (y, clk, wire1941, wire1940, wire1939, wire1938);
  output wire [(32'h247):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire1941;
  input wire signed [(3'h7):(1'h0)] wire1940;
  input wire signed [(3'h7):(1'h0)] wire1939;
  input wire signed [(5'h14):(1'h0)] wire1938;
  wire signed [(4'hf):(1'h0)] wire1995;
  wire [(4'h8):(1'h0)] wire1994;
  reg [(4'hb):(1'h0)] reg1993 = (1'h0);
  reg [(3'h5):(1'h0)] reg1992 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1991 = (1'h0);
  reg [(4'hf):(1'h0)] reg1990 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire1989;
  wire signed [(2'h3):(1'h0)] wire1988;
  reg signed [(2'h2):(1'h0)] reg1987 = (1'h0);
  reg [(5'h10):(1'h0)] reg1986 = (1'h0);
  reg [(4'ha):(1'h0)] reg1985 = (1'h0);
  reg [(3'h6):(1'h0)] reg1984 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1983 = (1'h0);
  reg [(3'h6):(1'h0)] reg1982 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1981 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1980 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1979 = (1'h0);
  wire [(4'h8):(1'h0)] wire1978;
  wire [(3'h7):(1'h0)] wire1977;
  reg [(4'he):(1'h0)] reg1976 = (1'h0);
  reg [(4'h8):(1'h0)] reg1975 = (1'h0);
  reg [(3'h4):(1'h0)] reg1974 = (1'h0);
  wire [(2'h3):(1'h0)] wire1973;
  wire [(4'hd):(1'h0)] wire1972;
  reg signed [(4'h9):(1'h0)] reg1971 = (1'h0);
  reg [(5'h12):(1'h0)] reg1970 = (1'h0);
  reg [(4'hd):(1'h0)] reg1969 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1968 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1967 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1966 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1965 = (1'h0);
  reg [(3'h4):(1'h0)] reg1964 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1963 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1962 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1961 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1960 = (1'h0);
  reg [(3'h7):(1'h0)] reg1959 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1958 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire1957;
  wire signed [(5'h11):(1'h0)] wire1956;
  wire [(2'h3):(1'h0)] wire1955;
  reg [(5'h15):(1'h0)] reg1954 = (1'h0);
  reg [(5'h12):(1'h0)] reg1953 = (1'h0);
  reg [(5'h15):(1'h0)] reg1952 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1951 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1950 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1949 = (1'h0);
  wire [(3'h4):(1'h0)] wire1948;
  reg [(4'he):(1'h0)] reg1947 = (1'h0);
  reg [(3'h5):(1'h0)] reg1946 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1945 = (1'h0);
  reg [(4'h9):(1'h0)] reg1944 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1943 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1942 = (1'h0);
  assign y = {wire1995,
                 wire1994,
                 reg1993,
                 reg1992,
                 reg1991,
                 reg1990,
                 wire1989,
                 wire1988,
                 reg1987,
                 reg1986,
                 reg1985,
                 reg1984,
                 forvar1983,
                 reg1982,
                 reg1981,
                 reg1980,
                 reg1979,
                 wire1978,
                 wire1977,
                 reg1976,
                 reg1975,
                 reg1974,
                 wire1973,
                 wire1972,
                 reg1971,
                 reg1970,
                 reg1969,
                 reg1968,
                 reg1967,
                 reg1966,
                 forvar1965,
                 reg1964,
                 reg1963,
                 reg1962,
                 forvar1961,
                 reg1960,
                 reg1959,
                 reg1958,
                 wire1957,
                 wire1956,
                 wire1955,
                 reg1954,
                 reg1953,
                 reg1952,
                 reg1951,
                 reg1950,
                 forvar1949,
                 wire1948,
                 reg1947,
                 reg1946,
                 reg1945,
                 reg1944,
                 forvar1943,
                 reg1942,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1942 <= $unsigned(({{{wire1939, wire1940}}, wire1940} < wire1940));
      for (forvar1943 = (1'h0); (forvar1943 < (1'h1)); forvar1943 = (forvar1943 + (1'h1)))
        begin
          reg1944 <= ({(~&($unsigned(reg1942) ^~ {(8'hbd)}))} <= $unsigned((^($signed(wire1939) & (7'h42)))));
        end
      reg1945 <= {$signed(($unsigned($signed(reg1942)) ?
              (((8'hac) ?
                  wire1938 : wire1939) >>> (wire1940 <<< forvar1943)) : (forvar1943 ?
                  forvar1943[(1'h0):(1'h0)] : $unsigned(wire1940))))};
      reg1946 <= (&(wire1938[(1'h1):(1'h0)] <<< $signed($signed($signed(wire1941)))));
      reg1947 = wire1941[(2'h2):(1'h1)];
    end
  assign wire1948 = ($signed((wire1938[(4'h9):(3'h5)] && ($signed(wire1938) ?
                            $signed((8'h9e)) : $signed(reg1947)))) ?
                        (8'haf) : $signed($signed($signed((7'h43)))));
  always
    @(posedge clk) begin
      for (forvar1949 = (1'h0); (forvar1949 < (3'h4)); forvar1949 = (forvar1949 + (1'h1)))
        begin
          reg1950 <= $signed((($unsigned({wire1939}) ?
                  ((reg1946 ?
                      reg1946 : forvar1949) && wire1940[(3'h5):(2'h3)]) : (8'hab)) ?
              {reg1944[(4'h8):(2'h3)]} : $unsigned(((forvar1943 | reg1947) ?
                  wire1938 : (+(8'hb2))))));
        end
      reg1951 <= ($unsigned((^~((|wire1948) * $unsigned(reg1950)))) << (^($signed(reg1945[(3'h4):(2'h3)]) ?
          (8'hbf) : (8'hb3))));
      reg1952 <= $signed((($signed({(8'ha7), wire1938}) ?
          (+wire1938) : ({(8'hb4)} + reg1944)) | ($unsigned((reg1950 == (8'hb3))) * (!$unsigned(reg1946)))));
      reg1953 <= reg1945[(3'h6):(3'h4)];
      reg1954 <= wire1948;
    end
  assign wire1955 = reg1950;
  assign wire1956 = wire1938;
  assign wire1957 = (((+wire1948) ?
                        wire1955[(1'h0):(1'h0)] : ($signed($signed(wire1941)) | (reg1950[(4'hd):(3'h7)] ^ {wire1939,
                            wire1940}))) + $signed((8'ha9)));
  always
    @(posedge clk) begin
      reg1958 = {$unsigned({(7'h40)})};
      reg1959 <= (forvar1943 ?
          $unsigned((reg1944[(4'h9):(3'h7)] > $unsigned((wire1939 ?
              wire1948 : forvar1943)))) : ({(|(wire1938 ?
                      wire1938 : wire1957))} ?
              forvar1943 : ($signed((&reg1952)) > (~forvar1949[(5'h10):(1'h0)]))));
      reg1960 <= (8'ha5);
      for (forvar1961 = (1'h0); (forvar1961 < (2'h2)); forvar1961 = (forvar1961 + (1'h1)))
        begin
          reg1962 = $unsigned((8'hb5));
          reg1963 = $unsigned((wire1941[(1'h1):(1'h0)] ?
              {(8'hb4)} : (|forvar1949[(5'h14):(5'h10)])));
          reg1964 = $unsigned({reg1960, wire1948});
          for (forvar1965 = (1'h0); (forvar1965 < (3'h4)); forvar1965 = (forvar1965 + (1'h1)))
            begin
              reg1966 <= reg1954[(5'h14):(5'h11)];
              reg1967 <= $signed($unsigned(reg1942[(3'h4):(1'h1)]));
              reg1968 <= reg1945;
              reg1969 <= (~^$unsigned(((!(~wire1957)) ?
                  ($signed((8'hb8)) ?
                      (wire1955 >>> (8'ha0)) : (8'hbc)) : ((forvar1943 ^ wire1938) ?
                      $unsigned((7'h43)) : reg1951[(1'h0):(1'h0)]))));
              reg1970 = (|(-$signed($unsigned(wire1941[(2'h3):(1'h0)]))));
            end
          reg1971 <= wire1939;
        end
    end
  assign wire1972 = (+(8'h9e));
  assign wire1973 = $signed(((~forvar1965[(1'h0):(1'h0)]) ?
                        reg1952[(4'hf):(3'h4)] : (reg1946[(3'h5):(1'h0)] && (reg1954[(3'h4):(3'h4)] || reg1964[(1'h0):(1'h0)]))));
  always
    @(posedge clk) begin
      reg1974 = ((-$unsigned((wire1938[(2'h2):(1'h0)] <<< forvar1949))) ?
          ($signed(reg1947) <= $signed((reg1944 ?
              $unsigned((8'ha0)) : $unsigned((8'hb3))))) : reg1966);
      reg1975 <= $signed($unsigned((reg1967[(4'ha):(2'h2)] ?
          wire1938 : $signed($unsigned(wire1972)))));
      reg1976 = $signed(($signed(($signed(reg1954) ?
          {reg1954} : ((8'ha1) <<< wire1948))) | (~|$unsigned($signed(reg1974)))));
    end
  assign wire1977 = reg1960[(3'h4):(1'h0)];
  assign wire1978 = (-{$unsigned(wire1956),
                        $unsigned((wire1973[(2'h2):(1'h0)] ?
                            forvar1961[(1'h1):(1'h0)] : (reg1946 ?
                                (8'hb7) : reg1969)))});
  always
    @(posedge clk) begin
      reg1979 = wire1973;
      reg1980 <= $signed(wire1941[(1'h1):(1'h0)]);
      reg1981 <= wire1977;
      reg1982 = (((reg1953 ? $signed((^reg1968)) : reg1981[(4'hc):(4'ha)]) ?
              $signed(reg1951) : (reg1952 && wire1972[(3'h5):(1'h1)])) ?
          {$unsigned($signed(reg1964[(2'h3):(1'h1)])),
              {((wire1956 ? reg1962 : (8'hb2)) ?
                      (reg1969 >>> reg1980) : (^(8'ha3)))}} : reg1974[(2'h3):(2'h3)]);
      for (forvar1983 = (1'h0); (forvar1983 < (3'h4)); forvar1983 = (forvar1983 + (1'h1)))
        begin
          reg1984 <= reg1959;
          reg1985 <= $unsigned({$unsigned(($signed(wire1938) + forvar1949))});
          reg1986 = (reg1947[(2'h2):(2'h2)] << (-$signed(($signed(wire1972) && $unsigned(forvar1965)))));
          reg1987 <= (^~$signed($unsigned(reg1958[(4'h8):(4'h8)])));
        end
    end
  assign wire1988 = wire1972[(1'h1):(1'h1)];
  assign wire1989 = ($signed({reg1950,
                        ((^reg1953) <<< (reg1970 == reg1979))}) | (8'hbd));
  always
    @(posedge clk) begin
      reg1990 = (($signed((!reg1960[(3'h7):(3'h5)])) ?
          reg1942[(4'h9):(1'h0)] : (~(&$unsigned(reg1969)))) & (~&reg1962));
      reg1991 <= ($unsigned(($unsigned($unsigned(reg1951)) ?
          (~^reg1990[(2'h2):(2'h2)]) : ($unsigned(wire1941) <<< reg1969))) >>> $signed($signed($unsigned(reg1963))));
      reg1992 <= reg1969;
      reg1993 <= {wire1948[(1'h0):(1'h0)]};
    end
  assign wire1994 = ({($unsigned($unsigned(wire1940)) ?
                                $signed($unsigned(reg1991)) : wire1977[(2'h2):(1'h0)]),
                            {{(reg1975 ? reg1990 : forvar1949)},
                                $unsigned((reg1976 ? forvar1965 : (8'hb5)))}} ?
                        (-{(-(~reg1991)),
                            (~|$unsigned(reg1993))}) : wire1988[(2'h2):(1'h1)]);
  assign wire1995 = $unsigned($signed(((reg1958[(2'h3):(2'h3)] - reg1963) ~^ (wire1940[(3'h4):(1'h1)] * (&wire1941)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2558
#( parameter param2603 = {((({(8'ha0)} || (^~(8'h9e))) ? {((7'h44) ? (8'hbd) : (8'h9d)), ((8'hb5) ^~ (8'hbd))} : ({(8'hb8)} ? (7'h40) : ((8'hac) ? (7'h42) : (8'h9d)))) ? (~&{((8'ha5) >= (8'had)), ((8'h9e) ? (8'hbb) : (8'hb3))}) : ((^~((8'hb9) >>> (8'ha6))) ? (((8'h9d) >>> (8'hbc)) * (~&(7'h40))) : {(&(8'hab))})), ((8'haa) & {(((8'hb6) && (8'hbc)) ? ((8'ha9) ? (8'hb9) : (7'h43)) : ((7'h42) >>> (8'haf)))})}
, parameter param2604 = param2603 )
(y, clk, wire2563, wire2562, wire2561, wire2560, wire2559);
  output wire [(32'h188):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire2563;
  input wire [(4'h9):(1'h0)] wire2562;
  input wire signed [(5'h13):(1'h0)] wire2561;
  input wire [(5'h14):(1'h0)] wire2560;
  input wire [(4'hd):(1'h0)] wire2559;
  reg signed [(4'hc):(1'h0)] reg2602 = (1'h0);
  reg [(4'ha):(1'h0)] reg2601 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire2600;
  wire [(3'h4):(1'h0)] wire2599;
  reg signed [(4'hb):(1'h0)] reg2598 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2597 = (1'h0);
  reg [(3'h6):(1'h0)] reg2596 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2595 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2594 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2593 = (1'h0);
  reg [(4'ha):(1'h0)] reg2592 = (1'h0);
  reg [(2'h3):(1'h0)] reg2591 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2590 = (1'h0);
  reg [(3'h4):(1'h0)] reg2589 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2588 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2587 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2586 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2585 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2584 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2583 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2582 = (1'h0);
  reg [(5'h15):(1'h0)] reg2581 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2580 = (1'h0);
  reg [(4'hb):(1'h0)] reg2579 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2578 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2577 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2576 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2575 = (1'h0);
  reg [(2'h3):(1'h0)] reg2574 = (1'h0);
  reg [(4'hb):(1'h0)] reg2573 = (1'h0);
  reg [(5'h12):(1'h0)] reg2572 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2571 = (1'h0);
  reg [(2'h3):(1'h0)] reg2570 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2569 = (1'h0);
  reg [(3'h5):(1'h0)] reg2568 = (1'h0);
  reg [(4'h9):(1'h0)] reg2567 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire2566;
  wire [(5'h13):(1'h0)] wire2565;
  wire [(3'h7):(1'h0)] wire2564;
  assign y = {reg2602,
                 reg2601,
                 wire2600,
                 wire2599,
                 reg2598,
                 reg2597,
                 reg2596,
                 reg2595,
                 reg2594,
                 forvar2593,
                 reg2592,
                 reg2591,
                 reg2590,
                 reg2589,
                 forvar2588,
                 reg2587,
                 reg2586,
                 forvar2585,
                 reg2584,
                 forvar2583,
                 reg2582,
                 reg2581,
                 reg2580,
                 reg2579,
                 forvar2578,
                 forvar2577,
                 reg2576,
                 reg2575,
                 reg2574,
                 reg2573,
                 reg2572,
                 forvar2571,
                 reg2570,
                 forvar2569,
                 reg2568,
                 reg2567,
                 wire2566,
                 wire2565,
                 wire2564,
                 (1'h0)};
  assign wire2564 = (wire2563[(1'h0):(1'h0)] ?
                        (wire2562 ?
                            $signed($unsigned((8'ha2))) : ($unsigned((wire2559 ?
                                    wire2560 : wire2561)) ?
                                (~(~wire2559)) : $unsigned((wire2563 || wire2559)))) : (({wire2560[(5'h13):(4'hf)],
                                    $unsigned(wire2559)} ?
                                ({wire2562} ?
                                    $unsigned(wire2561) : (-wire2562)) : wire2560) ?
                            $signed(wire2563[(1'h1):(1'h0)]) : $unsigned($unsigned(wire2563))));
  assign wire2565 = $signed(($signed(wire2560[(3'h7):(3'h5)]) >> (~&$signed(wire2563[(2'h3):(2'h2)]))));
  assign wire2566 = (+$unsigned($unsigned(wire2565)));
  always
    @(posedge clk) begin
      reg2567 = wire2562[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg2568 <= {((7'h41) < (&$signed(wire2565[(4'ha):(2'h2)])))};
      for (forvar2569 = (1'h0); (forvar2569 < (2'h2)); forvar2569 = (forvar2569 + (1'h1)))
        begin
          reg2570 <= reg2568;
          for (forvar2571 = (1'h0); (forvar2571 < (1'h1)); forvar2571 = (forvar2571 + (1'h1)))
            begin
              reg2572 = {$signed($signed(reg2568[(3'h5):(1'h0)]))};
              reg2573 = $unsigned({$unsigned(wire2563)});
              reg2574 = (($signed(((reg2572 >>> reg2568) ?
                      {reg2567, (8'hb5)} : (reg2572 ?
                          wire2561 : wire2564))) ^ (($signed((8'hab)) > (~|(8'hb0))) ?
                      ($unsigned(reg2570) >= (reg2572 ?
                          reg2573 : forvar2569)) : ((+wire2561) == $signed(wire2563)))) ?
                  reg2572[(1'h0):(1'h0)] : reg2570[(2'h2):(1'h1)]);
            end
        end
      reg2575 <= $signed((&reg2568));
      reg2576 <= $unsigned({wire2560[(4'hb):(2'h2)]});
    end
  always
    @(posedge clk) begin
      for (forvar2577 = (1'h0); (forvar2577 < (1'h1)); forvar2577 = (forvar2577 + (1'h1)))
        begin
          for (forvar2578 = (1'h0); (forvar2578 < (2'h3)); forvar2578 = (forvar2578 + (1'h1)))
            begin
              reg2579 <= $unsigned((($signed($signed(reg2573)) ?
                  (~^(&reg2575)) : $unsigned($unsigned(reg2574))) ~^ forvar2569));
              reg2580 <= reg2573[(1'h0):(1'h0)];
            end
          reg2581 = {(~&(^~reg2575[(4'h9):(1'h1)])), reg2576[(1'h0):(1'h0)]};
        end
      reg2582 = wire2565;
      for (forvar2583 = (1'h0); (forvar2583 < (2'h3)); forvar2583 = (forvar2583 + (1'h1)))
        begin
          reg2584 <= (8'ha7);
          for (forvar2585 = (1'h0); (forvar2585 < (2'h2)); forvar2585 = (forvar2585 + (1'h1)))
            begin
              reg2586 = reg2581;
            end
          reg2587 <= $signed($signed($unsigned({reg2576[(3'h4):(3'h4)],
              reg2574})));
        end
      for (forvar2588 = (1'h0); (forvar2588 < (2'h2)); forvar2588 = (forvar2588 + (1'h1)))
        begin
          reg2589 <= ($signed((8'haa)) ?
              reg2587 : ((forvar2578 ?
                  ((reg2587 ? reg2586 : reg2568) & ((8'hb9) ?
                      (8'hba) : forvar2571)) : ($unsigned(wire2563) ?
                      (&wire2559) : ((8'hbb) ~^ wire2560))) <<< ((~|(reg2581 ?
                  reg2580 : wire2561)) | $unsigned((wire2561 ?
                  reg2572 : reg2587)))));
          reg2590 <= (wire2564[(3'h6):(2'h3)] ?
              reg2574[(2'h3):(2'h3)] : wire2560);
          reg2591 <= reg2587[(1'h1):(1'h1)];
          reg2592 = $unsigned((forvar2577 < $signed(reg2586)));
          for (forvar2593 = (1'h0); (forvar2593 < (1'h0)); forvar2593 = (forvar2593 + (1'h1)))
            begin
              reg2594 <= $signed((+$unsigned(((+(8'hb4)) ?
                  reg2591 : $signed(forvar2577)))));
              reg2595 = (8'ha2);
              reg2596 <= (reg2567 ?
                  ($signed((reg2586[(3'h7):(3'h5)] ?
                          reg2579[(4'h8):(1'h0)] : forvar2588[(3'h7):(3'h4)])) ?
                      $unsigned(($unsigned(forvar2577) & {wire2565,
                          forvar2585})) : (8'hbf)) : (~^$signed(($signed((8'h9f)) < ((8'had) ?
                      reg2576 : reg2576)))));
              reg2597 <= ($signed(reg2568[(2'h2):(1'h1)]) ~^ wire2560[(4'h9):(1'h1)]);
              reg2598 <= reg2581[(1'h0):(1'h0)];
            end
        end
    end
  assign wire2599 = (^~reg2586[(3'h5):(3'h5)]);
  assign wire2600 = {((reg2579 >>> reg2568) + $unsigned({(~forvar2583)})),
                        $signed((~&$unsigned(wire2599[(2'h2):(1'h0)])))};
  always
    @(posedge clk) begin
      reg2601 <= ((~(!wire2559[(3'h6):(3'h6)])) ?
          $unsigned(($unsigned((~|reg2592)) || reg2595)) : ((reg2570 ?
              $signed($unsigned(reg2586)) : ($unsigned(wire2565) && (~reg2584))) & $unsigned($unsigned((^reg2595)))));
      reg2602 <= (-{$unsigned((((8'hb0) <<< wire2562) & reg2589)),
          (wire2562 | $signed(reg2598[(3'h7):(1'h1)]))});
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2491
#( parameter param2553 = ((((((8'ha2) ? (8'hbc) : (8'hbf)) ? (8'hb4) : (~^(8'hbe))) ? ((8'ha2) >> ((7'h42) & (7'h43))) : (^~(~|(8'hbd)))) & (^~(((8'h9d) ? (8'had) : (8'ha1)) >> {(8'hbe)}))) ? ((({(8'hb5)} >>> ((8'ha5) ? (8'ha3) : (8'ha8))) && ((+(8'ha0)) ? ((8'hb1) ? (8'hbc) : (8'hbb)) : ((7'h44) + (8'hab)))) ? (^~(~|((7'h43) ? (8'hba) : (8'ha7)))) : (((|(7'h42)) < {(8'ha2)}) ? ({(8'ha1), (8'hb6)} | ((8'hbc) ? (7'h43) : (8'ha4))) : (^~((8'hba) ? (8'hb3) : (8'hb9))))) : ((^~(8'ha1)) ^ ({((8'haa) >>> (8'ha4))} ? (^((8'hb6) <= (8'ha7))) : (((7'h40) ? (8'had) : (8'ha5)) ? {(8'ha1)} : (&(8'h9f))))))
, parameter param2554 = (~^(!param2553)) )
(y, clk, wire2496, wire2495, wire2494, wire2493, wire2492);
  output wire [(32'h251):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire2496;
  input wire [(3'h4):(1'h0)] wire2495;
  input wire signed [(4'hf):(1'h0)] wire2494;
  input wire signed [(5'h14):(1'h0)] wire2493;
  input wire [(2'h3):(1'h0)] wire2492;
  reg [(5'h12):(1'h0)] reg2552 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2551 = (1'h0);
  reg [(4'h9):(1'h0)] reg2550 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2549 = (1'h0);
  reg [(3'h4):(1'h0)] reg2548 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2547 = (1'h0);
  reg [(3'h4):(1'h0)] reg2546 = (1'h0);
  reg [(5'h13):(1'h0)] reg2545 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2544 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2543 = (1'h0);
  reg [(5'h13):(1'h0)] reg2542 = (1'h0);
  reg [(3'h5):(1'h0)] reg2541 = (1'h0);
  reg [(4'hd):(1'h0)] reg2540 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2539 = (1'h0);
  reg [(2'h3):(1'h0)] reg2538 = (1'h0);
  reg [(3'h7):(1'h0)] reg2537 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2536 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2535 = (1'h0);
  reg [(5'h12):(1'h0)] reg2534 = (1'h0);
  reg [(4'h8):(1'h0)] reg2533 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2532 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2531 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2530 = (1'h0);
  reg [(3'h4):(1'h0)] reg2529 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2528 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2527 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2526 = (1'h0);
  reg [(2'h2):(1'h0)] reg2525 = (1'h0);
  reg [(5'h15):(1'h0)] reg2524 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2523 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2522 = (1'h0);
  reg [(5'h11):(1'h0)] reg2521 = (1'h0);
  reg [(2'h3):(1'h0)] reg2520 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2519 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2518 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2517 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2516 = (1'h0);
  reg [(5'h11):(1'h0)] reg2515 = (1'h0);
  reg [(5'h14):(1'h0)] reg2514 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2513 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2512 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2511 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2510 = (1'h0);
  reg [(5'h10):(1'h0)] reg2509 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2508 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2507 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire2506;
  wire signed [(4'hc):(1'h0)] wire2505;
  reg signed [(5'h11):(1'h0)] reg2504 = (1'h0);
  reg [(4'h9):(1'h0)] reg2503 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire2502;
  reg [(4'hd):(1'h0)] reg2501 = (1'h0);
  reg [(4'he):(1'h0)] reg2500 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2499 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2498 = (1'h0);
  reg [(2'h2):(1'h0)] reg2497 = (1'h0);
  assign y = {reg2552,
                 reg2551,
                 reg2550,
                 forvar2549,
                 reg2548,
                 reg2547,
                 reg2546,
                 reg2545,
                 reg2544,
                 reg2543,
                 reg2542,
                 reg2541,
                 reg2540,
                 reg2539,
                 reg2538,
                 reg2537,
                 forvar2536,
                 reg2535,
                 reg2534,
                 reg2533,
                 reg2532,
                 reg2531,
                 forvar2530,
                 reg2529,
                 reg2528,
                 forvar2527,
                 reg2526,
                 reg2525,
                 reg2524,
                 reg2523,
                 forvar2522,
                 reg2521,
                 reg2520,
                 forvar2519,
                 reg2518,
                 reg2517,
                 reg2516,
                 reg2515,
                 reg2514,
                 reg2513,
                 reg2512,
                 forvar2511,
                 forvar2510,
                 reg2509,
                 reg2508,
                 forvar2507,
                 wire2506,
                 wire2505,
                 reg2504,
                 reg2503,
                 wire2502,
                 reg2501,
                 reg2500,
                 reg2499,
                 reg2498,
                 reg2497,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg2497 <= ((7'h42) ?
          $unsigned({wire2493,
              wire2494[(3'h4):(2'h3)]}) : (~$signed($unsigned((8'hba)))));
      reg2498 <= wire2494;
      reg2499 <= (~|{wire2495[(2'h3):(2'h3)]});
      if (reg2498[(1'h1):(1'h1)])
        begin
          reg2500 <= $signed(($signed((^~(wire2494 < reg2498))) >= (-wire2493)));
          reg2501 <= reg2497[(1'h1):(1'h1)];
        end
      else
        begin
          reg2500 <= ((|wire2496) ?
              (~$unsigned($unsigned($unsigned((8'ha9))))) : (($signed(((8'ha9) ?
                      wire2493 : wire2493)) ~^ $unsigned((~^reg2501))) ?
                  reg2497[(1'h0):(1'h0)] : reg2499[(3'h7):(3'h7)]));
        end
    end
  assign wire2502 = (~^(-((|(reg2501 | wire2493)) ?
                        ((reg2501 ? (8'hb7) : reg2497) == (wire2494 ?
                            wire2494 : reg2500)) : reg2499[(2'h2):(1'h1)])));
  always
    @(posedge clk) begin
      reg2503 = reg2500[(4'h8):(2'h3)];
      reg2504 <= $signed((wire2502 ~^ {{{wire2494, reg2498}}}));
    end
  assign wire2505 = ((~&(+({wire2492} && (~^wire2492)))) && (wire2493 ?
                        (wire2494[(3'h7):(1'h0)] - ((reg2501 >= reg2501) == $signed(reg2498))) : $unsigned(((reg2504 ?
                            wire2494 : wire2495) ^ wire2492))));
  assign wire2506 = (reg2498 >> wire2493);
  always
    @(posedge clk) begin
      for (forvar2507 = (1'h0); (forvar2507 < (3'h4)); forvar2507 = (forvar2507 + (1'h1)))
        begin
          reg2508 <= $signed({($signed($unsigned((8'ha2))) ?
                  (!reg2499[(3'h5):(3'h5)]) : reg2497[(1'h1):(1'h1)]),
              ((!$unsigned(reg2504)) ?
                  {{wire2506, wire2494},
                      $unsigned((8'hbb))} : (reg2497[(1'h1):(1'h1)] == (8'hba)))});
        end
      reg2509 <= (^~$signed(wire2492));
      for (forvar2510 = (1'h0); (forvar2510 < (2'h2)); forvar2510 = (forvar2510 + (1'h1)))
        begin
          for (forvar2511 = (1'h0); (forvar2511 < (2'h3)); forvar2511 = (forvar2511 + (1'h1)))
            begin
              reg2512 = $signed($signed($unsigned(((wire2496 ?
                      reg2503 : forvar2507) ?
                  (wire2496 | wire2492) : (wire2493 ^~ (8'hbe))))));
              reg2513 = $unsigned({(+$unsigned(reg2499[(1'h0):(1'h0)])),
                  reg2499});
              reg2514 <= forvar2510;
              reg2515 <= reg2499;
              reg2516 <= (8'hb7);
            end
          reg2517 <= (wire2493 >= reg2498[(2'h2):(1'h1)]);
          reg2518 <= (8'hab);
        end
      for (forvar2519 = (1'h0); (forvar2519 < (1'h0)); forvar2519 = (forvar2519 + (1'h1)))
        begin
          reg2520 <= (~reg2518);
        end
    end
  always
    @(posedge clk) begin
      reg2521 <= ($signed($signed($unsigned($unsigned(reg2518)))) - {$signed($signed($signed(forvar2511))),
          (|forvar2510[(3'h7):(3'h5)])});
      for (forvar2522 = (1'h0); (forvar2522 < (1'h0)); forvar2522 = (forvar2522 + (1'h1)))
        begin
          if ($unsigned($unsigned(reg2503[(3'h5):(3'h5)])))
            begin
              reg2523 <= $unsigned(($unsigned($unsigned(reg2517)) ?
                  ($signed(wire2492) ?
                      (~&{(8'hb4)}) : ((8'hb8) == (~reg2504))) : ((~^(-(8'hae))) ^~ ($unsigned(reg2518) << reg2513[(3'h7):(3'h5)]))));
              reg2524 = wire2502[(3'h7):(1'h1)];
              reg2525 <= $unsigned((wire2502[(4'h8):(3'h4)] ?
                  (((reg2517 ? reg2524 : reg2499) ^ (^~reg2508)) > ({reg2518,
                      (7'h41)} && $unsigned(wire2505))) : reg2514[(5'h10):(3'h6)]));
            end
          else
            begin
              reg2523 = ((+(|forvar2511[(2'h2):(1'h0)])) >= (!((~&$signed(reg2508)) == reg2501)));
              reg2524 <= (|(($signed((reg2514 ^~ forvar2510)) ?
                  {(8'hbe)} : $unsigned({forvar2507, wire2492})) == (8'hb5)));
              reg2525 = forvar2510;
              reg2526 <= (8'hb0);
            end
          for (forvar2527 = (1'h0); (forvar2527 < (1'h0)); forvar2527 = (forvar2527 + (1'h1)))
            begin
              reg2528 = (reg2523[(4'h8):(4'h8)] ?
                  {forvar2511[(4'h9):(1'h0)],
                      reg2513} : {reg2497[(1'h1):(1'h1)],
                      (-((forvar2519 ? (8'hb9) : wire2493) ?
                          reg2512 : (reg2526 ? reg2512 : reg2523)))});
            end
          reg2529 <= reg2514[(3'h4):(2'h3)];
          for (forvar2530 = (1'h0); (forvar2530 < (2'h2)); forvar2530 = (forvar2530 + (1'h1)))
            begin
              reg2531 <= reg2512;
              reg2532 = $signed((reg2523 ^ ($unsigned($unsigned(wire2492)) && {wire2495,
                  (wire2502 * reg2525)})));
              reg2533 <= $signed(reg2513);
              reg2534 = {($unsigned(((reg2514 ?
                      reg2514 : (7'h42)) + reg2517[(3'h7):(3'h5)])) ~^ (reg2512[(4'hd):(3'h7)] >>> wire2495[(2'h3):(2'h3)]))};
              reg2535 = {(!reg2518)};
            end
          for (forvar2536 = (1'h0); (forvar2536 < (3'h4)); forvar2536 = (forvar2536 + (1'h1)))
            begin
              reg2537 <= {{(&reg2497[(1'h0):(1'h0)])}, (8'ha6)};
              reg2538 <= ($signed($signed((~|reg2532))) ?
                  (reg2528 ?
                      (~$unsigned((-reg2513))) : $unsigned($signed((reg2532 ?
                          reg2534 : reg2501)))) : (reg2520[(2'h2):(1'h0)] ?
                      $signed(($unsigned(reg2513) ?
                          (reg2517 || reg2528) : $signed(reg2508))) : wire2493));
              reg2539 = $unsigned(reg2533[(4'h8):(2'h2)]);
              reg2540 <= reg2513;
              reg2541 <= forvar2536[(2'h2):(1'h1)];
            end
        end
      reg2542 <= {$unsigned(reg2538)};
      if (reg2534)
        begin
          reg2543 <= $signed((reg2500 <= reg2513[(3'h5):(3'h5)]));
          reg2544 <= (~|{reg2538[(2'h3):(2'h2)]});
          reg2545 = $signed($unsigned($signed((reg2501 << {reg2533}))));
          reg2546 <= reg2518[(1'h0):(1'h0)];
        end
      else
        begin
          reg2543 <= {$signed($unsigned(reg2509[(1'h0):(1'h0)])),
              reg2521[(3'h7):(2'h3)]};
          reg2544 <= $signed((~&(($unsigned(reg2521) >> (^~reg2534)) || (wire2493[(4'he):(4'h8)] ?
              wire2505[(4'h9):(2'h2)] : $unsigned(reg2513)))));
          reg2545 = $signed(reg2529[(1'h0):(1'h0)]);
          reg2546 = $signed(reg2516);
          reg2547 <= (reg2512[(4'hd):(4'hd)] ^ $signed((~(wire2493[(1'h0):(1'h0)] > (~&(7'h40))))));
        end
      reg2548 <= (reg2514[(1'h1):(1'h1)] ?
          (!$unsigned(forvar2511[(3'h5):(3'h5)])) : ((&(7'h42)) ?
              reg2545 : $unsigned($signed(reg2525))));
    end
  always
    @(posedge clk) begin
      for (forvar2549 = (1'h0); (forvar2549 < (3'h4)); forvar2549 = (forvar2549 + (1'h1)))
        begin
          reg2550 <= (8'haa);
          reg2551 <= (($unsigned((wire2493[(4'he):(4'hc)] ?
                  (|reg2513) : {reg2501, forvar2527})) ?
              reg2500 : (reg2513[(3'h5):(2'h3)] ?
                  ($signed(reg2546) ?
                      (|(8'ha1)) : (reg2515 >> wire2502)) : reg2545[(3'h5):(3'h4)])) ^ reg2542);
          reg2552 <= reg2518;
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2402  (y, clk, wire2407, wire2406, wire2405, wire2404, wire2403);
  output wire [(32'h371):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire2407;
  input wire signed [(4'hc):(1'h0)] wire2406;
  input wire [(4'h8):(1'h0)] wire2405;
  input wire signed [(3'h6):(1'h0)] wire2404;
  input wire signed [(4'hc):(1'h0)] wire2403;
  reg signed [(5'h13):(1'h0)] reg2488 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2487 = (1'h0);
  reg [(5'h12):(1'h0)] reg2486 = (1'h0);
  reg [(2'h2):(1'h0)] reg2485 = (1'h0);
  reg [(4'h8):(1'h0)] reg2484 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2483 = (1'h0);
  reg [(3'h4):(1'h0)] reg2482 = (1'h0);
  reg [(4'ha):(1'h0)] reg2481 = (1'h0);
  reg [(4'hd):(1'h0)] reg2480 = (1'h0);
  reg [(4'hb):(1'h0)] reg2479 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2478 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2477 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2476 = (1'h0);
  reg [(4'hd):(1'h0)] reg2475 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2474 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2473 = (1'h0);
  reg [(4'ha):(1'h0)] reg2472 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2471 = (1'h0);
  reg [(4'ha):(1'h0)] reg2470 = (1'h0);
  reg [(5'h13):(1'h0)] reg2469 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2468 = (1'h0);
  reg [(3'h6):(1'h0)] reg2467 = (1'h0);
  reg [(4'hb):(1'h0)] reg2466 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2465 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2464 = (1'h0);
  reg [(4'hd):(1'h0)] reg2463 = (1'h0);
  reg [(5'h12):(1'h0)] reg2462 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2461 = (1'h0);
  reg [(5'h14):(1'h0)] reg2460 = (1'h0);
  reg [(4'h8):(1'h0)] reg2459 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2458 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2457 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2456 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire2455;
  reg signed [(2'h2):(1'h0)] reg2454 = (1'h0);
  reg [(3'h4):(1'h0)] reg2453 = (1'h0);
  reg [(3'h7):(1'h0)] reg2452 = (1'h0);
  reg [(4'he):(1'h0)] reg2451 = (1'h0);
  reg [(4'h9):(1'h0)] reg2450 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2449 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire2448;
  reg signed [(3'h5):(1'h0)] reg2447 = (1'h0);
  reg [(3'h4):(1'h0)] reg2446 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2445 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2444 = (1'h0);
  reg [(4'hb):(1'h0)] reg2443 = (1'h0);
  reg [(4'ha):(1'h0)] reg2442 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2441 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2440 = (1'h0);
  reg [(2'h3):(1'h0)] reg2439 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2438 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2437 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2436 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2435 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2434 = (1'h0);
  wire [(2'h3):(1'h0)] wire2433;
  reg [(5'h12):(1'h0)] reg2432 = (1'h0);
  reg [(2'h2):(1'h0)] reg2431 = (1'h0);
  reg [(2'h2):(1'h0)] reg2430 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2429 = (1'h0);
  reg [(5'h13):(1'h0)] reg2428 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire2427;
  reg signed [(4'hf):(1'h0)] reg2426 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2425 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2424 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2423 = (1'h0);
  reg [(4'hb):(1'h0)] reg2422 = (1'h0);
  reg [(4'hb):(1'h0)] reg2421 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2420 = (1'h0);
  reg [(3'h4):(1'h0)] reg2419 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2418 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2417 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2416 = (1'h0);
  reg [(4'hd):(1'h0)] reg2415 = (1'h0);
  reg [(5'h10):(1'h0)] reg2414 = (1'h0);
  reg [(5'h13):(1'h0)] reg2413 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2412 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2411 = (1'h0);
  reg [(3'h6):(1'h0)] reg2410 = (1'h0);
  wire [(3'h4):(1'h0)] wire2409;
  wire signed [(5'h12):(1'h0)] wire2408;
  assign y = {reg2488,
                 reg2487,
                 reg2486,
                 reg2485,
                 reg2484,
                 reg2483,
                 reg2482,
                 reg2481,
                 reg2480,
                 reg2479,
                 forvar2478,
                 reg2477,
                 reg2476,
                 reg2475,
                 reg2474,
                 reg2473,
                 reg2472,
                 forvar2471,
                 reg2470,
                 reg2469,
                 reg2468,
                 reg2467,
                 reg2466,
                 forvar2465,
                 forvar2464,
                 reg2463,
                 reg2462,
                 reg2461,
                 reg2460,
                 reg2459,
                 reg2458,
                 reg2457,
                 reg2456,
                 wire2455,
                 reg2454,
                 reg2453,
                 reg2452,
                 reg2451,
                 reg2450,
                 forvar2449,
                 wire2448,
                 reg2447,
                 reg2446,
                 reg2445,
                 reg2444,
                 reg2443,
                 reg2442,
                 reg2441,
                 reg2440,
                 reg2439,
                 forvar2438,
                 reg2437,
                 reg2436,
                 forvar2435,
                 reg2434,
                 wire2433,
                 reg2432,
                 reg2431,
                 reg2430,
                 reg2429,
                 reg2428,
                 wire2427,
                 reg2426,
                 reg2425,
                 reg2424,
                 reg2423,
                 reg2422,
                 reg2421,
                 forvar2420,
                 reg2419,
                 forvar2418,
                 forvar2417,
                 reg2416,
                 reg2415,
                 reg2414,
                 reg2413,
                 forvar2412,
                 reg2411,
                 reg2410,
                 wire2409,
                 wire2408,
                 (1'h0)};
  assign wire2408 = wire2404;
  assign wire2409 = $unsigned(wire2404[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      reg2410 <= ((8'hb8) ^~ wire2406[(3'h6):(2'h3)]);
      reg2411 <= $unsigned(wire2404);
      for (forvar2412 = (1'h0); (forvar2412 < (3'h4)); forvar2412 = (forvar2412 + (1'h1)))
        begin
          reg2413 <= wire2406;
        end
      reg2414 <= wire2407[(4'h8):(4'h8)];
      reg2415 <= ($signed(((~&(wire2409 > reg2411)) ?
          (+$unsigned(forvar2412)) : ({forvar2412} ?
              $signed(wire2406) : (~^(8'haa))))) >> $signed((|({wire2407,
              reg2411} ?
          (wire2409 & wire2407) : $unsigned((8'hb2))))));
    end
  always
    @(posedge clk) begin
      reg2416 = (reg2411 + $signed((&reg2414)));
      for (forvar2417 = (1'h0); (forvar2417 < (1'h1)); forvar2417 = (forvar2417 + (1'h1)))
        begin
          for (forvar2418 = (1'h0); (forvar2418 < (1'h1)); forvar2418 = (forvar2418 + (1'h1)))
            begin
              reg2419 = $unsigned((reg2411[(1'h0):(1'h0)] >= wire2403));
            end
          for (forvar2420 = (1'h0); (forvar2420 < (3'h4)); forvar2420 = (forvar2420 + (1'h1)))
            begin
              reg2421 <= ((!wire2408) + (((8'ha9) ?
                      ({wire2405} <= (-wire2406)) : wire2404) ?
                  (wire2408 ^~ {{reg2419, reg2414},
                      $signed((8'ha2))}) : wire2408));
              reg2422 <= reg2410[(2'h3):(2'h2)];
              reg2423 = reg2415;
              reg2424 <= (|$signed(wire2409));
            end
        end
      reg2425 <= $signed($unsigned($unsigned((reg2411 || $unsigned(forvar2418)))));
      reg2426 <= ($unsigned(({$unsigned((8'hbe))} ?
          ((|reg2413) ?
              (^wire2403) : {wire2405}) : reg2422[(3'h6):(2'h3)])) ^ $signed((~&(&reg2411[(4'hc):(4'ha)]))));
    end
  assign wire2427 = reg2411;
  always
    @(posedge clk) begin
      reg2428 <= (($unsigned($unsigned($unsigned(reg2414))) ?
              reg2425[(2'h3):(2'h3)] : (8'hbd)) ?
          $unsigned($unsigned((^~wire2403[(3'h7):(1'h1)]))) : wire2406);
      reg2429 <= reg2423;
      reg2430 <= $unsigned(reg2428[(5'h12):(4'he)]);
      reg2431 <= (($unsigned($unsigned(((8'ha2) ?
              forvar2418 : wire2404))) < $signed((~(reg2421 ?
              forvar2418 : reg2416)))) ?
          (reg2428 ?
              forvar2420[(3'h4):(2'h3)] : (^((wire2407 ? reg2429 : (8'ha3)) ?
                  (~reg2423) : (reg2425 | wire2427)))) : $signed((({(8'hab)} ^ reg2421[(1'h0):(1'h0)]) ?
              {$signed(forvar2420)} : $signed({forvar2412}))));
    end
  always
    @(posedge clk) begin
      reg2432 <= $unsigned(reg2429[(4'hd):(1'h0)]);
    end
  assign wire2433 = reg2422;
  always
    @(posedge clk) begin
      reg2434 <= $signed($unsigned({$signed(wire2433),
          (~^(reg2414 >= reg2415))}));
      for (forvar2435 = (1'h0); (forvar2435 < (2'h2)); forvar2435 = (forvar2435 + (1'h1)))
        begin
          reg2436 = (reg2416[(4'h9):(3'h6)] ?
              $unsigned($unsigned($unsigned((reg2414 ?
                  forvar2435 : reg2419)))) : $unsigned(($signed((forvar2420 ?
                      (8'ha3) : wire2407)) ?
                  forvar2435 : ($unsigned(reg2419) ?
                      $signed(wire2403) : {wire2406}))));
          reg2437 = $signed({$unsigned({$signed(wire2406),
                  {forvar2417, wire2409}}),
              (reg2410 ?
                  {$unsigned(wire2433), wire2427} : $signed({forvar2412,
                      wire2403}))});
          for (forvar2438 = (1'h0); (forvar2438 < (2'h3)); forvar2438 = (forvar2438 + (1'h1)))
            begin
              reg2439 <= (forvar2438 ?
                  (reg2410[(1'h0):(1'h0)] ?
                      forvar2420 : reg2414) : $unsigned(((wire2404[(1'h1):(1'h1)] || (~(8'hba))) ?
                      ({(8'hbe)} ?
                          (&reg2428) : $unsigned(reg2422)) : reg2411)));
              reg2440 <= $signed(({wire2433[(1'h0):(1'h0)]} == reg2426));
              reg2441 <= $signed(forvar2412[(4'h9):(3'h4)]);
              reg2442 <= $unsigned((($unsigned(reg2425[(1'h0):(1'h0)]) || {{reg2413,
                      reg2429}}) == (!{forvar2420,
                  forvar2438[(4'he):(3'h5)]})));
            end
        end
      reg2443 <= (|$signed(($signed($unsigned(reg2416)) ?
          reg2415[(3'h5):(2'h3)] : $unsigned($signed(wire2433)))));
      reg2444 <= reg2423;
      reg2445 = wire2407;
    end
  always
    @(posedge clk) begin
      reg2446 <= (8'hb3);
      reg2447 <= reg2415;
    end
  assign wire2448 = $unsigned(wire2405[(3'h5):(2'h3)]);
  always
    @(posedge clk) begin
      for (forvar2449 = (1'h0); (forvar2449 < (2'h2)); forvar2449 = (forvar2449 + (1'h1)))
        begin
          reg2450 <= wire2404;
          reg2451 <= wire2405[(3'h6):(2'h2)];
        end
      reg2452 <= $unsigned((-$unsigned((reg2428[(2'h2):(2'h2)] ?
          forvar2438 : $signed(forvar2438)))));
      reg2453 <= {{($unsigned((8'ha4)) ? $signed((|(8'hbe))) : reg2443),
              (forvar2438 ? (~&$unsigned(reg2441)) : reg2429)},
          ($unsigned(reg2413) ?
              (((reg2434 << reg2425) ?
                      (wire2408 ? reg2439 : (7'h42)) : $unsigned(reg2429)) ?
                  (!{reg2424}) : ((wire2448 == forvar2449) >>> wire2403[(4'h8):(2'h2)])) : ($signed((reg2424 ?
                      reg2442 : forvar2417)) ?
                  $signed($unsigned((8'h9e))) : reg2451))};
      reg2454 <= wire2427[(1'h0):(1'h0)];
    end
  assign wire2455 = {wire2408[(4'h8):(1'h0)], $signed(wire2408[(2'h3):(1'h0)])};
  always
    @(posedge clk) begin
      reg2456 <= reg2447[(3'h4):(1'h1)];
      reg2457 <= ($unsigned($signed((8'ha6))) > wire2405[(1'h0):(1'h0)]);
      reg2458 <= forvar2420[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg2459 <= forvar2420;
      reg2460 <= {$unsigned($unsigned((!reg2411))),
          ($signed(forvar2438[(4'hb):(1'h1)]) >= (8'hba))};
      reg2461 <= wire2408;
      reg2462 = (~^$signed(reg2419[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg2463 <= ($signed((&(((8'hb9) + reg2416) ?
              ((8'ha4) ? (8'hbb) : reg2434) : reg2414[(4'hd):(4'hc)]))) ?
          wire2404 : (~^(((reg2431 ? (8'hb0) : reg2430) < (forvar2412 ?
              forvar2435 : forvar2449)) < ((forvar2449 >>> reg2443) ^ $signed(reg2461)))));
    end
  always
    @(posedge clk) begin
      for (forvar2464 = (1'h0); (forvar2464 < (2'h2)); forvar2464 = (forvar2464 + (1'h1)))
        begin
          for (forvar2465 = (1'h0); (forvar2465 < (2'h2)); forvar2465 = (forvar2465 + (1'h1)))
            begin
              reg2466 <= reg2463[(4'h9):(2'h3)];
              reg2467 <= reg2443;
              reg2468 <= {($unsigned(reg2432) < {((~reg2439) ?
                          {reg2456} : $unsigned(reg2434)),
                      $unsigned(((8'h9f) ? reg2459 : reg2461))}),
                  ((($signed(wire2403) ?
                              (reg2410 * reg2430) : (reg2429 ?
                                  reg2416 : wire2405)) ?
                          (&(wire2406 ?
                              (8'h9c) : reg2421)) : reg2430[(2'h2):(1'h0)]) ?
                      (~|(reg2439[(2'h3):(1'h0)] && reg2458[(4'hb):(2'h2)])) : reg2460)};
            end
        end
    end
  always
    @(posedge clk) begin
      reg2469 <= (reg2457 & $unsigned(((8'hbb) && reg2429[(4'ha):(4'h9)])));
    end
  always
    @(posedge clk) begin
      reg2470 <= $unsigned(reg2430[(1'h0):(1'h0)]);
      for (forvar2471 = (1'h0); (forvar2471 < (2'h3)); forvar2471 = (forvar2471 + (1'h1)))
        begin
          reg2472 = reg2422[(4'h9):(4'h9)];
          reg2473 <= {reg2467};
        end
      reg2474 <= (reg2443[(2'h3):(1'h1)] | (wire2408 ?
          $signed((~&reg2454[(2'h2):(1'h1)])) : $unsigned($signed(((8'hb6) ^ (8'hb7))))));
      reg2475 <= ((reg2439 ~^ (^reg2416[(4'ha):(3'h7)])) ?
          {reg2444} : {(~|$signed({(8'hbe), reg2436}))});
    end
  always
    @(posedge clk) begin
      reg2476 <= reg2457[(1'h1):(1'h1)];
      reg2477 <= {{$unsigned(reg2439), (^~wire2405)}};
      for (forvar2478 = (1'h0); (forvar2478 < (2'h2)); forvar2478 = (forvar2478 + (1'h1)))
        begin
          reg2479 = $signed(({$unsigned(forvar2417)} > reg2450));
          reg2480 <= (((((reg2454 >> reg2431) ?
              (wire2406 ?
                  (8'had) : reg2446) : ((8'hbf) ~^ reg2413)) << reg2468[(3'h5):(2'h3)]) >> (|wire2455[(3'h4):(2'h2)])) || (((|$unsigned(forvar2420)) ~^ reg2424[(3'h7):(3'h6)]) ?
              (!(^$signed(reg2413))) : (~|reg2446)));
          reg2481 = {reg2411};
        end
      reg2482 <= reg2481[(3'h6):(2'h2)];
      reg2483 <= (((^{forvar2418, {forvar2420, forvar2465}}) ?
              (reg2457 ?
                  ((reg2462 == reg2426) >>> (8'ha4)) : $unsigned($signed(reg2453))) : $unsigned((8'ha3))) ?
          reg2458 : ({($signed((8'ha4)) <<< $signed(reg2446))} >> reg2470[(3'h5):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg2484 = ((~wire2427[(1'h0):(1'h0)]) ?
          $signed(wire2405[(3'h7):(3'h5)]) : ((reg2470[(1'h0):(1'h0)] ^~ $signed($signed((8'hb9)))) ?
              (7'h40) : reg2466[(4'hb):(4'h8)]));
      reg2485 <= ((|$signed((~&reg2424[(3'h6):(3'h6)]))) ?
          ({$signed({forvar2449, (8'ha1)}), (8'h9d)} ?
              (($unsigned(reg2468) ^ $unsigned(wire2408)) ^ wire2433[(2'h2):(1'h0)]) : $signed(reg2428[(4'hd):(1'h0)])) : $unsigned(reg2462[(4'hf):(1'h1)]));
    end
  always
    @(posedge clk) begin
      reg2486 <= $unsigned(($signed($unsigned($signed((8'hb7)))) ?
          {forvar2471, $unsigned(forvar2449)} : (~|$signed((8'haf)))));
      reg2487 = {wire2448,
          $signed({reg2468, ($unsigned(wire2427) ? (-reg2429) : (8'had))})};
      reg2488 <= $signed(reg2486);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2375  (y, clk, wire2380, wire2379, wire2378, wire2377, wire2376);
  output wire [(32'h8b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire2380;
  input wire signed [(4'he):(1'h0)] wire2379;
  input wire [(5'h10):(1'h0)] wire2378;
  input wire signed [(5'h13):(1'h0)] wire2377;
  input wire [(3'h5):(1'h0)] wire2376;
  wire [(4'hc):(1'h0)] wire2392;
  wire [(5'h13):(1'h0)] wire2391;
  wire [(4'hb):(1'h0)] wire2390;
  wire signed [(4'hf):(1'h0)] wire2389;
  wire [(4'h9):(1'h0)] wire2388;
  reg [(4'hd):(1'h0)] reg2387 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire2386;
  reg [(2'h2):(1'h0)] reg2385 = (1'h0);
  reg [(5'h11):(1'h0)] reg2384 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2383 = (1'h0);
  reg [(2'h3):(1'h0)] reg2382 = (1'h0);
  wire [(5'h11):(1'h0)] wire2381;
  assign y = {wire2392,
                 wire2391,
                 wire2390,
                 wire2389,
                 wire2388,
                 reg2387,
                 wire2386,
                 reg2385,
                 reg2384,
                 reg2383,
                 reg2382,
                 wire2381,
                 (1'h0)};
  assign wire2381 = $signed($signed({$signed({wire2377}),
                        wire2380[(1'h0):(1'h0)]}));
  always
    @(posedge clk) begin
      reg2382 <= (-((^(((8'hb3) ? (8'had) : (8'hb6)) ?
              $unsigned(wire2379) : wire2378)) ?
          wire2381[(3'h7):(3'h4)] : wire2380[(1'h0):(1'h0)]));
      reg2383 = (!wire2381[(3'h7):(2'h3)]);
      reg2384 <= reg2382;
      reg2385 <= {(reg2383[(2'h2):(2'h2)] << $signed(reg2384)),
          ($unsigned((^~$signed(reg2382))) ?
              reg2382 : (~&{$unsigned(reg2384),
                  (wire2376 ? reg2383 : reg2384)}))};
    end
  assign wire2386 = reg2383;
  always
    @(posedge clk) begin
      reg2387 <= ($signed((~^((&wire2386) ?
          (wire2376 <<< wire2379) : wire2380))) - ($unsigned(wire2377[(3'h6):(3'h6)]) <= {reg2385,
          (wire2377[(4'h9):(4'h9)] ?
              ((8'hb7) < wire2381) : $unsigned(wire2379))}));
    end
  assign wire2388 = $signed((-$unsigned(wire2376)));
  assign wire2389 = (~reg2383);
  assign wire2390 = $unsigned(reg2382[(1'h1):(1'h0)]);
  assign wire2391 = {{wire2386[(3'h4):(3'h4)]}};
  assign wire2392 = ($signed(((wire2386 ?
                                $unsigned(reg2382) : $unsigned(wire2389)) ?
                            wire2389[(3'h7):(1'h0)] : {reg2382[(2'h3):(2'h3)],
                                (wire2381 ? reg2384 : wire2391)})) ?
                        (^$signed($signed(wire2391))) : wire2389);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2314
#( parameter param2363 = (~^(((((8'hbe) ? (8'haa) : (8'haf)) ? ((8'ha2) ? (8'hae) : (8'hbe)) : ((7'h42) ? (8'hb9) : (7'h42))) ^~ (((8'ha1) ? (8'hbc) : (8'hb6)) - ((8'ha9) << (8'hac)))) ^~ (^{(~|(8'hab)), ((8'ha0) >> (8'hae))}))) )
(y, clk, wire2319, wire2318, wire2317, wire2316, wire2315);
  output wire [(32'h1c3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire2319;
  input wire signed [(4'hc):(1'h0)] wire2318;
  input wire signed [(3'h5):(1'h0)] wire2317;
  input wire [(4'hb):(1'h0)] wire2316;
  input wire signed [(3'h5):(1'h0)] wire2315;
  reg [(4'hf):(1'h0)] reg2362 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2361 = (1'h0);
  reg [(2'h3):(1'h0)] reg2360 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2359 = (1'h0);
  reg [(4'he):(1'h0)] reg2358 = (1'h0);
  reg [(4'hf):(1'h0)] reg2357 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2356 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2355 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2354 = (1'h0);
  reg [(3'h7):(1'h0)] reg2353 = (1'h0);
  reg [(4'ha):(1'h0)] reg2352 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2351 = (1'h0);
  reg [(4'h8):(1'h0)] reg2350 = (1'h0);
  wire [(5'h12):(1'h0)] wire2349;
  reg signed [(5'h11):(1'h0)] reg2348 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2347 = (1'h0);
  reg [(3'h6):(1'h0)] reg2346 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2345 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2344 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2343 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2342 = (1'h0);
  reg [(4'hb):(1'h0)] reg2341 = (1'h0);
  wire [(4'he):(1'h0)] wire2340;
  wire signed [(4'h8):(1'h0)] wire2339;
  reg signed [(2'h3):(1'h0)] reg2338 = (1'h0);
  reg [(4'h9):(1'h0)] reg2337 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2336 = (1'h0);
  reg [(4'hf):(1'h0)] reg2335 = (1'h0);
  wire signed [(4'he):(1'h0)] wire2334;
  reg signed [(5'h13):(1'h0)] reg2333 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2332 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2331 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2330 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2329 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2328 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2327 = (1'h0);
  reg [(3'h6):(1'h0)] reg2326 = (1'h0);
  reg [(4'h8):(1'h0)] reg2325 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2324 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2323 = (1'h0);
  reg [(3'h7):(1'h0)] reg2322 = (1'h0);
  reg [(4'h9):(1'h0)] reg2321 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2320 = (1'h0);
  assign y = {reg2362,
                 reg2361,
                 reg2360,
                 reg2359,
                 reg2358,
                 reg2357,
                 reg2356,
                 reg2355,
                 reg2354,
                 reg2353,
                 reg2352,
                 reg2351,
                 reg2350,
                 wire2349,
                 reg2348,
                 reg2347,
                 reg2346,
                 forvar2345,
                 reg2344,
                 reg2343,
                 reg2342,
                 reg2341,
                 wire2340,
                 wire2339,
                 reg2338,
                 reg2337,
                 reg2336,
                 reg2335,
                 wire2334,
                 reg2333,
                 reg2332,
                 reg2331,
                 reg2330,
                 reg2329,
                 reg2328,
                 reg2327,
                 reg2326,
                 reg2325,
                 reg2324,
                 reg2323,
                 reg2322,
                 reg2321,
                 forvar2320,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar2320 = (1'h0); (forvar2320 < (2'h3)); forvar2320 = (forvar2320 + (1'h1)))
        begin
          if ((wire2318 * (+$signed({$signed((8'ha7)), $signed(forvar2320)}))))
            begin
              reg2321 = wire2318[(2'h3):(1'h0)];
            end
          else
            begin
              reg2321 <= (&$signed($unsigned(($signed(reg2321) ?
                  wire2317[(3'h4):(2'h2)] : wire2319[(3'h7):(2'h2)]))));
              reg2322 <= ((((wire2315 ?
                          forvar2320[(3'h6):(1'h0)] : (|reg2321)) ?
                      forvar2320 : forvar2320[(3'h7):(1'h1)]) << (&wire2318[(3'h4):(1'h0)])) ?
                  wire2318 : (-wire2316));
              reg2323 <= {{reg2321,
                      ($unsigned((wire2316 - forvar2320)) <<< wire2319)}};
              reg2324 <= $unsigned($unsigned({(8'hbd)}));
              reg2325 <= $signed($signed((7'h41)));
            end
          reg2326 <= (wire2317[(2'h2):(1'h0)] ?
              wire2319[(2'h3):(2'h3)] : reg2324[(3'h6):(2'h3)]);
          reg2327 <= $signed(({(&$signed((8'hab))),
              forvar2320[(1'h1):(1'h0)]} <<< ({$signed(wire2319),
              (~^(7'h43))} - ($unsigned(wire2315) ?
              ((8'ha6) ^ reg2325) : ((8'ha8) ? (8'ha9) : reg2326)))));
          reg2328 <= wire2319;
        end
      reg2329 <= (~^wire2319);
      reg2330 <= (8'hb5);
    end
  always
    @(posedge clk) begin
      reg2331 <= reg2323[(4'h9):(3'h6)];
      reg2332 = $signed($unsigned({(^(reg2331 ? reg2328 : (8'hbc)))}));
      reg2333 <= ($signed((reg2330[(4'he):(3'h4)] + wire2317)) >= {(~|reg2332[(4'ha):(1'h0)])});
    end
  assign wire2334 = $unsigned(reg2329);
  always
    @(posedge clk) begin
      reg2335 = $signed($unsigned({$unsigned((~|wire2317)), (^~reg2332)}));
    end
  always
    @(posedge clk) begin
      reg2336 <= ((($unsigned((wire2317 & reg2330)) ?
              reg2331[(2'h2):(1'h0)] : (-reg2330[(4'he):(1'h0)])) == reg2322) ?
          reg2323[(4'ha):(2'h3)] : (~^wire2318[(3'h7):(2'h3)]));
      reg2337 = {reg2326[(3'h4):(2'h3)], $unsigned(reg2332)};
      reg2338 <= (({reg2333[(5'h10):(3'h7)], forvar2320} ?
              (({reg2333, reg2337} ? $signed(reg2329) : $signed(reg2324)) ?
                  ((reg2337 * reg2335) ?
                      (^~wire2317) : $signed(reg2330)) : $unsigned(wire2316[(3'h4):(2'h2)])) : wire2317[(3'h5):(2'h2)]) ?
          {wire2317, $unsigned(wire2316)} : (~&wire2317));
    end
  assign wire2339 = reg2323[(1'h1):(1'h0)];
  assign wire2340 = (!(forvar2320 ?
                        (!$signed((reg2337 ?
                            (8'hbd) : reg2330))) : (reg2337 < $signed({reg2333,
                            reg2335}))));
  always
    @(posedge clk) begin
      reg2341 <= wire2316[(1'h0):(1'h0)];
      reg2342 = $unsigned((reg2328 ?
          ($signed((reg2338 >= reg2336)) && wire2315[(1'h0):(1'h0)]) : reg2324));
      reg2343 = $signed($signed(reg2333));
      reg2344 = {(^~reg2342[(2'h2):(1'h1)]),
          $unsigned(($signed($signed(wire2316)) ^~ $signed((!wire2339))))};
    end
  always
    @(posedge clk) begin
      for (forvar2345 = (1'h0); (forvar2345 < (1'h1)); forvar2345 = (forvar2345 + (1'h1)))
        begin
          reg2346 <= $unsigned($signed($signed($signed((~&wire2340)))));
        end
      reg2347 <= ((-((&wire2340) ?
          wire2317 : (8'haf))) ^~ $signed(((~&$signed(wire2319)) ?
          (8'ha4) : reg2338[(2'h3):(2'h3)])));
      reg2348 <= {wire2317[(1'h1):(1'h1)],
          (reg2342[(3'h4):(1'h0)] + (((wire2340 ? wire2340 : reg2337) ?
                  $signed((8'ha3)) : reg2344[(3'h6):(3'h4)]) ?
              reg2331 : (reg2344 <= $unsigned(reg2322))))};
    end
  assign wire2349 = $unsigned({($unsigned(reg2341[(3'h4):(1'h0)]) << reg2325),
                        (reg2322[(1'h1):(1'h0)] != wire2318)});
  always
    @(posedge clk) begin
      reg2350 <= ((8'hb7) <= $signed($signed(($signed(wire2349) ?
          (reg2327 ? reg2342 : reg2321) : reg2321[(3'h5):(1'h1)]))));
      reg2351 = (wire2315[(1'h1):(1'h1)] ?
          $signed(wire2334[(3'h7):(1'h1)]) : reg2344);
      reg2352 = $signed((((8'h9e) ?
          wire2315 : $signed(wire2316)) && ((~$unsigned(reg2333)) | (~^(wire2315 << forvar2345)))));
    end
  always
    @(posedge clk) begin
      reg2353 = $unsigned(((!reg2344) ?
          (reg2343[(3'h4):(1'h0)] != ($signed(reg2347) ?
              wire2339 : reg2350[(3'h7):(1'h0)])) : (reg2351 > (^~{wire2339,
              (8'hae)}))));
      if (($signed((+({wire2317, reg2342} ?
          (~^(7'h43)) : reg2329))) | (|$unsigned(wire2339[(3'h7):(3'h6)]))))
        begin
          reg2354 <= reg2353;
          reg2355 <= ($signed((!reg2350)) != $unsigned((~|$signed($signed(reg2352)))));
          reg2356 <= (8'h9c);
        end
      else
        begin
          reg2354 <= {reg2332};
          reg2355 <= $signed((~|$unsigned(reg2330)));
          reg2356 <= (^(-(&((~&(8'hb1)) ^~ wire2316))));
        end
      reg2357 <= ($unsigned((^{reg2347})) ?
          ((reg2321 >= reg2347[(3'h4):(1'h1)]) && $unsigned((&(reg2347 >> reg2342)))) : $unsigned($signed((+reg2325[(3'h4):(1'h1)]))));
    end
  always
    @(posedge clk) begin
      reg2358 <= (|$unsigned((reg2338[(2'h3):(2'h3)] ^~ (^{wire2316}))));
      reg2359 <= $unsigned((^$signed((reg2327[(1'h0):(1'h0)] ?
          reg2354[(5'h10):(1'h0)] : (8'hb6)))));
      reg2360 <= {$unsigned(reg2337[(1'h1):(1'h1)])};
      reg2361 = (-(~|$unsigned((+wire2349))));
      reg2362 <= ({forvar2320[(1'h1):(1'h1)]} >= $signed($signed(($signed(reg2354) + (wire2317 ?
          reg2351 : forvar2345)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2254  (y, clk, wire2259, wire2258, wire2257, wire2256, wire2255);
  output wire [(32'h26e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire2259;
  input wire signed [(4'ha):(1'h0)] wire2258;
  input wire [(2'h3):(1'h0)] wire2257;
  input wire signed [(5'h13):(1'h0)] wire2256;
  input wire [(2'h3):(1'h0)] wire2255;
  reg signed [(5'h15):(1'h0)] reg2306 = (1'h0);
  reg [(4'ha):(1'h0)] reg2305 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2304 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire2303;
  wire [(4'h9):(1'h0)] wire2302;
  reg [(5'h12):(1'h0)] reg2301 = (1'h0);
  wire [(5'h12):(1'h0)] wire2300;
  reg signed [(5'h13):(1'h0)] reg2299 = (1'h0);
  reg [(4'h8):(1'h0)] reg2298 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2297 = (1'h0);
  reg [(5'h12):(1'h0)] reg2296 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2295 = (1'h0);
  reg [(3'h7):(1'h0)] reg2294 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2293 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2292 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire2291;
  wire [(5'h15):(1'h0)] wire2290;
  reg [(3'h7):(1'h0)] reg2289 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2288 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2287 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2286 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2285 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2284 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2283 = (1'h0);
  reg [(4'hb):(1'h0)] reg2282 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2281 = (1'h0);
  reg [(5'h11):(1'h0)] reg2280 = (1'h0);
  wire [(3'h6):(1'h0)] wire2279;
  reg [(5'h12):(1'h0)] reg2278 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2277 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2276 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2275 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2274 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2273 = (1'h0);
  reg [(4'hd):(1'h0)] reg2272 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2271 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2270 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2269 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2268 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2267 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2266 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2265 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2264 = (1'h0);
  reg [(2'h2):(1'h0)] reg2263 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2262 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire2261;
  reg signed [(5'h13):(1'h0)] reg2260 = (1'h0);
  assign y = {reg2306,
                 reg2305,
                 reg2304,
                 wire2303,
                 wire2302,
                 reg2301,
                 wire2300,
                 reg2299,
                 reg2298,
                 reg2297,
                 reg2296,
                 reg2295,
                 reg2294,
                 forvar2293,
                 reg2292,
                 wire2291,
                 wire2290,
                 reg2289,
                 reg2288,
                 reg2287,
                 reg2286,
                 reg2285,
                 reg2284,
                 reg2283,
                 reg2282,
                 forvar2281,
                 reg2280,
                 wire2279,
                 reg2278,
                 reg2277,
                 reg2276,
                 forvar2275,
                 forvar2274,
                 reg2273,
                 reg2272,
                 reg2271,
                 reg2270,
                 reg2269,
                 forvar2268,
                 reg2267,
                 reg2266,
                 reg2265,
                 reg2264,
                 reg2263,
                 reg2262,
                 wire2261,
                 reg2260,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg2260 <= wire2258[(2'h2):(1'h1)];
    end
  assign wire2261 = $unsigned(((($signed((8'h9d)) >> (~wire2256)) ?
                        (~&(wire2256 < wire2257)) : ($signed(wire2256) << $unsigned(wire2259))) << reg2260));
  always
    @(posedge clk) begin
      reg2262 <= wire2258;
      reg2263 <= (reg2260 && reg2260[(4'he):(4'h8)]);
      reg2264 <= $unsigned((~|{(~|{wire2256}), reg2262}));
    end
  always
    @(posedge clk) begin
      reg2265 <= reg2264[(4'h8):(4'h8)];
      reg2266 <= (($unsigned({(~&wire2256),
          (wire2256 ?
              reg2262 : (8'hb8))}) | (8'h9e)) << $unsigned($signed($unsigned((~wire2257)))));
      reg2267 <= wire2255[(1'h0):(1'h0)];
      for (forvar2268 = (1'h0); (forvar2268 < (3'h4)); forvar2268 = (forvar2268 + (1'h1)))
        begin
          reg2269 = ($unsigned((((8'haf) ?
              wire2259[(2'h2):(1'h0)] : (^wire2257)) ~^ (^(wire2257 >> reg2263)))) | forvar2268[(3'h4):(3'h4)]);
          reg2270 <= $signed((-reg2266));
          reg2271 = {reg2269};
          reg2272 <= (^~$signed(reg2267));
          reg2273 <= ((($signed(wire2256) ?
                  wire2256 : ($unsigned((8'hb6)) && $unsigned(reg2269))) && ((reg2269[(3'h4):(3'h4)] ?
                      reg2264 : (wire2256 != (8'haf))) ?
                  reg2270 : (reg2269[(3'h7):(1'h0)] | reg2264[(3'h6):(3'h4)]))) ?
              (wire2261[(1'h0):(1'h0)] ?
                  $signed((((8'hb1) | reg2263) > (forvar2268 ?
                      reg2272 : wire2255))) : ((^$unsigned((8'ha0))) ^ $signed({wire2258}))) : ($signed(((reg2270 && reg2267) | reg2270)) - $unsigned(reg2263)));
        end
      for (forvar2274 = (1'h0); (forvar2274 < (2'h2)); forvar2274 = (forvar2274 + (1'h1)))
        begin
          for (forvar2275 = (1'h0); (forvar2275 < (1'h0)); forvar2275 = (forvar2275 + (1'h1)))
            begin
              reg2276 <= ($unsigned(reg2272) ?
                  (((^~wire2257) || $unsigned((reg2264 ?
                      reg2265 : wire2255))) <= wire2261) : $unsigned((&($signed((8'ha6)) ?
                      (~(8'hb9)) : (reg2265 ? wire2257 : reg2265)))));
              reg2277 <= $unsigned(reg2270[(3'h6):(3'h4)]);
            end
          reg2278 = wire2259[(1'h1):(1'h0)];
        end
    end
  assign wire2279 = {reg2260[(4'hd):(4'hc)]};
  always
    @(posedge clk) begin
      reg2280 <= wire2257[(2'h3):(1'h0)];
      for (forvar2281 = (1'h0); (forvar2281 < (2'h2)); forvar2281 = (forvar2281 + (1'h1)))
        begin
          reg2282 <= ($signed(reg2270[(4'h8):(3'h4)]) ?
              $signed((reg2272 <= (~&(forvar2274 + reg2267)))) : (+forvar2281[(3'h4):(1'h0)]));
          reg2283 <= reg2260;
          reg2284 <= reg2262[(5'h11):(5'h10)];
          reg2285 <= $unsigned(reg2262[(4'h9):(3'h7)]);
          reg2286 = (7'h42);
        end
      reg2287 <= ($unsigned((~^reg2282)) || (reg2283 <= ((+(wire2258 ?
          forvar2268 : reg2286)) || wire2261[(1'h1):(1'h0)])));
      reg2288 <= (!reg2262[(3'h5):(3'h5)]);
      reg2289 = (((~forvar2274[(1'h0):(1'h0)]) < (~&reg2287)) ?
          (8'ha5) : ($signed((~&(~^reg2273))) ?
              $signed(forvar2268) : {(-{reg2282}), reg2285[(4'hb):(3'h7)]}));
    end
  assign wire2290 = (^~{((reg2280 <<< $unsigned(wire2256)) ?
                            $unsigned(forvar2274) : $unsigned((reg2260 ?
                                wire2257 : reg2289))),
                        $signed(reg2286[(3'h4):(2'h2)])});
  assign wire2291 = $unsigned($unsigned($signed(reg2277[(5'h12):(4'h9)])));
  always
    @(posedge clk) begin
      reg2292 <= reg2266[(1'h0):(1'h0)];
      for (forvar2293 = (1'h0); (forvar2293 < (2'h2)); forvar2293 = (forvar2293 + (1'h1)))
        begin
          reg2294 <= reg2289[(3'h7):(3'h6)];
          reg2295 <= ((reg2278 ?
              reg2280 : ((~forvar2275[(2'h2):(2'h2)]) ?
                  $unsigned(forvar2281[(5'h14):(5'h13)]) : ({reg2292,
                      reg2263} ^ $unsigned(wire2279)))) < $signed($signed(reg2289)));
          reg2296 <= (^($unsigned((8'hb5)) ?
              reg2265[(3'h4):(2'h3)] : wire2257[(1'h0):(1'h0)]));
        end
      reg2297 <= {{($signed($unsigned(reg2284)) ?
                  $signed((reg2260 ? reg2263 : wire2291)) : (forvar2275 ?
                      $unsigned(reg2273) : reg2287)),
              $signed((((8'ha9) ? wire2259 : wire2290) > {reg2269}))}};
      reg2298 <= $signed(($signed(wire2258) == (~^($unsigned(wire2279) - $unsigned((8'ha0))))));
      reg2299 = $unsigned((8'hbf));
    end
  assign wire2300 = reg2267[(3'h6):(1'h0)];
  always
    @(posedge clk) begin
      reg2301 <= ((~{reg2295, (|$signed(reg2282))}) << reg2277);
    end
  assign wire2302 = (7'h40);
  assign wire2303 = (8'hbe);
  always
    @(posedge clk) begin
      reg2304 <= wire2303;
      reg2305 <= (!({(reg2282 <<< reg2292), reg2270} ?
          $signed(((reg2282 ?
              reg2267 : wire2259) >= reg2270)) : reg2298[(3'h6):(3'h6)]));
      reg2306 <= {wire2259,
          ({reg2304} ?
              (((~&reg2294) < (reg2271 ?
                  reg2305 : wire2290)) == forvar2293) : reg2292[(3'h4):(2'h2)])};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2229
#( parameter param2250 = (~&((8'ha7) ? (8'hb3) : ((~|((7'h44) ^ (8'ha1))) ^~ (((8'hb0) ? (8'h9d) : (8'ha3)) ? ((7'h44) ? (8'hba) : (8'ha0)) : ((8'hb1) && (8'h9d))))))
, parameter param2251 = (param2250 ? param2250 : (((~&(param2250 ? (8'h9e) : param2250)) ? param2250 : ((param2250 << param2250) ? (param2250 ? (8'ha4) : param2250) : (|param2250))) ? (((~&param2250) ? (param2250 ? param2250 : (8'ha9)) : (8'ha9)) ? (((8'ha8) - param2250) ? (~param2250) : ((8'hac) ? param2250 : param2250)) : (8'h9e)) : ({(^~param2250), (8'hb6)} ^ param2250))) )
(y, clk, wire2233, wire2232, wire2231, wire2230);
  output wire [(32'h7c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire2233;
  input wire [(2'h3):(1'h0)] wire2232;
  input wire signed [(4'ha):(1'h0)] wire2231;
  input wire signed [(3'h6):(1'h0)] wire2230;
  reg [(4'ha):(1'h0)] reg2249 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2248 = (1'h0);
  reg [(5'h12):(1'h0)] reg2247 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2246 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire2245;
  reg [(5'h14):(1'h0)] reg2244 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2243 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2242 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2241 = (1'h0);
  reg [(4'h8):(1'h0)] reg2240 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2239 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2238 = (1'h0);
  reg [(3'h4):(1'h0)] reg2237 = (1'h0);
  reg [(2'h3):(1'h0)] reg2236 = (1'h0);
  reg [(2'h2):(1'h0)] reg2235 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire2234;
  assign y = {reg2249,
                 reg2248,
                 reg2247,
                 reg2246,
                 wire2245,
                 reg2244,
                 forvar2243,
                 forvar2242,
                 reg2241,
                 reg2240,
                 reg2239,
                 reg2238,
                 reg2237,
                 reg2236,
                 reg2235,
                 wire2234,
                 (1'h0)};
  assign wire2234 = wire2233;
  always
    @(posedge clk) begin
      reg2235 <= wire2233[(5'h12):(4'hd)];
      reg2236 <= (~^reg2235);
    end
  always
    @(posedge clk) begin
      reg2237 <= $signed(wire2233[(3'h5):(2'h2)]);
      reg2238 <= ((+$signed({$signed((7'h40))})) ?
          (~^($unsigned($unsigned(wire2233)) | $signed((reg2236 ?
              wire2233 : wire2231)))) : {(7'h43)});
      reg2239 <= wire2230[(1'h1):(1'h0)];
      reg2240 = (&$unsigned(($unsigned($signed(reg2239)) - ((wire2231 - reg2235) ?
          wire2232[(1'h1):(1'h0)] : wire2233[(4'hf):(3'h4)]))));
    end
  always
    @(posedge clk) begin
      reg2241 = reg2240[(1'h0):(1'h0)];
      for (forvar2242 = (1'h0); (forvar2242 < (1'h1)); forvar2242 = (forvar2242 + (1'h1)))
        begin
          for (forvar2243 = (1'h0); (forvar2243 < (1'h1)); forvar2243 = (forvar2243 + (1'h1)))
            begin
              reg2244 <= $signed((|(~$signed($signed(wire2230)))));
            end
        end
    end
  assign wire2245 = $signed((({reg2241, (^forvar2243)} ?
                        $unsigned((|reg2237)) : $unsigned((reg2244 ?
                            forvar2242 : reg2244))) >> $signed(forvar2242)));
  always
    @(posedge clk) begin
      reg2246 <= ((forvar2242[(3'h4):(2'h3)] ?
          reg2238 : $unsigned({$unsigned(wire2234),
              (wire2232 >>> reg2237)})) || (-$signed($unsigned(reg2236[(2'h3):(1'h0)]))));
      reg2247 <= reg2236;
    end
  always
    @(posedge clk) begin
      reg2248 <= reg2241;
      reg2249 <= ((^$signed(reg2238)) - (!(~$signed($signed(reg2239)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2186
#( parameter param2226 = ((((^((8'hbc) ? (8'hb2) : (8'hb1))) ? ((~^(8'hb8)) != ((8'h9f) < (8'hb2))) : (~&{(8'ha4)})) ? ((((8'hb2) ~^ (8'h9f)) >= {(8'ha1)}) ? (~((8'hbe) ? (8'hb4) : (8'hab))) : {(+(8'hbe))}) : {((^(8'hb5)) | (~(8'haa))), ((~^(7'h44)) ? {(8'haf), (8'hb9)} : (~&(7'h43)))}) ? ((|(((8'hb9) ? (8'hb4) : (8'ha7)) ? ((8'hba) ? (8'hb5) : (8'hb9)) : ((8'ha4) ? (8'had) : (8'ha7)))) ? (((~|(8'h9d)) ^ (~^(8'ha5))) >>> (8'ha2)) : ((((8'hbe) ? (8'ha2) : (8'h9c)) ? {(8'ha1)} : (+(8'hbe))) & ((+(8'had)) ? ((8'hb7) != (8'ha0)) : ((8'ha0) ? (8'hb4) : (8'ha9))))) : {(((^(8'haa)) == ((8'ha6) ^ (8'ha0))) ? (((8'hb3) < (7'h40)) <<< ((8'hbf) ? (8'ha3) : (8'h9c))) : (((8'h9e) | (8'haa)) & ((7'h44) ^~ (8'hb5)))), (((8'ha1) ? ((8'hb1) <<< (8'hb2)) : (~&(8'ha8))) ? (((8'hbe) <= (8'hba)) ? {(8'ha5)} : {(7'h40), (8'ha5)}) : ((~(8'ha5)) <<< ((8'hbb) | (8'hbf))))}) )
(y, clk, wire2190, wire2189, wire2188, wire2187);
  output wire [(32'h179):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire2190;
  input wire [(5'h11):(1'h0)] wire2189;
  input wire [(3'h6):(1'h0)] wire2188;
  input wire [(4'h9):(1'h0)] wire2187;
  wire [(4'hd):(1'h0)] wire2225;
  reg signed [(5'h11):(1'h0)] reg2224 = (1'h0);
  wire [(5'h14):(1'h0)] wire2223;
  reg signed [(5'h15):(1'h0)] reg2222 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2221 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2220 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2219 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire2218;
  wire [(2'h3):(1'h0)] wire2217;
  wire [(5'h14):(1'h0)] wire2216;
  reg signed [(2'h2):(1'h0)] reg2215 = (1'h0);
  reg [(2'h2):(1'h0)] reg2214 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2213 = (1'h0);
  reg [(4'h9):(1'h0)] reg2212 = (1'h0);
  wire [(4'ha):(1'h0)] wire2211;
  wire [(4'hf):(1'h0)] wire2210;
  reg signed [(2'h3):(1'h0)] reg2209 = (1'h0);
  reg [(2'h3):(1'h0)] reg2208 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2207 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2206 = (1'h0);
  reg [(5'h14):(1'h0)] reg2205 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2204 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2203 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2202 = (1'h0);
  reg [(5'h11):(1'h0)] reg2201 = (1'h0);
  reg [(2'h3):(1'h0)] reg2200 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2199 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2198 = (1'h0);
  reg [(4'hc):(1'h0)] reg2197 = (1'h0);
  wire [(4'ha):(1'h0)] wire2196;
  wire signed [(2'h2):(1'h0)] wire2195;
  wire signed [(2'h3):(1'h0)] wire2194;
  wire [(4'hf):(1'h0)] wire2193;
  wire signed [(3'h4):(1'h0)] wire2192;
  wire [(2'h2):(1'h0)] wire2191;
  assign y = {wire2225,
                 reg2224,
                 wire2223,
                 reg2222,
                 reg2221,
                 reg2220,
                 reg2219,
                 wire2218,
                 wire2217,
                 wire2216,
                 reg2215,
                 reg2214,
                 reg2213,
                 reg2212,
                 wire2211,
                 wire2210,
                 reg2209,
                 reg2208,
                 reg2207,
                 reg2206,
                 reg2205,
                 reg2204,
                 forvar2203,
                 reg2202,
                 reg2201,
                 reg2200,
                 reg2199,
                 forvar2198,
                 reg2197,
                 wire2196,
                 wire2195,
                 wire2194,
                 wire2193,
                 wire2192,
                 wire2191,
                 (1'h0)};
  assign wire2191 = wire2187[(3'h5):(2'h2)];
  assign wire2192 = (7'h44);
  assign wire2193 = $signed(wire2189);
  assign wire2194 = (((~&wire2192[(3'h4):(2'h3)]) > $unsigned(wire2191)) ?
                        wire2190 : ($signed(wire2190) ?
                            ({(&wire2192),
                                ((8'h9f) | wire2190)} - ($signed(wire2193) && (~(8'hae)))) : {wire2190}));
  assign wire2195 = (+$unsigned($signed((wire2192[(3'h4):(1'h1)] * $unsigned(wire2194)))));
  assign wire2196 = $signed($unsigned($signed($unsigned(wire2191))));
  always
    @(posedge clk) begin
      reg2197 = $unsigned($signed((&wire2187[(3'h5):(2'h2)])));
      for (forvar2198 = (1'h0); (forvar2198 < (2'h3)); forvar2198 = (forvar2198 + (1'h1)))
        begin
          reg2199 <= {(8'had)};
          reg2200 = ((!((~$unsigned(wire2196)) == wire2194[(2'h2):(1'h1)])) != (-{((wire2193 != wire2196) >> (wire2189 ?
                  wire2188 : reg2197))}));
          reg2201 <= wire2188[(3'h5):(2'h3)];
          reg2202 = (((^(~|reg2201[(3'h6):(3'h4)])) ?
              ($signed($signed(reg2199)) ?
                  ((reg2199 || reg2200) ^ (!(8'ha3))) : (~&(wire2195 || wire2190))) : (-$unsigned((wire2191 >= wire2193)))) <<< reg2200);
          for (forvar2203 = (1'h0); (forvar2203 < (2'h3)); forvar2203 = (forvar2203 + (1'h1)))
            begin
              reg2204 = (~|{wire2188[(2'h2):(1'h0)]});
              reg2205 <= wire2193;
              reg2206 = reg2205[(3'h4):(2'h3)];
              reg2207 <= ($signed(((wire2192[(2'h2):(1'h0)] << $signed(reg2200)) ?
                      wire2196[(2'h3):(1'h0)] : reg2202)) ?
                  wire2191 : forvar2198[(1'h0):(1'h0)]);
            end
        end
      reg2208 <= ($unsigned((forvar2203[(1'h0):(1'h0)] ~^ (-$signed(wire2189)))) ~^ $unsigned(((-reg2201[(5'h11):(3'h6)]) ?
          ((reg2207 << wire2192) ~^ reg2205[(4'hb):(4'h9)]) : ((reg2202 != wire2192) ~^ {wire2194}))));
      reg2209 <= $unsigned((~|(reg2199[(3'h7):(3'h6)] + reg2207[(3'h7):(3'h6)])));
    end
  assign wire2210 = reg2201[(2'h3):(1'h0)];
  assign wire2211 = wire2192;
  always
    @(posedge clk) begin
      reg2212 <= $unsigned(wire2195[(1'h1):(1'h1)]);
      reg2213 <= $unsigned(forvar2203);
    end
  always
    @(posedge clk) begin
      reg2214 = ((!(reg2202 >>> $unsigned($unsigned(wire2195)))) ?
          {$unsigned(wire2193),
              (({(8'ha0)} ? (~wire2194) : $signed(reg2208)) ?
                  reg2213 : $unsigned((~^wire2192)))} : ({((wire2191 ?
                          reg2206 : reg2204) ?
                      $signed((8'ha0)) : reg2200[(2'h2):(1'h0)]),
                  (forvar2203 ?
                      (wire2194 ? reg2206 : reg2200) : {wire2191, (8'ha2)})} ?
              reg2202[(1'h0):(1'h0)] : ($signed($unsigned(wire2195)) ?
                  reg2207[(1'h0):(1'h0)] : (|(wire2190 && reg2199)))));
      reg2215 <= reg2199;
    end
  assign wire2216 = ((~&reg2205[(4'hf):(3'h7)]) ?
                        forvar2198[(2'h2):(2'h2)] : wire2187[(3'h4):(1'h0)]);
  assign wire2217 = ((((7'h44) << (((8'ha2) < reg2201) ?
                            $unsigned(wire2192) : $signed(wire2187))) ?
                        {(((8'hb4) ? (7'h44) : (8'hbd)) - wire2190),
                            (^forvar2198)} : $signed({$signed(wire2216),
                            (reg2204 + forvar2198)})) >>> wire2193);
  assign wire2218 = reg2214;
  always
    @(posedge clk) begin
      reg2219 = $unsigned(((reg2215[(1'h0):(1'h0)] ?
          (-(wire2192 ?
              reg2208 : reg2202)) : ($signed(wire2217) - wire2196)) << $unsigned(((wire2188 ?
              (8'hae) : reg2200) ?
          $unsigned(reg2204) : $signed(reg2215)))));
      reg2220 <= wire2217;
      reg2221 = {($unsigned(($unsigned(reg2201) ?
              (^reg2214) : (reg2209 ? reg2207 : reg2202))) & $signed(reg2212)),
          forvar2198};
    end
  always
    @(posedge clk) begin
      reg2222 <= ({(wire2190[(3'h4):(2'h3)] ?
                  $unsigned(reg2220[(1'h0):(1'h0)]) : (8'hab))} ?
          wire2193 : $unsigned({(wire2192 ?
                  (reg2215 & wire2190) : $unsigned(wire2218)),
              reg2202[(3'h4):(3'h4)]}));
    end
  assign wire2223 = (wire2192 ~^ $unsigned({(+{wire2196, reg2213})}));
  always
    @(posedge clk) begin
      reg2224 <= (reg2212[(4'h9):(2'h3)] ?
          (wire2194 ?
              $unsigned((-(~|wire2187))) : (({(8'h9f), wire2223} ?
                      $unsigned((8'hbd)) : $signed(wire2191)) ?
                  wire2196 : ($signed((8'ha7)) ?
                      reg2219 : (|(8'hb7))))) : (wire2193 ?
              (reg2222[(1'h0):(1'h0)] ?
                  ($unsigned(reg2212) != wire2196[(3'h5):(2'h2)]) : reg2199[(4'hf):(4'h8)]) : (|$signed((+(7'h43))))));
    end
  assign wire2225 = ({wire2223[(4'ha):(1'h0)],
                        (((wire2190 ? reg2209 : reg2197) + $unsigned(reg2205)) ?
                            $unsigned(((8'ha2) || wire2218)) : reg2200[(2'h2):(1'h1)])} & (-(wire2223[(3'h4):(3'h4)] > reg2222)));
endmodule