(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h55f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire4;
  input wire [(5'h13):(1'h0)] wire3;
  input wire [(4'he):(1'h0)] wire2;
  input wire signed [(4'hd):(1'h0)] wire1;
  input wire signed [(5'h14):(1'h0)] wire0;
  wire signed [(3'h6):(1'h0)] wire927;
  reg signed [(2'h2):(1'h0)] reg122 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg121 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg120 = (1'h0);
  reg [(4'hb):(1'h0)] reg119 = (1'h0);
  reg [(3'h6):(1'h0)] reg118 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar117 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire116;
  wire [(3'h4):(1'h0)] wire115;
  reg signed [(3'h5):(1'h0)] reg114 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg113 = (1'h0);
  reg [(5'h12):(1'h0)] reg112 = (1'h0);
  reg [(5'h12):(1'h0)] reg111 = (1'h0);
  reg [(5'h12):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg108 = (1'h0);
  reg [(4'he):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg106 = (1'h0);
  reg [(3'h5):(1'h0)] reg105 = (1'h0);
  reg signed [(4'he):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar103 = (1'h0);
  reg [(4'h8):(1'h0)] reg102 = (1'h0);
  reg [(4'he):(1'h0)] reg101 = (1'h0);
  reg [(5'h17):(1'h0)] reg100 = (1'h0);
  reg [(5'h13):(1'h0)] reg99 = (1'h0);
  reg [(5'h14):(1'h0)] reg98 = (1'h0);
  reg [(4'he):(1'h0)] reg97 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg96 = (1'h0);
  reg [(4'hc):(1'h0)] forvar95 = (1'h0);
  reg [(4'h8):(1'h0)] reg94 = (1'h0);
  reg [(3'h7):(1'h0)] reg93 = (1'h0);
  reg [(3'h4):(1'h0)] reg92 = (1'h0);
  reg [(5'h15):(1'h0)] reg91 = (1'h0);
  reg [(4'hb):(1'h0)] reg90 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar89 = (1'h0);
  reg [(4'h8):(1'h0)] forvar88 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg87 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar86 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar85 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg84 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg83 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg82 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg81 = (1'h0);
  reg [(4'hc):(1'h0)] reg80 = (1'h0);
  reg [(5'h14):(1'h0)] reg79 = (1'h0);
  reg [(4'ha):(1'h0)] forvar78 = (1'h0);
  reg [(4'hd):(1'h0)] reg77 = (1'h0);
  reg [(3'h5):(1'h0)] forvar76 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg72 = (1'h0);
  reg signed [(4'he):(1'h0)] reg71 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar70 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar69 = (1'h0);
  reg [(4'hc):(1'h0)] reg68 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg67 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg66 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar65 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg64 = (1'h0);
  reg [(2'h2):(1'h0)] reg63 = (1'h0);
  reg [(4'h8):(1'h0)] forvar62 = (1'h0);
  reg [(4'h8):(1'h0)] reg61 = (1'h0);
  reg [(4'ha):(1'h0)] reg60 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar55 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg54 = (1'h0);
  reg [(2'h2):(1'h0)] reg53 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg52 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg51 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg50 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar49 = (1'h0);
  reg [(2'h3):(1'h0)] reg48 = (1'h0);
  reg [(2'h2):(1'h0)] reg47 = (1'h0);
  reg [(4'hc):(1'h0)] reg46 = (1'h0);
  reg [(5'h17):(1'h0)] reg45 = (1'h0);
  reg [(5'h10):(1'h0)] forvar44 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg43 = (1'h0);
  reg [(3'h7):(1'h0)] forvar42 = (1'h0);
  reg [(5'h13):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar40 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg39 = (1'h0);
  reg [(4'h8):(1'h0)] reg38 = (1'h0);
  reg [(4'hd):(1'h0)] reg37 = (1'h0);
  reg [(5'h10):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg35 = (1'h0);
  reg [(2'h3):(1'h0)] reg34 = (1'h0);
  reg [(2'h2):(1'h0)] reg33 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg32 = (1'h0);
  reg [(4'hd):(1'h0)] reg31 = (1'h0);
  reg [(4'h9):(1'h0)] reg30 = (1'h0);
  reg [(5'h10):(1'h0)] reg29 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg28 = (1'h0);
  reg [(5'h17):(1'h0)] reg27 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg26 = (1'h0);
  reg [(4'hd):(1'h0)] reg25 = (1'h0);
  reg [(3'h7):(1'h0)] forvar21 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg24 = (1'h0);
  reg [(3'h6):(1'h0)] reg23 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg22 = (1'h0);
  reg [(4'hd):(1'h0)] reg21 = (1'h0);
  reg [(5'h13):(1'h0)] reg20 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar19 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg17 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg16 = (1'h0);
  reg [(2'h2):(1'h0)] reg15 = (1'h0);
  reg [(4'h9):(1'h0)] reg14 = (1'h0);
  reg [(3'h4):(1'h0)] reg13 = (1'h0);
  reg [(4'hb):(1'h0)] reg12 = (1'h0);
  reg [(2'h3):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg10 = (1'h0);
  reg [(4'h8):(1'h0)] forvar9 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar8 = (1'h0);
  reg [(5'h15):(1'h0)] reg7 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6 = (1'h0);
  reg [(5'h12):(1'h0)] forvar5 = (1'h0);
  assign y = {wire927,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 forvar117,
                 wire116,
                 wire115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 forvar103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 forvar95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 forvar89,
                 forvar88,
                 reg87,
                 forvar86,
                 forvar85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 forvar78,
                 reg77,
                 forvar76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 forvar70,
                 forvar69,
                 reg68,
                 reg67,
                 reg66,
                 forvar65,
                 reg64,
                 reg63,
                 forvar62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 forvar55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 forvar49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 forvar44,
                 reg43,
                 forvar42,
                 reg41,
                 forvar40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 forvar21,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 forvar19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 forvar9,
                 forvar8,
                 reg7,
                 forvar6,
                 forvar5,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar5 = (1'h0); (forvar5 < (1'h0)); forvar5 = (forvar5 + (1'h1)))
        begin
          for (forvar6 = (1'h0); (forvar6 < (2'h2)); forvar6 = (forvar6 + (1'h1)))
            begin
              reg7 <= wire0[(2'h3):(1'h0)];
            end
          for (forvar8 = (1'h0); (forvar8 < (1'h1)); forvar8 = (forvar8 + (1'h1)))
            begin
              for (forvar9 = (1'h0); (forvar9 < (3'h4)); forvar9 = (forvar9 + (1'h1)))
                begin
                  reg10 <= forvar6;
                  reg11 <= ("riwPwp" | ("5sb3ZhNfwb" ?
                      (~^"J17VbeWrErBnS") : wire3[(3'h6):(2'h3)]));
                end
            end
          reg12 <= {(reg11[(1'h0):(1'h0)] ?
                  (^$signed(wire4[(4'h9):(4'h9)])) : forvar5)};
          reg13 <= (($unsigned(wire4) ?
              {wire2[(3'h7):(3'h7)], $signed($signed(reg7))} : ((-(~&reg10)) ?
                  ($unsigned(wire3) | $signed(wire3)) : (!$unsigned(forvar6)))) ~^ (($unsigned((~&reg12)) ?
              $signed(reg10) : forvar6[(1'h1):(1'h0)]) + (8'h9f)));
        end
    end
  always
    @(posedge clk) begin
      reg14 = {$unsigned((~&{"vfnHH8bHekCiFHnKy", (reg12 || reg11)}))};
      reg15 = ((($signed(forvar5[(4'hd):(3'h5)]) << wire4[(3'h7):(1'h1)]) ?
              (((8'hbb) ? forvar9 : wire3[(3'h7):(1'h0)]) ?
                  $signed($signed(wire0)) : $signed((forvar6 ?
                      wire3 : reg13))) : (($signed(reg14) ?
                      $signed(forvar8) : (wire2 ? reg13 : reg7)) ?
                  "rC3qhS" : ((wire2 ? forvar9 : reg10) ?
                      "VylUJ2AN" : (reg13 ? forvar6 : forvar6)))) ?
          (($unsigned(reg10[(4'he):(3'h5)]) ~^ $signed((^~reg10))) ?
              {{(^wire4), (reg12 ? reg7 : wire3)},
                  (!"6pGhr")} : reg7[(2'h2):(2'h2)]) : "Ks5");
      reg16 <= {("KE" < "PwrWuEZEaXZ")};
    end
  always
    @(posedge clk) begin
      reg17 <= reg11[(1'h1):(1'h0)];
      reg18 <= wire1;
    end
  always
    @(posedge clk) begin
      for (forvar19 = (1'h0); (forvar19 < (3'h4)); forvar19 = (forvar19 + (1'h1)))
        begin
          if ((reg17 * ($unsigned({$unsigned(reg10),
              (~reg12)}) >>> ({(forvar8 ~^ reg16),
              wire1[(4'hc):(2'h3)]} ~^ $signed(forvar5)))))
            begin
              reg20 <= "uTJQYiPXXQ6rXfzcSy";
              reg21 <= $unsigned(wire4[(4'h9):(3'h6)]);
              reg22 <= ((~&$signed(("6k8i8r8tfdYJHX5GiZ" ?
                      wire0 : "0FRxmXdPRMsEvhiWs0f"))) ?
                  (&{{reg18}, (^~$unsigned((8'h9e)))}) : $signed(reg17));
              reg23 <= $unsigned(forvar19);
              reg24 = wire0[(3'h7):(1'h1)];
            end
          else
            begin
              reg20 <= reg12;
              if (((~|{(~|(reg20 << reg16)), (forvar9 != ((8'h9c) > wire0))}) ?
                  $unsigned(({{forvar19},
                      reg15} * reg20[(4'h9):(4'h8)])) : ($unsigned(reg20[(4'ha):(4'ha)]) ?
                      wire3 : reg11[(2'h2):(1'h1)])))
                begin
                  for (forvar21 = (1'h0); (forvar21 < (1'h0)); forvar21 = (forvar21 + (1'h1)))
                    begin
                      reg22 <= (wire0[(4'h9):(4'h8)] ?
                          $signed(wire3[(1'h1):(1'h0)]) : "82WbKnlCaWZ");
                      reg23 = reg20;
                      reg24 <= forvar5[(1'h1):(1'h1)];
                      reg25 = $unsigned((^wire1[(4'hb):(2'h3)]));
                      reg26 <= (("aX1S" ^ ($signed($unsigned(wire0)) ?
                              ({reg15} || $signed((8'ha9))) : {$signed(forvar21),
                                  $unsigned(reg21)})) ?
                          {(reg7 && "Ihi0Tz8tXtNqW5Uw"),
                              (wire4 + {$unsigned((7'h48))})} : ($signed(("ePCxqV09paXIiFA5VKb2" <<< reg17)) ?
                              {$signed($unsigned(forvar9)),
                                  $signed(((8'hbc) - wire0))} : {(forvar19 ?
                                      $signed(reg24) : (wire4 != forvar5)),
                                  ($unsigned(reg25) - (^reg12))}));
                    end
                  reg27 <= $unsigned($unsigned(((~|(~&wire2)) ^~ forvar21)));
                  reg28 = $unsigned($signed($unsigned((^~(|forvar6)))));
                  reg29 = (reg24[(2'h3):(2'h2)] >>> (wire2[(4'hd):(1'h1)] >= (reg15 ?
                      ($signed((8'hab)) ? reg21 : $unsigned(wire4)) : reg17)));
                end
              else
                begin
                  reg21 <= $signed($unsigned(reg17));
                end
              reg30 = ($signed(reg7) >>> $unsigned((|(|(!reg27)))));
              reg31 <= (^forvar19);
            end
          reg32 = (("WO" <= "A") ?
              ((forvar9[(3'h6):(3'h6)] + {$signed(wire3)}) && "0eQQ8VTfYxzz3VDUR") : $signed(($signed((8'hbe)) ^ reg26)));
          reg33 <= {reg10[(3'h6):(2'h2)], reg18};
          reg34 = "IrVdbSw3AlDNo5W";
        end
      reg35 = "8vIGB9eb99xbwPvW";
      reg36 <= $unsigned((($signed(reg14[(2'h2):(1'h0)]) - ("RallC5lASQnSG6t7" - (^reg34))) >= ($unsigned($unsigned(reg15)) ?
          $signed($signed(reg14)) : reg24[(3'h4):(2'h3)])));
      reg37 <= reg10[(4'h8):(1'h1)];
      reg38 <= $signed($unsigned($unsigned({$unsigned((8'hab))})));
    end
  always
    @(posedge clk) begin
      reg39 = (-("BtMh" ?
          (($signed(reg14) ? (^wire2) : $signed(forvar21)) >>> "0C9") : "UrP"));
      for (forvar40 = (1'h0); (forvar40 < (3'h4)); forvar40 = (forvar40 + (1'h1)))
        begin
          reg41 = (reg23[(2'h2):(1'h1)] >>> (8'hb0));
          for (forvar42 = (1'h0); (forvar42 < (2'h3)); forvar42 = (forvar42 + (1'h1)))
            begin
              reg43 = reg39;
              for (forvar44 = (1'h0); (forvar44 < (1'h1)); forvar44 = (forvar44 + (1'h1)))
                begin
                  reg45 = $signed((reg36[(3'h4):(1'h0)] * (-$signed("z3MbGT"))));
                  reg46 <= (~("3XGT92r5u" ~^ (8'hb9)));
                  reg47 <= forvar8;
                  reg48 = "kbXQ8RkaYp4m";
                  for (forvar49 = (1'h0); (forvar49 < (3'h4)); forvar49 = (forvar49 + (1'h1)))
                    begin
                      reg50 <= $signed((reg24 ?
                          {(forvar42 <= (^~reg46)),
                              wire3[(1'h1):(1'h1)]} : reg15[(2'h2):(2'h2)]));
                      reg51 <= (~^$signed(reg16[(1'h1):(1'h1)]));
                      reg52 = reg30[(1'h1):(1'h0)];
                      reg53 <= {((|reg46) * (|"kO7Lz5VUGkpi"))};
                      reg54 <= $signed($signed(((8'hb5) ?
                          reg13[(2'h3):(1'h1)] : (reg45 ?
                              "Ro0AaBPui0OPhtUvVYq" : $signed(reg28)))));
                    end
                end
            end
          for (forvar55 = (1'h0); (forvar55 < (3'h4)); forvar55 = (forvar55 + (1'h1)))
            begin
              reg56 <= (|wire1);
              reg57 <= $signed("gYBXvmY");
              reg58 <= $unsigned({("pO0oB37CkzwyBom6" ?
                      $unsigned($unsigned(reg14)) : forvar5),
                  reg7});
              reg59 <= {$signed(reg12[(4'ha):(1'h1)])};
              reg60 <= (!({$unsigned(reg21)} ?
                  (-(~&"NgawVYZHx98pqMAsXUngm")) : (+"FRDyXtfawMvVKPMmROS")));
            end
          reg61 = "Y12";
        end
      for (forvar62 = (1'h0); (forvar62 < (3'h4)); forvar62 = (forvar62 + (1'h1)))
        begin
          reg63 <= forvar5;
          reg64 <= $signed((^~forvar9));
          for (forvar65 = (1'h0); (forvar65 < (1'h0)); forvar65 = (forvar65 + (1'h1)))
            begin
              reg66 = $signed(reg39);
              reg67 <= "w10ASCIRx4UFG5hlvKmBm";
              reg68 <= forvar49;
              for (forvar69 = (1'h0); (forvar69 < (1'h0)); forvar69 = (forvar69 + (1'h1)))
                begin
                  for (forvar70 = (1'h0); (forvar70 < (1'h0)); forvar70 = (forvar70 + (1'h1)))
                    begin
                      reg71 <= reg35;
                      reg72 = ((8'hb8) < (^"nGJv"));
                    end
                  reg73 = reg20;
                end
            end
        end
    end
  always
    @(posedge clk) begin
      reg74 <= (^{$signed($signed((^~forvar62)))});
      reg75 <= reg28[(5'h14):(1'h1)];
      for (forvar76 = (1'h0); (forvar76 < (1'h1)); forvar76 = (forvar76 + (1'h1)))
        begin
          reg77 <= $unsigned((reg23[(2'h2):(2'h2)] & (+$unsigned((reg53 ?
              reg17 : reg61)))));
        end
      for (forvar78 = (1'h0); (forvar78 < (1'h1)); forvar78 = (forvar78 + (1'h1)))
        begin
          reg79 = ($signed($signed($unsigned((forvar78 - (7'h44))))) ?
              (7'h46) : (8'hb2));
          reg80 <= (({"gg2PL19gpS", "c9Ugdl2rhKPo4Zw"} ?
                  "yv7uzJQcdW9" : reg29[(4'ha):(3'h7)]) ?
              (8'hb5) : {reg26});
          reg81 <= reg37[(1'h0):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      reg82 <= $unsigned(({((reg64 <<< reg29) ?
              $unsigned(forvar55) : (reg73 ?
                  forvar8 : reg12))} >> (+reg48[(2'h3):(1'h1)])));
      reg83 = $signed($unsigned((8'hb1)));
      reg84 <= (&reg52[(4'he):(4'ha)]);
      for (forvar85 = (1'h0); (forvar85 < (2'h3)); forvar85 = (forvar85 + (1'h1)))
        begin
          for (forvar86 = (1'h0); (forvar86 < (3'h4)); forvar86 = (forvar86 + (1'h1)))
            begin
              reg87 <= ($unsigned({$signed($unsigned(reg81))}) ?
                  $signed("fz4SIrRSuFLuqlTKfkYXL") : ($signed(($unsigned(wire4) | {reg35,
                          forvar69})) ?
                      $unsigned($unsigned((reg54 ?
                          reg34 : reg77))) : ($unsigned((forvar69 ?
                              wire0 : reg16)) ?
                          (forvar76[(2'h3):(1'h1)] ?
                              {reg75} : $signed(forvar86)) : (((7'h43) ?
                                  reg63 : reg63) ?
                              forvar62 : $unsigned(reg15)))));
              for (forvar88 = (1'h0); (forvar88 < (2'h2)); forvar88 = (forvar88 + (1'h1)))
                begin
                  for (forvar89 = (1'h0); (forvar89 < (2'h2)); forvar89 = (forvar89 + (1'h1)))
                    begin
                      reg90 <= (reg13[(3'h4):(1'h1)] < wire2[(3'h7):(1'h0)]);
                      reg91 = ((~^((reg15 >>> $signed(reg37)) >> $unsigned($unsigned((8'ha1))))) ?
                          {(($unsigned(wire1) * {reg27}) ~^ $signed((&reg34)))} : $signed(reg56[(4'h9):(3'h7)]));
                      reg92 = (reg72[(5'h10):(4'hd)] || forvar9[(3'h4):(1'h0)]);
                      reg93 <= "lfNZRJ19Oln7A0EqQNF";
                      reg94 = reg48;
                    end
                end
            end
          for (forvar95 = (1'h0); (forvar95 < (1'h1)); forvar95 = (forvar95 + (1'h1)))
            begin
              reg96 <= (~&reg90);
              reg97 <= (reg54 ? $signed(reg45) : reg80);
            end
          reg98 <= reg52;
          reg99 = $unsigned({{(forvar55[(4'hb):(4'h9)] ?
                      (reg77 ? (8'haa) : reg73) : ((8'ha0) << reg16))},
              $signed("NZNqaHxxp9ihdw")});
        end
    end
  always
    @(posedge clk) begin
      reg100 <= ($signed(reg13[(1'h0):(1'h0)]) ?
          reg43 : $unsigned(("0ee3y15779" ~^ ((~|forvar5) >= $unsigned(forvar9)))));
      reg101 = (^~((reg81 >= ((!reg66) ?
          $signed((8'hb2)) : (forvar44 <<< (8'hbf)))) ~^ forvar86[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg102 <= (~&((reg21 ?
              (reg12 ? "r2lAaWI" : forvar86) : $unsigned("NFUe")) ?
          (reg74[(5'h11):(4'ha)] - (^(8'ha1))) : "lvnMLtnGJX"));
      for (forvar103 = (1'h0); (forvar103 < (2'h2)); forvar103 = (forvar103 + (1'h1)))
        begin
          reg104 <= (~&("h21" & (|$unsigned("Zw1De"))));
          reg105 = reg94;
          reg106 = (~|reg67);
        end
    end
  always
    @(posedge clk) begin
      if (reg59)
        begin
          reg107 = ((("EfyLQ0lL9A4qK7o" ~^ wire2) ?
              ("cleY77oSbTiJTCBitJxS" ?
                  ($signed(reg84) >>> wire1) : reg99[(4'ha):(3'h7)]) : (wire0 + $signed(wire3))) ^ reg82);
          reg108 <= "M";
          reg109 <= $unsigned($signed(reg11));
          reg110 = (forvar76 ?
              (~&$unsigned(({reg100, forvar21} ?
                  {(8'ha3),
                      (7'h43)} : (~reg39)))) : $signed(reg106[(3'h5):(2'h2)]));
          reg111 <= $unsigned((^reg99));
        end
      else
        begin
          reg107 = "caSXKahMzeadx";
          reg108 <= {(~^($signed(((7'h44) ~^ forvar5)) ?
                  $signed((reg54 ? reg99 : reg56)) : $signed((forvar85 ?
                      reg53 : (7'h40)))))};
          reg109 <= (8'h9c);
          reg110 <= $unsigned(("I41MyNxmn" ~^ (|reg26)));
          reg111 <= {{("Dud" ?
                      ((reg43 ? (8'h9f) : reg92) >> (forvar21 ?
                          reg79 : forvar69)) : reg71[(4'hc):(4'hb)])}};
        end
      reg112 = "GtvkrnVogPvqUs0CgbT";
      reg113 <= "YVdB0b";
      reg114 = reg18;
    end
  assign wire115 = $signed({(~|wire3), reg87});
  assign wire116 = {($signed(reg92) ~^ ("M9cvsMOtHOa" ?
                           (-((8'hac) | reg113)) : reg59)),
                       "xffn7cMh2TET0xcbkm"};
  always
    @(posedge clk) begin
      for (forvar117 = (1'h0); (forvar117 < (2'h3)); forvar117 = (forvar117 + (1'h1)))
        begin
          reg118 <= reg59[(1'h1):(1'h0)];
        end
      reg119 <= ({$signed((~&$unsigned(reg22)))} >>> reg97);
      reg120 <= reg17[(2'h3):(1'h0)];
      reg121 <= (!((reg101[(2'h2):(1'h1)] ? ((^~reg79) | {reg77}) : reg82) ?
          {$unsigned((reg113 ? forvar6 : reg84)),
              (^~(reg87 ? forvar95 : reg39))} : ("sKJN" ?
              (!$unsigned(reg97)) : $unsigned($signed(reg11)))));
    end
  always
    @(posedge clk) begin
      reg122 <= (~^$unsigned("o1ZtEE"));
    end
  module123 modinst928 (.wire127(reg23), .y(wire927), .wire125(reg26), .clk(clk), .wire126(reg58), .wire124(reg108));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module123  (y, clk, wire124, wire125, wire126, wire127);
  output wire [(32'h401):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire124;
  input wire signed [(4'hc):(1'h0)] wire125;
  input wire signed [(5'h15):(1'h0)] wire126;
  input wire signed [(3'h6):(1'h0)] wire127;
  reg [(5'h10):(1'h0)] reg926 = (1'h0);
  reg [(3'h4):(1'h0)] reg925 = (1'h0);
  reg signed [(4'he):(1'h0)] reg924 = (1'h0);
  reg [(3'h6):(1'h0)] reg923 = (1'h0);
  reg [(4'h8):(1'h0)] reg922 = (1'h0);
  reg [(5'h12):(1'h0)] reg921 = (1'h0);
  reg [(4'hc):(1'h0)] reg920 = (1'h0);
  reg [(3'h6):(1'h0)] reg919 = (1'h0);
  reg [(3'h5):(1'h0)] reg918 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar917 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar916 = (1'h0);
  reg [(3'h7):(1'h0)] reg915 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg914 = (1'h0);
  reg [(4'h8):(1'h0)] reg913 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar912 = (1'h0);
  reg [(3'h7):(1'h0)] reg911 = (1'h0);
  reg [(5'h10):(1'h0)] forvar910 = (1'h0);
  reg [(4'hd):(1'h0)] reg909 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg908 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg907 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar906 = (1'h0);
  reg [(4'hd):(1'h0)] forvar905 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg904 = (1'h0);
  reg [(4'ha):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg902 = (1'h0);
  reg [(2'h2):(1'h0)] reg901 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire900;
  reg signed [(4'hd):(1'h0)] reg899 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg898 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg128 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg129 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg130 = (1'h0);
  reg [(5'h15):(1'h0)] reg131 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg132 = (1'h0);
  reg [(5'h12):(1'h0)] forvar133 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg135 = (1'h0);
  reg [(5'h11):(1'h0)] reg136 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar137 = (1'h0);
  reg [(5'h16):(1'h0)] forvar138 = (1'h0);
  reg [(4'he):(1'h0)] reg139 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg140 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg141 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar142 = (1'h0);
  reg [(4'hc):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg144 = (1'h0);
  reg [(4'hc):(1'h0)] reg145 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg146 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg147 = (1'h0);
  reg [(5'h15):(1'h0)] reg148 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg149 = (1'h0);
  reg [(4'hc):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar151 = (1'h0);
  reg [(2'h2):(1'h0)] reg152 = (1'h0);
  reg [(5'h10):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg154 = (1'h0);
  reg [(5'h17):(1'h0)] reg155 = (1'h0);
  reg [(4'h9):(1'h0)] reg156 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg157 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg159 = (1'h0);
  wire [(5'h13):(1'h0)] wire160;
  reg signed [(5'h15):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg162 = (1'h0);
  reg [(5'h12):(1'h0)] reg163 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar164 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg165 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg166 = (1'h0);
  reg [(5'h10):(1'h0)] reg167 = (1'h0);
  reg [(5'h14):(1'h0)] reg168 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg169 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg170 = (1'h0);
  reg [(5'h15):(1'h0)] forvar171 = (1'h0);
  reg [(3'h6):(1'h0)] reg172 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg173 = (1'h0);
  reg [(5'h15):(1'h0)] reg174 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg176 = (1'h0);
  wire [(5'h10):(1'h0)] wire896;
  assign y = {reg926,
                 reg925,
                 reg924,
                 reg923,
                 reg922,
                 reg921,
                 reg920,
                 reg919,
                 reg918,
                 forvar917,
                 forvar916,
                 reg915,
                 reg914,
                 reg913,
                 forvar912,
                 reg911,
                 forvar910,
                 reg909,
                 reg908,
                 reg907,
                 forvar906,
                 forvar905,
                 reg904,
                 reg903,
                 reg902,
                 reg901,
                 wire900,
                 reg899,
                 reg898,
                 reg128,
                 reg129,
                 reg130,
                 reg131,
                 reg132,
                 forvar133,
                 reg134,
                 reg135,
                 reg136,
                 forvar137,
                 forvar138,
                 reg139,
                 reg140,
                 reg141,
                 forvar142,
                 reg143,
                 reg144,
                 reg145,
                 reg146,
                 reg147,
                 reg148,
                 reg149,
                 reg150,
                 forvar151,
                 reg152,
                 reg153,
                 reg154,
                 reg155,
                 reg156,
                 reg157,
                 reg158,
                 reg159,
                 wire160,
                 reg161,
                 reg162,
                 reg163,
                 forvar164,
                 reg165,
                 reg166,
                 reg167,
                 reg168,
                 reg169,
                 reg170,
                 forvar171,
                 reg172,
                 reg173,
                 reg174,
                 reg175,
                 reg176,
                 wire896,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg128 = (wire126[(4'hd):(3'h7)] ?
          (8'haf) : ((wire127[(3'h5):(3'h5)] - (~&{wire127,
              wire127})) | ((~|"") < "YQJD8PeH7RP3Cpo2J2UnR")));
      reg129 <= wire127[(3'h5):(3'h5)];
      reg130 <= ((8'ha6) ?
          (($signed((wire126 && wire125)) ?
                  ($signed(wire124) ?
                      wire127[(1'h1):(1'h0)] : $unsigned(wire126)) : "c4iAe1Ug2hIu") ?
              wire124 : ($signed($signed(wire126)) && $unsigned(reg129[(1'h1):(1'h0)]))) : ({("2XC" + {wire126,
                  (8'ha0)}),
              "9iVNGpY3KMdpMG"} * (("39AU1lgJTTMTsfIH7RfS" ?
                  $signed(reg129) : wire127) ?
              (~^"gcdnNgiL") : $unsigned($unsigned(wire125)))));
      reg131 = $signed(reg130[(2'h3):(2'h3)]);
      reg132 = $signed($signed(reg130));
    end
  always
    @(posedge clk) begin
      for (forvar133 = (1'h0); (forvar133 < (2'h3)); forvar133 = (forvar133 + (1'h1)))
        begin
          reg134 <= $signed("gKNvhGgE2PzCczakTHY");
        end
      reg135 = $unsigned({((^$unsigned(reg130)) ^ $unsigned("a4XO5piPSkokFk6AkMpR2U"))});
      if ($unsigned($unsigned((7'h44))))
        begin
          reg136 <= forvar133;
        end
      else
        begin
          reg136 <= forvar133[(1'h1):(1'h1)];
          for (forvar137 = (1'h0); (forvar137 < (2'h3)); forvar137 = (forvar137 + (1'h1)))
            begin
              for (forvar138 = (1'h0); (forvar138 < (3'h4)); forvar138 = (forvar138 + (1'h1)))
                begin
                  reg139 <= wire125;
                  reg140 = $signed({$signed({(~&wire125),
                          (reg129 != forvar138)})});
                  reg141 <= reg136[(4'hc):(3'h4)];
                end
              for (forvar142 = (1'h0); (forvar142 < (1'h0)); forvar142 = (forvar142 + (1'h1)))
                begin
                  reg143 <= "l9fbxY";
                  if (reg131[(4'ha):(2'h3)])
                    begin
                      reg144 <= wire124[(2'h2):(1'h0)];
                      reg145 <= ($unsigned(((~&reg129[(1'h1):(1'h1)]) ^~ $signed((forvar133 || reg144)))) - $unsigned(reg143[(3'h4):(2'h3)]));
                      reg146 <= (-($unsigned({reg141[(2'h3):(1'h0)]}) ~^ "Eh2K"));
                    end
                  else
                    begin
                      reg144 <= {reg146};
                      reg145 <= wire125;
                      reg146 <= ("CJnHilcZHKFnt7he" ?
                          {(((8'h9c) ~^ reg128) >>> $unsigned("CxEO1aE")),
                              reg129[(2'h3):(1'h1)]} : (("Rh8VVCJFWIcANkwog" | (reg130[(2'h3):(2'h2)] ?
                                  "B" : ((8'hae) & wire126))) ?
                              (^~(+{reg130})) : ((-(reg128 ?
                                  reg130 : reg132)) <= $signed(forvar137))));
                    end
                  reg147 <= reg132;
                  reg148 <= ($unsigned(($unsigned(reg145[(4'hc):(1'h0)]) & $signed("iMxudV97YZw8pVAUaF"))) <= {($unsigned((reg136 > (7'h43))) != "2iy9xVYSZhNtcQ"),
                      (reg139 ? reg128 : "J")});
                  reg149 <= $unsigned(("WrZse09tZn" ?
                      ({reg146, wire124} ?
                          (~&(reg130 ?
                              reg128 : reg147)) : reg140) : "whLEZ69rkiBpLo7QiBdC"));
                end
            end
          reg150 <= "";
          for (forvar151 = (1'h0); (forvar151 < (2'h3)); forvar151 = (forvar151 + (1'h1)))
            begin
              reg152 <= {"qcrwpLui0", "IrbEPIYeE3JgdXXlb"};
              reg153 = forvar133;
            end
        end
      reg154 = "kMLm8oAEJ";
      reg155 <= ("pqi9fOEAq" >>> "sMrh5UzHlnz8XGTHOGnL");
    end
  always
    @(posedge clk) begin
      reg156 <= (&("u" ~^ $signed("vARmV6rA")));
      reg157 = (reg150 ?
          (^((^~(reg135 ? reg130 : (7'h43))) ~^ ((reg152 * (8'hb5)) ?
              reg136[(3'h4):(1'h0)] : wire124))) : wire126[(2'h2):(1'h0)]);
      reg158 <= $unsigned(wire124[(2'h2):(1'h0)]);
      reg159 <= "UvDi03AL7H8yqF";
    end
  assign wire160 = (8'ha8);
  always
    @(posedge clk) begin
      reg161 <= (("Z" ?
              wire126 : ($unsigned($signed((8'ha1))) ?
                  (&"CnDl3OqAU9na3TNyyUUO") : reg156)) ?
          ((reg159[(4'h9):(3'h7)] >> reg149[(2'h2):(2'h2)]) ^ "FYmRdwN") : reg153);
      reg162 <= {((!((forvar151 ? forvar133 : reg154) ?
                  $signed(reg159) : (reg154 << reg129))) ?
              $unsigned(wire124[(1'h0):(1'h0)]) : ((8'hac) >= reg152))};
      reg163 = "";
    end
  always
    @(posedge clk) begin
      for (forvar164 = (1'h0); (forvar164 < (2'h2)); forvar164 = (forvar164 + (1'h1)))
        begin
          reg165 <= reg153[(3'h5):(3'h5)];
          reg166 <= {"0QrJhIsEY4uudECYMNP", "2ED"};
          reg167 <= (^~(($unsigned({forvar142}) ?
                  reg161[(4'he):(3'h7)] : (reg154 ?
                      (reg145 ? reg154 : reg134) : (-reg150))) ?
              $signed(reg150) : (($signed(reg128) ^~ "lzZnF0BnGGfBB6GcHhQ") > "loI")));
          reg168 <= ($unsigned("VM0") ?
              ($signed((~|reg154)) ^~ $signed(("yRgk4" ?
                  $signed(reg130) : $unsigned(reg163)))) : ($signed(((^forvar138) != (reg141 ?
                  reg132 : forvar142))) || $unsigned((^$unsigned(reg167)))));
          reg169 <= {$unsigned("WJnD7y9QHZmkotYUVHd"), "tslTkv0Yzmi"};
        end
      reg170 = $signed(({$unsigned($signed(reg168)), (~&reg136)} ?
          "NnKlvWMNqH8ZloVvu" : "399yRH0bxyonlUt"));
      for (forvar171 = (1'h0); (forvar171 < (2'h3)); forvar171 = (forvar171 + (1'h1)))
        begin
          reg172 = (^((+({reg154, reg149} <= reg131[(4'h8):(3'h4)])) ?
              ("crJ6ZMKDeni" <= (~&(reg141 ?
                  reg129 : reg152))) : $signed({(!reg130)})));
          reg173 <= {{$signed("6n2Egz36Ovy"), forvar142}};
          reg174 <= $signed("ZIVoUGJSKyh6IAGy4ZkOm");
          reg175 = "C4A9EWvrM0qXoHPWY9FTX";
        end
      reg176 = (wire125[(1'h0):(1'h0)] * $signed(reg169[(3'h5):(1'h0)]));
    end
  module177 modinst897 (wire896, clk, reg168, reg155, reg130, reg144, reg162);
  always
    @(posedge clk) begin
      reg898 <= $unsigned($signed(("46AorK5l16HVwV9rW6uqe" ?
          ("WDd9YJuasV4136iCi8" <= "") : forvar133)));
    end
  always
    @(posedge clk) begin
      reg899 <= $unsigned(reg168[(4'hb):(2'h2)]);
    end
  assign wire900 = ("" ? ({reg155} ~^ wire126) : reg158[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      reg901 <= "z1HaS3uo1";
      reg902 = reg135;
      reg903 <= (reg165 ? $signed(reg129[(2'h2):(1'h0)]) : reg136);
      reg904 = ($unsigned(((~|(reg132 >= (8'ha9))) || $signed(reg157))) ?
          $unsigned(forvar142) : {{$unsigned(((8'hb2) ? reg135 : (8'had)))}});
    end
  always
    @(posedge clk) begin
      for (forvar905 = (1'h0); (forvar905 < (2'h3)); forvar905 = (forvar905 + (1'h1)))
        begin
          for (forvar906 = (1'h0); (forvar906 < (3'h4)); forvar906 = (forvar906 + (1'h1)))
            begin
              reg907 <= {$unsigned($signed(((forvar133 ~^ reg159) ~^ reg155)))};
              reg908 = reg143[(1'h0):(1'h0)];
              reg909 = "wOA5oUPO";
              for (forvar910 = (1'h0); (forvar910 < (2'h2)); forvar910 = (forvar910 + (1'h1)))
                begin
                  reg911 <= reg175[(1'h1):(1'h0)];
                end
            end
          for (forvar912 = (1'h0); (forvar912 < (1'h0)); forvar912 = (forvar912 + (1'h1)))
            begin
              reg913 <= $unsigned(($unsigned(("m" ?
                      (^~reg156) : $signed(wire125))) ?
                  (reg155 ?
                      $unsigned($unsigned(reg136)) : reg908) : (reg157[(3'h5):(3'h4)] < {"wGcv4b"})));
              reg914 <= (|$signed(reg162[(4'he):(3'h7)]));
              reg915 <= reg145;
              for (forvar916 = (1'h0); (forvar916 < (2'h2)); forvar916 = (forvar916 + (1'h1)))
                begin
                  for (forvar917 = (1'h0); (forvar917 < (1'h0)); forvar917 = (forvar917 + (1'h1)))
                    begin
                      reg918 <= $unsigned($unsigned($signed(($unsigned(reg909) != {reg136,
                          reg150}))));
                    end
                  reg919 = $unsigned("Tt1o77xq");
                  reg920 <= reg161[(5'h13):(4'he)];
                  reg921 <= (reg919 ? "InUtOtNqGJc4wH" : (7'h47));
                  reg922 = reg170[(3'h5):(2'h3)];
                end
              reg923 <= (-(~&("XiZK9UNAEflb0" - $signed({wire900,
                  forvar905}))));
            end
        end
      reg924 <= "";
      reg925 <= $unsigned(($signed($unsigned("pwaSGogo")) | "dEYNPdomwdPhQUZtTSN"));
      reg926 <= {"VqSvD", wire124};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module177
#( parameter param894 = (((^({(8'h9e)} ? {(8'hb5)} : ((8'hb1) >> (8'hb5)))) ? (|({(8'haa)} ? (^(8'h9c)) : ((8'ha2) ? (7'h42) : (8'hb7)))) : (^~((^~(8'h9f)) * ((8'ha8) <= (8'hb2))))) ? (({(-(8'ha4)), ((7'h47) >> (8'h9d))} + {(-(8'hb6))}) & ((8'ha1) ? (^~(~^(8'hab))) : {(|(8'hab)), (~^(7'h47))})) : (^(~(~&((8'ha6) >>> (8'hb3))))))
, parameter param895 = {(((8'hbb) ? param894 : ((~param894) ? (~&(8'hb8)) : (~^param894))) || ({(param894 ? param894 : (7'h42)), {param894, param894}} ? {(param894 ? param894 : param894)} : {{param894, param894}})), param894} )
(y, clk, wire182, wire181, wire180, wire179, wire178);
  output wire [(32'h5ca):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire182;
  input wire signed [(5'h17):(1'h0)] wire181;
  input wire [(5'h15):(1'h0)] wire180;
  input wire signed [(4'hb):(1'h0)] wire179;
  input wire signed [(5'h11):(1'h0)] wire178;
  wire [(3'h6):(1'h0)] wire893;
  reg [(2'h3):(1'h0)] reg892 = (1'h0);
  reg [(5'h16):(1'h0)] reg891 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar890 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg889 = (1'h0);
  reg [(5'h14):(1'h0)] reg888 = (1'h0);
  reg [(5'h17):(1'h0)] reg887 = (1'h0);
  reg [(3'h6):(1'h0)] reg886 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar885 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg884 = (1'h0);
  reg [(2'h3):(1'h0)] reg883 = (1'h0);
  reg [(2'h3):(1'h0)] reg882 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg881 = (1'h0);
  reg [(4'hc):(1'h0)] forvar880 = (1'h0);
  reg [(3'h7):(1'h0)] reg879 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg878 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg877 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar876 = (1'h0);
  reg [(3'h4):(1'h0)] reg875 = (1'h0);
  reg [(4'hb):(1'h0)] forvar874 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg873 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar872 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg871 = (1'h0);
  reg [(5'h16):(1'h0)] reg870 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar869 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg868 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg867 = (1'h0);
  reg [(2'h3):(1'h0)] reg866 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg865 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg864 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg863 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar862 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar861 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar860 = (1'h0);
  reg [(5'h13):(1'h0)] reg859 = (1'h0);
  reg [(4'h9):(1'h0)] reg858 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar853 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg857 = (1'h0);
  reg [(5'h15):(1'h0)] reg856 = (1'h0);
  reg [(5'h12):(1'h0)] reg855 = (1'h0);
  reg signed [(4'he):(1'h0)] reg854 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg853 = (1'h0);
  reg [(4'ha):(1'h0)] reg852 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire851;
  reg [(3'h7):(1'h0)] reg850 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg849 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg848 = (1'h0);
  reg [(4'hb):(1'h0)] reg847 = (1'h0);
  wire [(4'h9):(1'h0)] wire845;
  reg signed [(4'ha):(1'h0)] reg247 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire246;
  reg [(5'h11):(1'h0)] reg240 = (1'h0);
  reg [(4'hf):(1'h0)] reg245 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg244 = (1'h0);
  reg [(5'h12):(1'h0)] reg243 = (1'h0);
  reg [(4'h8):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg241 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar240 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg239 = (1'h0);
  reg [(4'hd):(1'h0)] reg238 = (1'h0);
  reg [(4'ha):(1'h0)] reg237 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg236 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar235 = (1'h0);
  reg [(3'h7):(1'h0)] reg234 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire233;
  reg [(5'h14):(1'h0)] reg232 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg231 = (1'h0);
  reg [(3'h6):(1'h0)] forvar230 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg229 = (1'h0);
  reg [(2'h2):(1'h0)] reg228 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar227 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar226 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg225 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg224 = (1'h0);
  reg [(5'h17):(1'h0)] reg223 = (1'h0);
  reg [(5'h12):(1'h0)] reg222 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg221 = (1'h0);
  reg [(5'h13):(1'h0)] reg220 = (1'h0);
  reg [(4'hb):(1'h0)] forvar219 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg218 = (1'h0);
  reg [(5'h15):(1'h0)] forvar217 = (1'h0);
  reg [(4'hf):(1'h0)] forvar216 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg215 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar214 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg213 = (1'h0);
  reg [(5'h17):(1'h0)] reg212 = (1'h0);
  reg [(5'h13):(1'h0)] reg211 = (1'h0);
  reg [(4'ha):(1'h0)] reg210 = (1'h0);
  reg [(3'h4):(1'h0)] reg209 = (1'h0);
  reg [(4'hd):(1'h0)] forvar208 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg207 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg205 = (1'h0);
  reg [(5'h14):(1'h0)] reg204 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg203 = (1'h0);
  reg signed [(4'he):(1'h0)] reg202 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar201 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg200 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg199 = (1'h0);
  reg [(5'h13):(1'h0)] reg198 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar197 = (1'h0);
  reg [(2'h2):(1'h0)] forvar196 = (1'h0);
  reg [(5'h17):(1'h0)] reg195 = (1'h0);
  reg [(5'h15):(1'h0)] reg194 = (1'h0);
  reg [(4'hc):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar192 = (1'h0);
  reg [(5'h10):(1'h0)] reg191 = (1'h0);
  reg [(4'ha):(1'h0)] forvar190 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg189 = (1'h0);
  reg [(5'h14):(1'h0)] reg188 = (1'h0);
  reg signed [(4'he):(1'h0)] reg187 = (1'h0);
  reg [(5'h14):(1'h0)] reg186 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar185 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg184 = (1'h0);
  reg [(4'ha):(1'h0)] reg183 = (1'h0);
  assign y = {wire893,
                 reg892,
                 reg891,
                 forvar890,
                 reg889,
                 reg888,
                 reg887,
                 reg886,
                 forvar885,
                 reg884,
                 reg883,
                 reg882,
                 reg881,
                 forvar880,
                 reg879,
                 reg878,
                 reg877,
                 forvar876,
                 reg875,
                 forvar874,
                 reg873,
                 forvar872,
                 reg871,
                 reg870,
                 forvar869,
                 reg868,
                 reg867,
                 reg866,
                 reg865,
                 reg864,
                 reg863,
                 forvar862,
                 forvar861,
                 forvar860,
                 reg859,
                 reg858,
                 forvar853,
                 reg857,
                 reg856,
                 reg855,
                 reg854,
                 reg853,
                 reg852,
                 wire851,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 wire845,
                 reg247,
                 wire246,
                 reg240,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 forvar240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 forvar235,
                 reg234,
                 wire233,
                 reg232,
                 reg231,
                 forvar230,
                 reg229,
                 reg228,
                 forvar227,
                 forvar226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 forvar219,
                 reg218,
                 forvar217,
                 forvar216,
                 reg215,
                 forvar214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 forvar208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 forvar201,
                 reg200,
                 reg199,
                 reg198,
                 forvar197,
                 forvar196,
                 reg195,
                 reg194,
                 reg193,
                 forvar192,
                 reg191,
                 forvar190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 forvar185,
                 reg184,
                 reg183,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg183 <= {"z8MY8L9HIUpXau"};
      reg184 <= wire181[(3'h4):(1'h0)];
      for (forvar185 = (1'h0); (forvar185 < (1'h1)); forvar185 = (forvar185 + (1'h1)))
        begin
          reg186 <= (forvar185[(4'h8):(2'h3)] ?
              wire182[(5'h13):(4'hc)] : (&((^(|reg183)) + $unsigned("He"))));
          reg187 <= (((((wire178 == reg183) | $signed(reg183)) - forvar185[(4'hb):(4'h8)]) * wire179[(3'h5):(2'h3)]) ?
              "VAdL1Jut7Dop4xNO" : $unsigned("2HIma57vACRE"));
          reg188 <= forvar185[(3'h6):(2'h2)];
        end
      reg189 <= $unsigned(reg186);
      for (forvar190 = (1'h0); (forvar190 < (1'h1)); forvar190 = (forvar190 + (1'h1)))
        begin
          reg191 <= wire181[(3'h5):(3'h5)];
          for (forvar192 = (1'h0); (forvar192 < (2'h3)); forvar192 = (forvar192 + (1'h1)))
            begin
              reg193 = forvar185[(4'ha):(2'h3)];
              reg194 <= reg193;
              reg195 <= reg187[(3'h7):(3'h6)];
              for (forvar196 = (1'h0); (forvar196 < (2'h3)); forvar196 = (forvar196 + (1'h1)))
                begin
                  for (forvar197 = (1'h0); (forvar197 < (2'h2)); forvar197 = (forvar197 + (1'h1)))
                    begin
                      reg198 <= $unsigned({(+(~^(forvar185 ?
                              wire182 : (8'hb4))))});
                      reg199 <= (reg191[(2'h2):(2'h2)] ?
                          ((8'ha9) ?
                              forvar197 : forvar185[(4'hc):(3'h7)]) : "5IWWcUw5BFC1oDP");
                      reg200 = "B3zQ";
                    end
                  for (forvar201 = (1'h0); (forvar201 < (3'h4)); forvar201 = (forvar201 + (1'h1)))
                    begin
                      reg202 <= ((~&$signed((-$unsigned(reg195)))) ?
                          reg189 : (!$unsigned(wire180[(4'h9):(3'h4)])));
                      reg203 <= wire182[(5'h13):(3'h6)];
                      reg204 <= $unsigned($unsigned(reg187));
                      reg205 <= $signed($signed((~reg187)));
                    end
                end
              reg206 <= "";
            end
          reg207 <= (&({(+$signed(reg205)), (^forvar197[(4'ha):(1'h1)])} ?
              forvar192 : {$signed(forvar192), ""}));
          for (forvar208 = (1'h0); (forvar208 < (3'h4)); forvar208 = (forvar208 + (1'h1)))
            begin
              reg209 = ((-(!($signed(reg184) ?
                      wire180[(1'h0):(1'h0)] : $unsigned(forvar190)))) ?
                  $unsigned(((|$signed(reg199)) < ($signed((8'hb4)) ^ ((7'h40) ?
                      reg198 : forvar192)))) : wire178[(1'h1):(1'h1)]);
              reg210 <= ("EUp" ?
                  (-((reg205 + (~^(7'h42))) ?
                      {reg202[(2'h3):(2'h2)],
                          $unsigned((8'haf))} : forvar201)) : (~&reg207));
              reg211 <= $unsigned((^{forvar208[(3'h4):(2'h2)]}));
              reg212 <= {{($unsigned($signed(reg211)) ?
                          reg194[(4'ha):(4'ha)] : "CUK3P3bVKHPzrOhlK6"),
                      $unsigned((~|$unsigned(reg204)))},
                  $unsigned(("ZwfxTDqrkE" ?
                      (reg187 & $unsigned(reg195)) : (~|{reg211, reg193})))};
            end
          reg213 <= forvar201[(4'h8):(1'h1)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar214 = (1'h0); (forvar214 < (3'h4)); forvar214 = (forvar214 + (1'h1)))
        begin
          reg215 <= $unsigned(reg187);
          for (forvar216 = (1'h0); (forvar216 < (1'h1)); forvar216 = (forvar216 + (1'h1)))
            begin
              for (forvar217 = (1'h0); (forvar217 < (2'h2)); forvar217 = (forvar217 + (1'h1)))
                begin
                  reg218 <= (reg206[(3'h7):(1'h1)] ?
                      (reg205 <<< reg213) : (&(((reg203 ?
                          (8'hb5) : wire180) ^ (wire180 ?
                          reg191 : reg186)) || "UrQJVLWz")));
                  for (forvar219 = (1'h0); (forvar219 < (1'h1)); forvar219 = (forvar219 + (1'h1)))
                    begin
                      reg220 <= forvar196;
                      reg221 <= (-$unsigned($signed(((forvar192 > (8'hbd)) ?
                          (reg184 != reg186) : (!reg183)))));
                      reg222 = reg207[(3'h6):(1'h1)];
                    end
                  reg223 <= (reg204[(3'h5):(1'h1)] <<< $unsigned("S3pdh6Usdf6"));
                end
            end
          reg224 = $unsigned("JBHkrIrfg");
        end
      reg225 <= (reg191 ?
          $signed($unsigned(reg203[(1'h1):(1'h0)])) : forvar196);
      for (forvar226 = (1'h0); (forvar226 < (2'h2)); forvar226 = (forvar226 + (1'h1)))
        begin
          for (forvar227 = (1'h0); (forvar227 < (1'h1)); forvar227 = (forvar227 + (1'h1)))
            begin
              reg228 <= {$signed(((^(reg202 < forvar219)) || (~&(~|forvar226))))};
              reg229 = (8'hb2);
            end
          for (forvar230 = (1'h0); (forvar230 < (2'h2)); forvar230 = (forvar230 + (1'h1)))
            begin
              reg231 = $unsigned($unsigned((~&$unsigned($signed(forvar214)))));
            end
          reg232 <= forvar227[(3'h4):(3'h4)];
        end
    end
  assign wire233 = ((("dW7Pcr6HqQUH" ~^ ((^~(8'ha7)) ^~ forvar192)) | (~|(^"Kwn5UK2nrA"))) << "R9NZnvJdnXrJWdA9oT");
  always
    @(posedge clk) begin
      reg234 <= $signed("QrDvvmJrOL3Pp");
      for (forvar235 = (1'h0); (forvar235 < (2'h3)); forvar235 = (forvar235 + (1'h1)))
        begin
          reg236 = ({("nXgS" ?
                      $signed((reg187 ?
                          wire180 : forvar227)) : $unsigned($unsigned(reg210))),
                  (~{$signed(reg210), $signed((8'hbc))})} ?
              ((reg220[(1'h1):(1'h1)] || ((reg225 ?
                  (8'ha5) : reg189) >> reg221[(2'h3):(1'h1)])) != {forvar214}) : (8'hba));
          reg237 = {(~^reg236[(5'h12):(4'hf)]), (~|(&forvar230))};
        end
      reg238 <= forvar226;
      reg239 <= $signed($signed($unsigned(reg220)));
      if ({(-($signed((reg220 ?
              forvar230 : reg212)) <<< ("sGWdyxW" <= reg213[(4'h8):(3'h6)])))})
        begin
          for (forvar240 = (1'h0); (forvar240 < (1'h1)); forvar240 = (forvar240 + (1'h1)))
            begin
              reg241 <= "4";
              reg242 = $unsigned(reg228);
              reg243 <= reg206[(1'h1):(1'h0)];
              reg244 <= reg183;
              reg245 <= reg234;
            end
        end
      else
        begin
          reg240 <= $signed((+(!wire178)));
          reg241 <= $signed((reg243 ~^ "N9JWO6tiCBeqmVZ79LOBb"));
          reg242 <= "Ds4uREsv4TlpwDQRV06Ry";
          reg243 = $signed(reg193[(3'h4):(3'h4)]);
        end
    end
  assign wire246 = "qnp";
  always
    @(posedge clk) begin
      reg247 = reg222;
    end
  module248 modinst846 (wire845, clk, reg204, forvar227, wire181, wire182);
  always
    @(posedge clk) begin
      reg847 = ({"1g1fD2NHs9eD2f4dJfac"} + $signed($signed(forvar219[(4'h8):(4'h8)])));
      reg848 = {$signed("Nyblq8qsXwnUl01GFJ"), "VyQB8nB1G"};
      reg849 <= forvar230[(3'h4):(2'h2)];
    end
  always
    @(posedge clk) begin
      reg850 <= $signed(((^$signed($signed(forvar196))) ?
          {forvar208[(4'hb):(3'h5)]} : {(reg205[(4'hd):(4'hc)] ?
                  "YvzPECSDFd" : ((8'haf) < reg237))}));
    end
  assign wire851 = ((~|"nZHE9l7kSvGLhnn5ug") ?
                       {($signed("A") ? "V9ppAoiZ" : "TcwTTOGWy6tHwAIBd1zZ"),
                           (~&({reg238} ?
                               (reg210 ?
                                   reg228 : wire182) : $unsigned(reg202)))} : reg194);
  always
    @(posedge clk) begin
      reg852 <= $signed((wire851 ?
          reg200[(3'h6):(3'h6)] : $signed("U1Rmc6TGZ8xVRDH7")));
      if ($signed((forvar208 ?
          (($signed(forvar192) * (forvar214 >>> (8'hbc))) ?
              ($signed(reg200) ?
                  "" : "a2R6Ab6rPHS5qS") : (~^(reg207 << reg186))) : ($unsigned(reg849[(3'h4):(2'h2)]) == (reg207[(3'h7):(3'h4)] ^ (wire181 ?
              forvar196 : forvar214))))))
        begin
          reg853 = $unsigned(({forvar190[(4'ha):(3'h6)]} ^ "42rG5UNkoDKUsKvwHB"));
          reg854 <= (($signed($unsigned($unsigned(reg223))) >> $unsigned({$signed(forvar235),
                  reg195[(3'h7):(1'h1)]})) ?
              $signed($unsigned("Z9BHW1pRiacY")) : (~&reg849));
          reg855 <= ($unsigned(reg199) ?
              reg232[(5'h14):(1'h1)] : $signed((&$unsigned((^~wire851)))));
          reg856 = "tMbvvdvxEdhgc";
          reg857 <= $unsigned(wire246[(1'h0):(1'h0)]);
        end
      else
        begin
          for (forvar853 = (1'h0); (forvar853 < (1'h0)); forvar853 = (forvar853 + (1'h1)))
            begin
              reg854 = $signed(((wire180[(1'h0):(1'h0)] ^~ "yEURIbbx") ^~ ($unsigned($unsigned((8'hbc))) > $unsigned($signed(reg855)))));
              reg855 <= $unsigned(($signed((~"wB0vQ0Zu70zQ041")) && reg207));
              reg856 <= (^~forvar190[(1'h1):(1'h1)]);
              reg857 = ((+$signed((&forvar190[(1'h1):(1'h1)]))) || ($unsigned(reg212[(4'hc):(4'h8)]) || wire246));
              reg858 <= forvar219;
            end
          reg859 <= $signed(reg204[(1'h0):(1'h0)]);
          for (forvar860 = (1'h0); (forvar860 < (2'h3)); forvar860 = (forvar860 + (1'h1)))
            begin
              for (forvar861 = (1'h0); (forvar861 < (2'h2)); forvar861 = (forvar861 + (1'h1)))
                begin
                  for (forvar862 = (1'h0); (forvar862 < (1'h0)); forvar862 = (forvar862 + (1'h1)))
                    begin
                      reg863 = $signed((~^("1y00qIt47SMqMcFYlBagOp" ?
                          (reg245[(4'h9):(4'h8)] != reg199[(2'h3):(1'h1)]) : reg857[(4'hd):(4'ha)])));
                      reg864 = {$signed(reg206), (~(~&"33Tb"))};
                      reg865 = ({reg863, reg243} ?
                          {reg234,
                              ((&(forvar197 ?
                                  reg215 : reg203)) > ($unsigned(forvar190) ?
                                  (reg210 ? (8'hac) : (7'h47)) : (forvar201 ?
                                      forvar235 : (8'haa))))} : (&({"BHzo8BdlFxHB2KCQ8wHeJ1",
                                  $unsigned((7'h45))} ?
                              $signed((reg241 >>> reg852)) : reg218[(1'h0):(1'h0)])));
                    end
                end
              reg866 <= (($signed(((~|reg184) ?
                  reg200 : $unsigned(reg848))) == "p5") != reg247);
              reg867 <= ((!$unsigned(reg238[(3'h6):(1'h0)])) ?
                  reg229[(2'h2):(1'h0)] : $signed({(forvar219[(4'h8):(2'h2)] < (reg199 * reg242))}));
            end
        end
      reg868 <= wire233;
      for (forvar869 = (1'h0); (forvar869 < (1'h1)); forvar869 = (forvar869 + (1'h1)))
        begin
          reg870 <= reg215;
        end
    end
  always
    @(posedge clk) begin
      reg871 = reg205[(3'h5):(2'h3)];
    end
  always
    @(posedge clk) begin
      for (forvar872 = (1'h0); (forvar872 < (3'h4)); forvar872 = (forvar872 + (1'h1)))
        begin
          reg873 <= {({($signed(reg849) ?
                      $unsigned(forvar853) : reg204)} * "RdNhDDBw1Hu")};
        end
      for (forvar874 = (1'h0); (forvar874 < (2'h2)); forvar874 = (forvar874 + (1'h1)))
        begin
          reg875 <= (reg184 ? reg242[(1'h1):(1'h0)] : (~^(reg849 <<< "zUMi")));
          for (forvar876 = (1'h0); (forvar876 < (2'h3)); forvar876 = (forvar876 + (1'h1)))
            begin
              reg877 = reg212[(5'h17):(3'h6)];
              reg878 <= $unsigned($signed(reg228[(1'h0):(1'h0)]));
              reg879 = $signed($signed(reg877));
              for (forvar880 = (1'h0); (forvar880 < (2'h3)); forvar880 = (forvar880 + (1'h1)))
                begin
                  reg881 <= $signed(((|forvar196) ?
                      $signed(("GNVZeGH" > reg223)) : reg878));
                  reg882 = $signed("N6dbYH");
                  reg883 <= reg213;
                  reg884 = (+$unsigned("xJgD4OhOPCXmUfYMDam"));
                end
            end
        end
      for (forvar885 = (1'h0); (forvar885 < (1'h0)); forvar885 = (forvar885 + (1'h1)))
        begin
          reg886 <= $signed(reg857[(2'h2):(1'h1)]);
        end
    end
  always
    @(posedge clk) begin
      reg887 <= reg873[(3'h4):(3'h4)];
    end
  always
    @(posedge clk) begin
      reg888 <= (-forvar240);
      reg889 <= "CWqsCies7ACUR";
      for (forvar890 = (1'h0); (forvar890 < (2'h2)); forvar890 = (forvar890 + (1'h1)))
        begin
          reg891 <= {(((^~forvar217[(3'h4):(2'h3)]) | $signed((~^reg229))) ?
                  "wL3" : "ydAJXs50C3VU8JOwFI0p")};
        end
      reg892 <= {reg206[(3'h6):(3'h4)],
          $unsigned($unsigned($unsigned(reg209[(3'h4):(2'h3)])))};
    end
  assign wire893 = $unsigned(reg220[(2'h3):(1'h1)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module248
#( parameter param844 = (((((+(8'hab)) ? ((8'ha3) ? (8'hab) : (8'hb7)) : ((7'h41) ? (8'ha4) : (7'h46))) ? (8'hb3) : (((7'h43) - (8'hb8)) <<< ((8'hb9) << (8'ha3)))) ? (8'hac) : (((&(7'h46)) ? ((8'hae) ? (8'hb2) : (8'ha9)) : (8'hb4)) ? {((8'hbc) ? (7'h41) : (8'ha7))} : (^((8'hb1) <= (8'hae))))) ? ((~^(((8'h9c) ? (8'h9d) : (8'ha5)) ? (-(8'hb8)) : (~^(7'h46)))) | ({{(8'hb0)}} | (~^(&(8'h9e))))) : {((^((8'haa) ? (8'hb8) : (7'h45))) ? ({(8'hbe)} << {(8'h9e), (8'ha5)}) : (8'haf)), (((+(8'h9d)) ? ((8'ha2) >> (8'ha8)) : ((8'h9d) ? (7'h44) : (7'h47))) ? (7'h48) : (!{(8'hbb)}))}) )
(y, clk, wire252, wire251, wire250, wire249);
  output wire [(32'h321):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire252;
  input wire [(4'h8):(1'h0)] wire251;
  input wire [(5'h17):(1'h0)] wire250;
  input wire signed [(4'hb):(1'h0)] wire249;
  wire signed [(5'h17):(1'h0)] wire778;
  wire [(3'h7):(1'h0)] wire303;
  reg signed [(4'he):(1'h0)] reg302 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg301 = (1'h0);
  reg [(4'hf):(1'h0)] reg300 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg299 = (1'h0);
  reg [(3'h7):(1'h0)] reg298 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg297 = (1'h0);
  reg [(5'h16):(1'h0)] reg296 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg295 = (1'h0);
  wire [(5'h11):(1'h0)] wire294;
  reg [(4'h9):(1'h0)] reg293 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg292 = (1'h0);
  reg signed [(4'he):(1'h0)] reg291 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar290 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg289 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg288 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg287 = (1'h0);
  reg [(3'h4):(1'h0)] reg286 = (1'h0);
  reg [(4'h9):(1'h0)] reg285 = (1'h0);
  reg [(5'h10):(1'h0)] reg284 = (1'h0);
  reg [(4'hb):(1'h0)] forvar283 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg282 = (1'h0);
  reg [(5'h12):(1'h0)] reg281 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg280 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar279 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire278;
  wire signed [(4'ha):(1'h0)] wire277;
  reg signed [(3'h6):(1'h0)] reg276 = (1'h0);
  reg [(3'h7):(1'h0)] reg275 = (1'h0);
  reg [(5'h14):(1'h0)] reg274 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg273 = (1'h0);
  reg [(5'h17):(1'h0)] reg272 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg271 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar270 = (1'h0);
  reg [(5'h12):(1'h0)] reg269 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar268 = (1'h0);
  reg [(4'he):(1'h0)] reg267 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar266 = (1'h0);
  reg [(5'h17):(1'h0)] reg265 = (1'h0);
  reg [(4'h9):(1'h0)] reg264 = (1'h0);
  reg [(5'h13):(1'h0)] reg263 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg262 = (1'h0);
  wire [(4'h8):(1'h0)] wire261;
  reg [(3'h4):(1'h0)] reg260 = (1'h0);
  reg [(4'hc):(1'h0)] reg259 = (1'h0);
  reg [(4'hd):(1'h0)] reg258 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar257 = (1'h0);
  reg [(4'hd):(1'h0)] reg256 = (1'h0);
  reg [(4'ha):(1'h0)] reg255 = (1'h0);
  reg [(5'h14):(1'h0)] reg254 = (1'h0);
  reg [(4'hf):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg780 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg781 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg782 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg783 = (1'h0);
  reg [(4'h9):(1'h0)] reg784 = (1'h0);
  reg [(5'h12):(1'h0)] reg785 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg786 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg787 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg788 = (1'h0);
  reg [(5'h10):(1'h0)] reg789 = (1'h0);
  wire signed [(4'he):(1'h0)] wire842;
  assign y = {wire778,
                 wire303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 wire294,
                 reg293,
                 reg292,
                 reg291,
                 forvar290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 forvar283,
                 reg282,
                 reg281,
                 reg280,
                 forvar279,
                 wire278,
                 wire277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 forvar270,
                 reg269,
                 forvar268,
                 reg267,
                 forvar266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 wire261,
                 reg260,
                 reg259,
                 reg258,
                 forvar257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg780,
                 reg781,
                 reg782,
                 reg783,
                 reg784,
                 reg785,
                 reg786,
                 reg787,
                 reg788,
                 reg789,
                 wire842,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg253 = ((8'ha0) ?
          "DP" : ((^wire250) ? $signed($signed("OXJrYvRhVVx")) : wire250));
      reg254 <= reg253[(1'h0):(1'h0)];
      reg255 = (~^((~^(-$signed(reg254))) == (~|$unsigned(((8'ha8) >= wire252)))));
      reg256 <= (wire249 ?
          "4hffCHr1E4STEfDyz9" : ((8'h9e) ?
              (&reg254) : ($signed(wire251) > ("2xJ4ZlU3QnEH" == wire252))));
      for (forvar257 = (1'h0); (forvar257 < (1'h0)); forvar257 = (forvar257 + (1'h1)))
        begin
          reg258 <= $unsigned(("PH0V0EsogLW2Vete9J1itw" > (((reg256 - wire249) ?
                  (8'hb1) : reg255) ?
              (reg255[(1'h0):(1'h0)] ?
                  "9Mv" : ((8'hb5) || reg256)) : ({reg254} >= {reg256}))));
          reg259 = {"vU8M"};
          reg260 <= ($unsigned((((reg259 ? wire249 : (7'h45)) - {wire251,
                      wire251}) ?
                  (7'h43) : (reg254[(3'h4):(1'h0)] != "C"))) ?
              "FiLQ63pO45M1ALz" : $signed("CLgg"));
        end
    end
  assign wire261 = $unsigned(((((|reg254) ~^ $signed(reg253)) <= ($signed((7'h40)) | "0PqIqbXJmeANXx92H")) ?
                       "1JBIX3giKO" : wire250[(4'he):(4'hc)]));
  always
    @(posedge clk) begin
      if ((~&$signed(reg255)))
        begin
          reg262 <= reg255;
          reg263 = "fg3UTp4wLQ0KbK4cShy";
          reg264 <= (^~$unsigned(wire249));
          reg265 <= ($signed(wire251) << (reg256[(3'h6):(3'h4)] ?
              ((reg263[(4'he):(1'h1)] & "6pPWtGGcfrBb5yfczeo") + (^~(wire252 && reg256))) : (-((~|reg260) ?
                  (forvar257 ? (8'hb0) : reg263) : $unsigned(reg255)))));
          for (forvar266 = (1'h0); (forvar266 < (1'h1)); forvar266 = (forvar266 + (1'h1)))
            begin
              reg267 <= (!((&((wire261 ? wire252 : reg260) ?
                  (reg260 ?
                      reg254 : reg256) : wire249[(4'h8):(3'h6)])) ^~ $signed(((reg260 ?
                  forvar257 : wire252) != (~forvar266)))));
              for (forvar268 = (1'h0); (forvar268 < (1'h1)); forvar268 = (forvar268 + (1'h1)))
                begin
                  reg269 = ({wire261,
                      (+{"DdyvaGSWNasZhtA9Lm6SvO",
                          (reg258 ?
                              wire251 : wire251)})} == forvar257[(3'h6):(1'h0)]);
                  for (forvar270 = (1'h0); (forvar270 < (2'h2)); forvar270 = (forvar270 + (1'h1)))
                    begin
                      reg271 <= (8'hb5);
                      reg272 = $signed({(wire250 >= "H99Zu52Iq3RYypoJd2"),
                          {(wire251[(3'h7):(3'h7)] >>> $unsigned(reg269)),
                              ((^~reg260) > "WsID5qkBl")}});
                      reg273 <= reg263;
                    end
                end
              reg274 <= "C7gNGKn";
              reg275 = $unsigned((~^wire251[(2'h3):(2'h3)]));
              reg276 <= {forvar268[(4'hf):(2'h2)]};
            end
        end
      else
        begin
          reg262 = reg260[(1'h0):(1'h0)];
        end
    end
  assign wire277 = $unsigned($unsigned(""));
  assign wire278 = (!reg255[(2'h3):(2'h2)]);
  always
    @(posedge clk) begin
      for (forvar279 = (1'h0); (forvar279 < (2'h2)); forvar279 = (forvar279 + (1'h1)))
        begin
          reg280 <= ((({"DL82ll", reg258[(1'h1):(1'h1)]} ?
                      reg260[(3'h4):(3'h4)] : (~^{reg259})) ?
                  ($signed(((8'ha3) <= (8'ha9))) <= wire261[(3'h6):(3'h5)]) : ("KywhEF3B7" >> (|$unsigned((8'ha9))))) ?
              {$unsigned(wire277),
                  $signed(((wire249 ?
                      reg263 : (8'hbb)) < wire261))} : "odGkzqrPBI");
          reg281 <= ("8HbFh3T" ?
              {$unsigned((|reg253[(2'h2):(1'h1)]))} : reg264[(4'h9):(1'h1)]);
        end
      reg282 <= ($signed((^~$unsigned(reg271[(2'h2):(1'h0)]))) > $signed(reg267));
      for (forvar283 = (1'h0); (forvar283 < (1'h1)); forvar283 = (forvar283 + (1'h1)))
        begin
          reg284 <= reg255;
        end
      reg285 <= $signed(reg281);
      reg286 <= $signed($unsigned($signed({$signed(reg265)})));
    end
  always
    @(posedge clk) begin
      reg287 <= $signed(((&(^(reg285 != reg253))) <= (&reg269)));
      reg288 <= $unsigned((((reg260 ? (~|reg282) : (&wire250)) ?
              (^~reg263[(5'h11):(4'h9)]) : $unsigned((wire261 & reg267))) ?
          forvar266 : (forvar268 ?
              ((+reg256) ?
                  "NeyaQZaBvI" : "wJebINnl3RqBXX") : ((~|reg281) >= $signed(reg272)))));
      reg289 <= ($unsigned(forvar279) ?
          $signed({$unsigned(wire277)}) : (+forvar257));
      for (forvar290 = (1'h0); (forvar290 < (3'h4)); forvar290 = (forvar290 + (1'h1)))
        begin
          reg291 = {"EHhRQECeHMqH099k", "CO2xGJy4"};
          reg292 = $unsigned($signed(("czcpO1sNGlB3tH7kUspvk" ?
              forvar257[(4'h8):(2'h2)] : (+wire261[(1'h1):(1'h1)]))));
          reg293 <= ((~^(|"NDZOaRMwg")) <= forvar290);
        end
    end
  assign wire294 = (&("MwH" || $signed(wire261)));
  always
    @(posedge clk) begin
      reg295 <= $unsigned(wire250[(4'hd):(4'ha)]);
      reg296 <= $signed(((+(~&$unsigned(reg288))) & forvar283));
      reg297 <= ("Wc97f3K19Ez" < (reg265[(3'h7):(3'h7)] && reg291[(1'h0):(1'h0)]));
      reg298 <= (!(&$unsigned(reg262[(3'h4):(1'h1)])));
    end
  always
    @(posedge clk) begin
      reg299 <= reg296[(1'h0):(1'h0)];
      reg300 <= "SiT3m1XJO1NAWKvu7onA";
      reg301 <= reg258[(4'hb):(3'h4)];
      reg302 = forvar283;
    end
  assign wire303 = wire252[(3'h6):(3'h5)];
  module304 modinst779 (.y(wire778), .clk(clk), .wire306(reg265), .wire307(reg259), .wire308(reg253), .wire305(reg286), .wire309(reg272));
  always
    @(posedge clk) begin
      reg780 <= forvar257[(1'h0):(1'h0)];
      reg781 <= forvar270[(4'ha):(2'h2)];
      reg782 = (~&$unsigned($unsigned(reg281[(4'hf):(4'h8)])));
    end
  always
    @(posedge clk) begin
      reg783 <= $unsigned({"k63", reg253});
      reg784 <= "clSXP77Ifa6VFCO88t0qK3";
    end
  always
    @(posedge clk) begin
      reg785 = $signed($signed($unsigned({$unsigned(reg302), forvar279})));
      reg786 <= $unsigned((~&($signed({reg295,
          wire261}) || ({(8'h9e)} >> $signed(reg275)))));
      reg787 <= {(wire278[(2'h2):(2'h2)] ?
              $signed((reg260[(1'h0):(1'h0)] ?
                  (reg299 & reg255) : (reg260 ?
                      reg782 : wire251))) : (~reg785))};
    end
  always
    @(posedge clk) begin
      reg788 <= $signed(((~&("EG5JAJz6HSd7eOv0" & reg260)) ?
          ($unsigned(((8'ha8) ?
              reg291 : reg267)) < $unsigned($unsigned(reg272))) : ((~"FXFNbo9gyJitacpyu") ?
              "DBbL4L2X3ShHlRYUV" : reg296)));
    end
  always
    @(posedge clk) begin
      reg789 <= reg787[(4'h9):(4'h9)];
    end
  module790 modinst843 (wire842, clk, reg263, reg787, reg272, wire778, reg265);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module790
#( parameter param841 = ({(^(((8'hae) ? (8'ha3) : (8'hb1)) + ((8'hbd) ? (8'hac) : (7'h44)))), (8'hb1)} ? (((((8'h9f) ? (8'h9f) : (8'haf)) * {(7'h46)}) == (((7'h48) | (8'hbd)) ? (!(8'h9e)) : {(8'ha4)})) ? ((7'h40) ? (~^((8'h9f) == (8'ha1))) : ((!(8'hb6)) - ((8'haf) <= (8'hb7)))) : ((!((8'hae) <= (8'hae))) + (&{(8'hbd)}))) : (7'h42)) )
(y, clk, wire795, wire794, wire793, wire792, wire791);
  output wire [(32'h1fd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire795;
  input wire signed [(3'h6):(1'h0)] wire794;
  input wire signed [(5'h17):(1'h0)] wire793;
  input wire signed [(5'h17):(1'h0)] wire792;
  input wire signed [(5'h17):(1'h0)] wire791;
  reg signed [(3'h6):(1'h0)] reg840 = (1'h0);
  reg [(3'h4):(1'h0)] forvar839 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg838 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg837 = (1'h0);
  reg [(5'h17):(1'h0)] reg836 = (1'h0);
  reg [(4'hb):(1'h0)] reg835 = (1'h0);
  reg [(3'h4):(1'h0)] reg834 = (1'h0);
  reg [(4'hb):(1'h0)] forvar833 = (1'h0);
  reg [(5'h14):(1'h0)] reg832 = (1'h0);
  reg [(5'h15):(1'h0)] reg831 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg830 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg829 = (1'h0);
  reg [(5'h12):(1'h0)] reg828 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg827 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg826 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg825 = (1'h0);
  reg [(5'h14):(1'h0)] reg824 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar823 = (1'h0);
  reg [(3'h4):(1'h0)] reg822 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg821 = (1'h0);
  reg [(5'h11):(1'h0)] reg820 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg819 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar818 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg817 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg816 = (1'h0);
  reg [(3'h6):(1'h0)] reg815 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg814 = (1'h0);
  reg [(4'hc):(1'h0)] reg813 = (1'h0);
  reg [(4'h9):(1'h0)] reg812 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire811;
  reg signed [(5'h11):(1'h0)] reg810 = (1'h0);
  reg [(4'h9):(1'h0)] reg809 = (1'h0);
  reg [(3'h5):(1'h0)] reg808 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire807;
  reg [(4'ha):(1'h0)] reg806 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg805 = (1'h0);
  reg [(2'h3):(1'h0)] reg804 = (1'h0);
  reg [(4'hb):(1'h0)] reg803 = (1'h0);
  reg [(2'h2):(1'h0)] reg802 = (1'h0);
  reg [(3'h5):(1'h0)] reg801 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire800;
  reg signed [(4'he):(1'h0)] reg799 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg798 = (1'h0);
  reg [(2'h2):(1'h0)] reg797 = (1'h0);
  wire [(3'h5):(1'h0)] wire796;
  assign y = {reg840,
                 forvar839,
                 reg838,
                 reg837,
                 reg836,
                 reg835,
                 reg834,
                 forvar833,
                 reg832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 reg827,
                 reg826,
                 reg825,
                 reg824,
                 forvar823,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 forvar818,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 reg812,
                 wire811,
                 reg810,
                 reg809,
                 reg808,
                 wire807,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg802,
                 reg801,
                 wire800,
                 reg799,
                 reg798,
                 reg797,
                 wire796,
                 (1'h0)};
  assign wire796 = (+"UNx9FL0AHchOU");
  always
    @(posedge clk) begin
      reg797 = "2Yl7iINZLl5D";
      reg798 = reg797[(2'h2):(1'h0)];
      reg799 <= $unsigned($signed({"zqxR41zE8"}));
    end
  assign wire800 = $unsigned("71TP8iCoEyzf");
  always
    @(posedge clk) begin
      reg801 <= ((+wire796[(3'h4):(1'h0)]) ~^ (^~"5a18KabE7sgbUkI0Hf"));
      reg802 = wire796[(3'h5):(3'h5)];
      reg803 <= (~&(+wire800));
    end
  always
    @(posedge clk) begin
      reg804 = wire795[(4'h8):(4'h8)];
      reg805 = "EiNzcH5pN2THpC4h94";
      reg806 = $signed(reg804[(1'h1):(1'h1)]);
    end
  assign wire807 = $signed(((+(^~{reg798})) & (~^((reg799 << wire796) ?
                       {(7'h45)} : (wire795 ? reg803 : reg802)))));
  always
    @(posedge clk) begin
      reg808 <= "CesoNYam7Wxot";
      reg809 = ((reg803 >> (({(8'hb0), wire793} < reg804[(1'h1):(1'h1)]) ?
              wire807[(4'ha):(3'h7)] : "A9RAOXBYbUKO7dGip0Ic")) ?
          ((~(-$unsigned(wire791))) ^ {"oMRLEsZWap",
              reg803}) : {$signed(wire793[(4'ha):(4'h9)]),
              "9Q1eCdvipJUuyyfLM155o"});
      reg810 <= $signed("yoPBOZOTrVcFRe");
    end
  assign wire811 = $signed(wire795);
  always
    @(posedge clk) begin
      reg812 <= {$signed((wire795[(5'h11):(3'h7)] ?
              $unsigned(reg799[(1'h1):(1'h0)]) : $unsigned($unsigned(wire793)))),
          reg798[(3'h7):(3'h4)]};
      reg813 <= "eW3B7M";
      reg814 <= ((reg812[(3'h4):(2'h2)] ?
              (wire793 ?
                  $unsigned((reg812 << (8'hac))) : $unsigned(reg798)) : $unsigned(reg809[(3'h5):(3'h5)])) ?
          ($unsigned("eIlQHAEZdhxWi") ?
              (7'h40) : (!{(reg797 - reg802),
                  (reg803 ?
                      wire807 : wire792)})) : $signed(($signed($unsigned(reg806)) ?
              {"", (8'hb0)} : ((wire791 ~^ reg809) ?
                  reg810[(1'h0):(1'h0)] : (reg809 > reg809)))));
    end
  always
    @(posedge clk) begin
      reg815 <= reg809;
    end
  always
    @(posedge clk) begin
      reg816 <= (~|wire795[(5'h10):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg817 = $unsigned(reg815);
    end
  always
    @(posedge clk) begin
      for (forvar818 = (1'h0); (forvar818 < (2'h2)); forvar818 = (forvar818 + (1'h1)))
        begin
          reg819 <= $signed({(~$unsigned((wire792 ? reg799 : wire811))),
              reg808});
          reg820 <= $signed($unsigned("iW"));
          reg821 <= (({$unsigned($unsigned(reg799))} < ({$unsigned(wire792),
                  "hWu2zqfYtZf3YMpns"} ?
              "AtT" : $unsigned((wire792 ^ wire795)))) >> "h7dZbny");
          reg822 <= wire811[(1'h1):(1'h1)];
        end
      for (forvar823 = (1'h0); (forvar823 < (2'h2)); forvar823 = (forvar823 + (1'h1)))
        begin
          if ($signed((~reg802)))
            begin
              reg824 = reg797[(1'h0):(1'h0)];
              reg825 <= $signed($signed(($unsigned((&reg808)) == reg808)));
              reg826 <= $unsigned((^~(wire792[(4'hc):(3'h4)] >> $signed($unsigned(wire792)))));
              reg827 = wire807[(4'h9):(2'h2)];
              reg828 = (-reg799);
            end
          else
            begin
              reg824 = "dA1mXlOPhMIKLs";
              reg825 <= $unsigned("X8PoUdl");
            end
          reg829 <= {"cZJNW2gOflwmvqFNI4HJL",
              $unsigned($unsigned(("IFhL4lQ" ?
                  $signed(reg820) : reg828[(3'h4):(1'h0)])))};
          reg830 <= "GHikWkm5aAhD";
          reg831 <= (reg825 ? $unsigned("O") : $signed((!reg809)));
          reg832 <= (+(~&(~reg804)));
        end
      for (forvar833 = (1'h0); (forvar833 < (3'h4)); forvar833 = (forvar833 + (1'h1)))
        begin
          reg834 <= $signed($unsigned({(^~reg819)}));
          reg835 <= (~reg801[(2'h2):(1'h1)]);
          reg836 = (+$signed($unsigned((^wire811[(3'h4):(2'h3)]))));
          reg837 <= ({(^($signed(reg825) <= (wire791 < (8'hbd))))} ?
              (!$signed(reg813[(4'h9):(3'h6)])) : "s");
          reg838 = ($unsigned(reg831) <= $unsigned({(8'hb9)}));
        end
      for (forvar839 = (1'h0); (forvar839 < (1'h1)); forvar839 = (forvar839 + (1'h1)))
        begin
          reg840 = $unsigned(reg820);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module304
#( parameter param776 = ((-((((8'haf) ? (8'hbf) : (8'ha7)) ? (~^(7'h47)) : {(8'ha3)}) == (((8'hbb) + (7'h43)) & (~(7'h44))))) == {(((-(8'ha2)) < (|(7'h45))) ^ (^((7'h41) ? (8'ha5) : (8'h9d)))), ((^(~(7'h40))) ? (&((8'hb1) ? (8'hb6) : (8'ha6))) : (|((8'hb5) ? (8'hb3) : (8'ha3))))})
, parameter param777 = {(({((8'hac) ^ (8'hbd))} * param776) != {(8'hbf), (|param776)}), (!(8'hb5))} )
(y, clk, wire305, wire306, wire307, wire308, wire309);
  output wire [(32'h56a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire305;
  input wire [(4'hb):(1'h0)] wire306;
  input wire signed [(4'h8):(1'h0)] wire307;
  input wire [(4'hf):(1'h0)] wire308;
  input wire signed [(2'h2):(1'h0)] wire309;
  reg [(5'h15):(1'h0)] reg775 = (1'h0);
  reg [(2'h3):(1'h0)] reg774 = (1'h0);
  reg signed [(4'he):(1'h0)] reg773 = (1'h0);
  reg [(4'hf):(1'h0)] reg772 = (1'h0);
  reg [(5'h11):(1'h0)] reg771 = (1'h0);
  reg [(4'he):(1'h0)] forvar770 = (1'h0);
  reg [(4'hc):(1'h0)] forvar769 = (1'h0);
  reg [(4'ha):(1'h0)] reg768 = (1'h0);
  reg [(5'h10):(1'h0)] reg767 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg766 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg765 = (1'h0);
  reg [(3'h6):(1'h0)] forvar764 = (1'h0);
  reg [(4'h9):(1'h0)] reg763 = (1'h0);
  reg [(3'h7):(1'h0)] reg762 = (1'h0);
  reg [(2'h2):(1'h0)] reg761 = (1'h0);
  reg [(5'h12):(1'h0)] forvar760 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg759 = (1'h0);
  reg [(3'h5):(1'h0)] reg758 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg757 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg756 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar755 = (1'h0);
  reg [(5'h15):(1'h0)] forvar754 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg753 = (1'h0);
  reg [(4'ha):(1'h0)] reg752 = (1'h0);
  reg [(5'h11):(1'h0)] reg751 = (1'h0);
  reg [(2'h3):(1'h0)] forvar310 = (1'h0);
  reg [(4'h9):(1'h0)] reg311 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg312 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg313 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar315 = (1'h0);
  reg [(4'h9):(1'h0)] reg316 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg317 = (1'h0);
  reg [(4'hd):(1'h0)] reg318 = (1'h0);
  wire [(3'h4):(1'h0)] wire319;
  wire [(5'h11):(1'h0)] wire320;
  reg signed [(3'h6):(1'h0)] reg321 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar322 = (1'h0);
  reg [(5'h14):(1'h0)] forvar323 = (1'h0);
  reg [(5'h10):(1'h0)] forvar324 = (1'h0);
  reg [(4'he):(1'h0)] reg325 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar326 = (1'h0);
  reg [(5'h13):(1'h0)] reg327 = (1'h0);
  reg [(4'he):(1'h0)] reg328 = (1'h0);
  reg [(4'h8):(1'h0)] reg329 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg330 = (1'h0);
  reg signed [(4'he):(1'h0)] reg331 = (1'h0);
  reg [(5'h15):(1'h0)] forvar332 = (1'h0);
  reg [(4'ha):(1'h0)] reg333 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg334 = (1'h0);
  reg [(3'h7):(1'h0)] reg335 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg336 = (1'h0);
  reg [(5'h14):(1'h0)] reg337 = (1'h0);
  reg [(3'h7):(1'h0)] reg338 = (1'h0);
  reg [(5'h15):(1'h0)] reg339 = (1'h0);
  reg [(4'hf):(1'h0)] reg340 = (1'h0);
  reg [(4'hf):(1'h0)] reg341 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar342 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg344 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg345 = (1'h0);
  reg [(3'h4):(1'h0)] reg346 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg347 = (1'h0);
  reg [(5'h11):(1'h0)] reg348 = (1'h0);
  reg [(3'h5):(1'h0)] reg349 = (1'h0);
  reg [(5'h11):(1'h0)] reg350 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg351 = (1'h0);
  wire [(3'h6):(1'h0)] wire352;
  reg signed [(4'ha):(1'h0)] reg353 = (1'h0);
  reg [(5'h14):(1'h0)] reg354 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg355 = (1'h0);
  reg [(5'h15):(1'h0)] reg356 = (1'h0);
  reg [(4'h8):(1'h0)] reg357 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg358 = (1'h0);
  reg [(4'h9):(1'h0)] reg359 = (1'h0);
  reg [(3'h5):(1'h0)] reg360 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar361 = (1'h0);
  reg [(3'h6):(1'h0)] reg362 = (1'h0);
  reg [(5'h12):(1'h0)] reg363 = (1'h0);
  reg [(5'h17):(1'h0)] forvar364 = (1'h0);
  reg [(5'h16):(1'h0)] reg365 = (1'h0);
  reg [(5'h13):(1'h0)] reg366 = (1'h0);
  reg [(4'hf):(1'h0)] forvar367 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg368 = (1'h0);
  reg [(2'h2):(1'h0)] reg369 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar370 = (1'h0);
  reg [(4'he):(1'h0)] reg371 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg372 = (1'h0);
  reg [(4'hb):(1'h0)] reg373 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg374 = (1'h0);
  reg [(4'hc):(1'h0)] reg375 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg376 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar377 = (1'h0);
  reg signed [(4'he):(1'h0)] reg378 = (1'h0);
  reg [(5'h17):(1'h0)] reg379 = (1'h0);
  reg [(5'h12):(1'h0)] forvar380 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg381 = (1'h0);
  reg [(3'h4):(1'h0)] reg382 = (1'h0);
  reg [(5'h15):(1'h0)] reg383 = (1'h0);
  reg [(5'h12):(1'h0)] reg384 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg385 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg386 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire387;
  wire [(3'h5):(1'h0)] wire388;
  reg [(5'h12):(1'h0)] reg389 = (1'h0);
  reg [(4'h8):(1'h0)] reg390 = (1'h0);
  reg [(4'hb):(1'h0)] reg391 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg392 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg393 = (1'h0);
  reg [(4'hd):(1'h0)] reg394 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire749;
  assign y = {reg775,
                 reg774,
                 reg773,
                 reg772,
                 reg771,
                 forvar770,
                 forvar769,
                 reg768,
                 reg767,
                 reg766,
                 reg765,
                 forvar764,
                 reg763,
                 reg762,
                 reg761,
                 forvar760,
                 reg759,
                 reg758,
                 reg757,
                 reg756,
                 forvar755,
                 forvar754,
                 reg753,
                 reg752,
                 reg751,
                 forvar310,
                 reg311,
                 reg312,
                 reg313,
                 reg314,
                 forvar315,
                 reg316,
                 reg317,
                 reg318,
                 wire319,
                 wire320,
                 reg321,
                 forvar322,
                 forvar323,
                 forvar324,
                 reg325,
                 forvar326,
                 reg327,
                 reg328,
                 reg329,
                 reg330,
                 reg331,
                 forvar332,
                 reg333,
                 reg334,
                 reg335,
                 reg336,
                 reg337,
                 reg338,
                 reg339,
                 reg340,
                 reg341,
                 forvar342,
                 reg343,
                 reg344,
                 reg345,
                 reg346,
                 reg347,
                 reg348,
                 reg349,
                 reg350,
                 reg351,
                 wire352,
                 reg353,
                 reg354,
                 reg355,
                 reg356,
                 reg357,
                 reg358,
                 reg359,
                 reg360,
                 forvar361,
                 reg362,
                 reg363,
                 forvar364,
                 reg365,
                 reg366,
                 forvar367,
                 reg368,
                 reg369,
                 forvar370,
                 reg371,
                 reg372,
                 reg373,
                 reg374,
                 reg375,
                 reg376,
                 forvar377,
                 reg378,
                 reg379,
                 forvar380,
                 reg381,
                 reg382,
                 reg383,
                 reg384,
                 reg385,
                 reg386,
                 wire387,
                 wire388,
                 reg389,
                 reg390,
                 reg391,
                 reg392,
                 reg393,
                 reg394,
                 wire749,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar310 = (1'h0); (forvar310 < (1'h0)); forvar310 = (forvar310 + (1'h1)))
        begin
          reg311 <= (wire309[(2'h2):(2'h2)] <<< $unsigned($signed($unsigned((wire308 <= (8'hba))))));
          reg312 <= wire305[(2'h2):(1'h1)];
        end
      reg313 <= $signed((7'h47));
      reg314 <= $signed($unsigned("etmBp5"));
      for (forvar315 = (1'h0); (forvar315 < (3'h4)); forvar315 = (forvar315 + (1'h1)))
        begin
          reg316 = wire309[(1'h1):(1'h1)];
          reg317 <= {{wire306},
              $unsigned(((~^$signed(wire309)) ?
                  $signed((reg312 & reg311)) : "va"))};
          reg318 = $signed($unsigned($signed($signed((wire305 >> forvar315)))));
        end
    end
  assign wire319 = $unsigned((($unsigned((wire308 & wire305)) ?
                           $unsigned({reg316, reg314}) : "13RXa") ?
                       reg311[(4'h9):(4'h8)] : (reg312 ?
                           $unsigned({reg312}) : "NJezLQV9MENmsX9i")));
  assign wire320 = $unsigned(($unsigned({{wire309},
                       $signed(wire319)}) && forvar315));
  always
    @(posedge clk) begin
      reg321 <= (|$signed((&$signed($signed(wire308)))));
      for (forvar322 = (1'h0); (forvar322 < (3'h4)); forvar322 = (forvar322 + (1'h1)))
        begin
          for (forvar323 = (1'h0); (forvar323 < (2'h3)); forvar323 = (forvar323 + (1'h1)))
            begin
              for (forvar324 = (1'h0); (forvar324 < (1'h1)); forvar324 = (forvar324 + (1'h1)))
                begin
                  reg325 = "AX";
                  for (forvar326 = (1'h0); (forvar326 < (2'h2)); forvar326 = (forvar326 + (1'h1)))
                    begin
                      reg327 <= ((!$signed(("2OSzf1hPD7BVtf" & ((8'ha1) * (8'hb7))))) ^ "efoWYyu19g");
                      reg328 <= "DSX70hptYBu0herWf";
                      reg329 = ("EXQmgF2TwFici5XbD" ~^ reg313);
                    end
                  reg330 <= $signed("KZMUF5G1s");
                end
              reg331 <= ({(|$unsigned("adePoYfG1O")), "SLcAoUKN4mK"} ?
                  wire309[(1'h1):(1'h1)] : {reg311});
              for (forvar332 = (1'h0); (forvar332 < (1'h0)); forvar332 = (forvar332 + (1'h1)))
                begin
                  reg333 <= (~|(^(+$unsigned({wire320}))));
                  reg334 <= (reg327[(2'h3):(2'h3)] ^~ ($unsigned("yD") <<< $unsigned({$unsigned(reg328),
                      $unsigned(forvar326)})));
                  reg335 = reg317[(3'h5):(2'h2)];
                  reg336 <= "bhYGNKDfYWhwBzNI3";
                end
              reg337 = $signed((&"bPxV"));
            end
          reg338 <= "s9chx7";
        end
      reg339 <= (reg314[(4'hc):(2'h2)] ?
          $signed((-reg338)) : ("qn4FfZz8vxRAVByE3qJ0IL" >= (^$signed((8'ha5)))));
      reg340 = $unsigned({"Abdqsaz8UwOnELDLpAwEwi"});
    end
  always
    @(posedge clk) begin
      reg341 <= $unsigned((~&(-reg316[(2'h2):(2'h2)])));
    end
  always
    @(posedge clk) begin
      for (forvar342 = (1'h0); (forvar342 < (2'h3)); forvar342 = (forvar342 + (1'h1)))
        begin
          reg343 = $unsigned($signed((-(7'h43))));
        end
      reg344 <= "CVy1leY";
      reg345 <= $unsigned("");
      reg346 <= reg318[(2'h3):(1'h1)];
      reg347 = (reg334 ? (-reg339[(4'ha):(3'h6)]) : reg312);
    end
  always
    @(posedge clk) begin
      reg348 <= ($signed((&(8'haa))) ?
          ($signed((^~((8'hbc) ?
              reg317 : reg344))) == {forvar324[(1'h1):(1'h1)],
              ($signed(wire309) ? reg346 : (^reg331))}) : {(8'hb4)});
      reg349 <= $signed($signed($signed($signed("vruX39FArDPugWYgOAcJLh"))));
      reg350 <= reg318[(3'h5):(2'h3)];
      reg351 <= (((wire320[(4'he):(4'ha)] * ((reg348 ? reg336 : (8'ha5)) ?
              $signed(forvar332) : (~reg350))) ?
          ((|(&reg334)) ?
              $unsigned("hiK2n") : ((reg336 ? wire307 : wire320) ?
                  reg328 : (^~reg318))) : reg316) ^ reg347[(2'h3):(2'h3)]);
    end
  assign wire352 = "lCSrYzffLMWh9P0K";
  always
    @(posedge clk) begin
      reg353 <= {$unsigned("CUIRUIfiScW7"),
          (-((+"pP") ? reg335[(2'h2):(2'h2)] : wire319[(1'h1):(1'h0)]))};
      reg354 <= reg339;
      reg355 = (($signed((^~(~^reg325))) ?
              (^((reg314 <<< (8'h9e)) != $unsigned(reg354))) : forvar315) ?
          ($unsigned(reg350) ?
              ({forvar323} != ((^~reg314) ?
                  reg329[(2'h2):(1'h0)] : wire320[(3'h6):(2'h2)])) : $unsigned(((wire307 < reg312) ?
                  forvar315 : ((8'ha0) == reg331)))) : (~^forvar315[(4'he):(2'h3)]));
      reg356 <= ($unsigned((wire305 > reg337[(4'h8):(2'h2)])) ~^ reg337[(5'h13):(3'h5)]);
    end
  always
    @(posedge clk) begin
      reg357 <= "XQNhAYh";
      reg358 = reg316;
      reg359 <= (-((^~"THrBX7UD") ?
          $unsigned(($unsigned(reg338) < $unsigned(reg343))) : wire319));
      reg360 <= $signed(reg330[(4'ha):(3'h4)]);
    end
  always
    @(posedge clk) begin
      for (forvar361 = (1'h0); (forvar361 < (2'h3)); forvar361 = (forvar361 + (1'h1)))
        begin
          reg362 <= (-($unsigned((!$signed(reg328))) ?
              reg338[(1'h1):(1'h1)] : ((forvar332 - "PC") ?
                  (-$unsigned((8'hbd))) : wire352)));
        end
      reg363 <= (~$unsigned($unsigned(((forvar326 >>> reg312) || $unsigned(wire319)))));
      for (forvar364 = (1'h0); (forvar364 < (1'h0)); forvar364 = (forvar364 + (1'h1)))
        begin
          reg365 = "3BLzrzhX";
          reg366 <= (((reg335 ?
              reg340[(1'h0):(1'h0)] : (wire307[(1'h0):(1'h0)] ?
                  reg330 : $signed(reg328))) <= reg363) < (forvar324[(3'h5):(1'h1)] ?
              (~(wire306 ?
                  "5" : {forvar342,
                      wire320})) : {$unsigned("TnM26Qntn7VM2KI1K4biHu")}));
          for (forvar367 = (1'h0); (forvar367 < (2'h2)); forvar367 = (forvar367 + (1'h1)))
            begin
              reg368 = forvar324[(2'h3):(2'h2)];
              reg369 <= reg330[(3'h6):(2'h2)];
              for (forvar370 = (1'h0); (forvar370 < (1'h1)); forvar370 = (forvar370 + (1'h1)))
                begin
                  reg371 <= ((($signed($unsigned(reg333)) ~^ {forvar364[(3'h6):(3'h4)],
                              (~|wire307)}) ?
                          (forvar324 ?
                              $unsigned($unsigned(reg360)) : ((~forvar322) ?
                                  (8'h9c) : "EpZgx6xPIanBNv2G")) : $unsigned(forvar367[(2'h2):(1'h0)])) ?
                      $signed($unsigned($unsigned(reg327))) : "vQU8cR");
                  reg372 = $unsigned((!$unsigned("R7z6w3XGybnJBEKaocbA")));
                  reg373 <= $signed(forvar310[(1'h1):(1'h0)]);
                  reg374 <= (forvar364 ?
                      (|"9fxechCueszt") : (-$signed(reg359)));
                end
              reg375 <= {{{"tfedQKfqKztdRWP", forvar332[(3'h7):(3'h5)]},
                      {reg327}}};
              reg376 <= $unsigned("VJVxO0gp9IBgJdKiJiN");
            end
        end
      for (forvar377 = (1'h0); (forvar377 < (1'h1)); forvar377 = (forvar377 + (1'h1)))
        begin
          reg378 <= "2QooxoWGOvVOdu";
          reg379 <= {$unsigned(reg321[(2'h2):(1'h1)]),
              $unsigned(wire319[(2'h2):(2'h2)])};
          for (forvar380 = (1'h0); (forvar380 < (2'h3)); forvar380 = (forvar380 + (1'h1)))
            begin
              reg381 = {(~reg371[(3'h7):(3'h7)]),
                  ((("rxvrp" & reg351[(2'h3):(1'h0)]) & $unsigned((~wire307))) ?
                      (^($signed(reg318) == reg337)) : ({$unsigned(reg333)} | {reg351}))};
              reg382 = ("iUT" ? reg318[(3'h5):(1'h1)] : "4xdLs002PrkMu1tUc");
              reg383 = (|"d");
              reg384 = forvar332[(4'hc):(2'h2)];
            end
          reg385 = "y";
        end
      reg386 <= $unsigned(((&$unsigned((7'h42))) >> forvar332));
    end
  assign wire387 = ($signed($unsigned($unsigned((&(8'haf))))) ?
                       "dp1" : ({(-"9eem791axd29eF74a")} ?
                           {$unsigned({(8'haa), (8'hb6)}), reg379} : reg376));
  assign wire388 = forvar361;
  always
    @(posedge clk) begin
      reg389 <= $unsigned(((8'ha9) ? "cH" : $unsigned("3doRB")));
    end
  always
    @(posedge clk) begin
      reg390 <= ((!"EVJ29eSMQ") ?
          $unsigned($unsigned($signed(forvar370))) : "e4iKl2QIq3176aS1");
      reg391 = ($signed((~|($signed(reg354) ?
              {reg353, (7'h44)} : $signed((8'hb9))))) ?
          $signed($signed((reg329[(2'h2):(1'h1)] ?
              (reg344 << reg346) : reg316[(1'h1):(1'h0)]))) : "V3qQapE5");
      reg392 = (("m1LPYcmkYXmKJFmaKahNZ" && {reg328[(4'h8):(3'h4)],
              ((reg312 ? reg311 : wire320) == reg339[(4'hc):(4'h9)])}) ?
          $unsigned((~forvar315)) : (reg363 < $unsigned(forvar332[(2'h3):(2'h2)])));
      reg393 <= $signed($unsigned(reg389[(1'h0):(1'h0)]));
      reg394 = ($signed(reg311[(4'h8):(3'h7)]) ?
          $signed("rDbothGu0knMR2p3GcV90y") : $signed($signed($signed((forvar377 ?
              wire307 : reg325)))));
    end
  module395 modinst750 (wire749, clk, reg385, reg331, reg313, reg356, forvar324);
  always
    @(posedge clk) begin
      reg751 <= $unsigned({(^~{(reg389 ? reg350 : reg393),
              (reg384 >>> reg312)})});
      reg752 <= $signed((("fpAUckqo5vqZD" + $unsigned((|reg353))) & (+reg393)));
      reg753 = (8'ha6);
      for (forvar754 = (1'h0); (forvar754 < (1'h0)); forvar754 = (forvar754 + (1'h1)))
        begin
          for (forvar755 = (1'h0); (forvar755 < (3'h4)); forvar755 = (forvar755 + (1'h1)))
            begin
              reg756 <= (^~$signed(reg329));
              reg757 <= ({(~&$unsigned((reg351 ? reg321 : forvar754))),
                      $unsigned(reg389)} ?
                  $unsigned($signed(($signed(reg331) + reg337))) : ($signed(((wire309 ^ reg386) <= (reg355 ?
                      wire309 : (8'hb6)))) != (~^("Q6b" ?
                      (+reg360) : $unsigned(reg366)))));
              reg758 <= (((8'h9c) ~^ "2xPMGp3u0") ?
                  (7'h45) : reg384[(4'hd):(2'h3)]);
              reg759 = (|reg393[(3'h4):(2'h3)]);
            end
          for (forvar760 = (1'h0); (forvar760 < (2'h2)); forvar760 = (forvar760 + (1'h1)))
            begin
              reg761 = "H7d";
              reg762 <= $unsigned("rW6QtSagFh");
              reg763 <= wire749;
              for (forvar764 = (1'h0); (forvar764 < (3'h4)); forvar764 = (forvar764 + (1'h1)))
                begin
                  reg765 <= (!forvar764);
                  reg766 <= ((~&reg761[(2'h2):(1'h1)]) ^ $unsigned(reg375[(2'h3):(2'h2)]));
                  reg767 <= forvar764;
                  reg768 = $unsigned((&(reg313[(3'h5):(2'h2)] <<< $signed($signed(forvar377)))));
                end
            end
        end
      for (forvar769 = (1'h0); (forvar769 < (1'h0)); forvar769 = (forvar769 + (1'h1)))
        begin
          for (forvar770 = (1'h0); (forvar770 < (3'h4)); forvar770 = (forvar770 + (1'h1)))
            begin
              reg771 <= $signed($unsigned($signed((reg354 & wire306))));
              reg772 <= reg759[(2'h2):(1'h0)];
            end
          reg773 = (forvar367 - ((((|(8'hae)) ?
              (reg354 > wire352) : (reg366 >= reg757)) < $signed({forvar361})) & $unsigned(($unsigned(reg316) ?
              "0IW" : forvar342))));
          reg774 <= $unsigned($signed($unsigned(($unsigned((8'hb4)) | (reg758 | reg390)))));
          reg775 = {reg340};
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module395  (y, clk, wire396, wire397, wire398, wire399, wire400);
  output wire [(32'h3cc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire396;
  input wire signed [(4'he):(1'h0)] wire397;
  input wire [(3'h5):(1'h0)] wire398;
  input wire [(5'h15):(1'h0)] wire399;
  input wire signed [(5'h10):(1'h0)] wire400;
  reg signed [(2'h3):(1'h0)] reg748 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg747 = (1'h0);
  reg [(3'h4):(1'h0)] reg746 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg745 = (1'h0);
  reg [(3'h5):(1'h0)] reg744 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg743 = (1'h0);
  reg signed [(4'he):(1'h0)] reg742 = (1'h0);
  reg [(2'h2):(1'h0)] reg741 = (1'h0);
  reg [(4'hf):(1'h0)] reg740 = (1'h0);
  reg [(3'h5):(1'h0)] reg739 = (1'h0);
  reg [(2'h3):(1'h0)] reg738 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg737 = (1'h0);
  reg [(4'he):(1'h0)] reg736 = (1'h0);
  reg [(3'h5):(1'h0)] reg735 = (1'h0);
  reg [(4'hd):(1'h0)] forvar734 = (1'h0);
  reg [(5'h15):(1'h0)] forvar733 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire732;
  reg signed [(4'hf):(1'h0)] reg731 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg730 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg401 = (1'h0);
  reg [(5'h14):(1'h0)] reg402 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar403 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg404 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg405 = (1'h0);
  reg [(5'h11):(1'h0)] reg406 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg407 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg408 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar409 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg410 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg411 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg412 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg413 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg414 = (1'h0);
  reg [(4'he):(1'h0)] forvar415 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg417 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg418 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg419 = (1'h0);
  reg [(5'h12):(1'h0)] reg420 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg421 = (1'h0);
  reg [(5'h16):(1'h0)] forvar422 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg423 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar424 = (1'h0);
  reg [(5'h17):(1'h0)] reg425 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg426 = (1'h0);
  reg [(5'h13):(1'h0)] reg427 = (1'h0);
  reg [(4'hf):(1'h0)] forvar428 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg429 = (1'h0);
  reg [(3'h6):(1'h0)] reg430 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg431 = (1'h0);
  reg [(4'hc):(1'h0)] reg432 = (1'h0);
  reg [(4'hc):(1'h0)] reg422 = (1'h0);
  reg [(3'h5):(1'h0)] reg433 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg434 = (1'h0);
  reg [(5'h10):(1'h0)] reg435 = (1'h0);
  reg [(4'h8):(1'h0)] reg436 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg437 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire438;
  reg [(2'h2):(1'h0)] reg439 = (1'h0);
  reg [(5'h11):(1'h0)] forvar440 = (1'h0);
  reg [(3'h5):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg442 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg443 = (1'h0);
  reg [(4'hb):(1'h0)] reg444 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar445 = (1'h0);
  reg [(5'h10):(1'h0)] forvar446 = (1'h0);
  reg [(2'h3):(1'h0)] forvar447 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg448 = (1'h0);
  reg [(5'h14):(1'h0)] reg449 = (1'h0);
  reg [(2'h3):(1'h0)] reg450 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg451 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg452 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg453 = (1'h0);
  reg [(5'h14):(1'h0)] forvar454 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg455 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg456 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg457 = (1'h0);
  reg [(4'hb):(1'h0)] reg458 = (1'h0);
  wire [(3'h7):(1'h0)] wire459;
  reg signed [(5'h11):(1'h0)] reg460 = (1'h0);
  wire [(3'h6):(1'h0)] wire728;
  assign y = {reg748,
                 reg747,
                 reg746,
                 reg745,
                 reg744,
                 reg743,
                 reg742,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 reg735,
                 forvar734,
                 forvar733,
                 wire732,
                 reg731,
                 reg730,
                 reg401,
                 reg402,
                 forvar403,
                 reg404,
                 reg405,
                 reg406,
                 reg407,
                 reg408,
                 forvar409,
                 reg410,
                 reg411,
                 reg412,
                 reg413,
                 reg414,
                 forvar415,
                 reg416,
                 reg417,
                 reg418,
                 reg419,
                 reg420,
                 reg421,
                 forvar422,
                 reg423,
                 forvar424,
                 reg425,
                 reg426,
                 reg427,
                 forvar428,
                 reg429,
                 reg430,
                 reg431,
                 reg432,
                 reg422,
                 reg433,
                 reg434,
                 reg435,
                 reg436,
                 reg437,
                 wire438,
                 reg439,
                 forvar440,
                 reg441,
                 reg442,
                 reg443,
                 reg444,
                 forvar445,
                 forvar446,
                 forvar447,
                 reg448,
                 reg449,
                 reg450,
                 reg451,
                 reg452,
                 reg453,
                 forvar454,
                 reg455,
                 reg456,
                 reg457,
                 reg458,
                 wire459,
                 reg460,
                 wire728,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg401 <= {$unsigned((&wire396[(1'h0):(1'h0)]))};
      reg402 <= ((&{(8'ha5), {reg401}}) <<< (|(8'ha5)));
    end
  always
    @(posedge clk) begin
      for (forvar403 = (1'h0); (forvar403 < (2'h3)); forvar403 = (forvar403 + (1'h1)))
        begin
          reg404 <= (wire399[(2'h3):(2'h3)] ?
              (wire396 ?
                  {reg402[(4'hf):(3'h4)],
                      $unsigned($signed(wire396))} : ($signed(((7'h46) > reg401)) != (8'ha4))) : (8'ha4));
        end
      reg405 <= wire398[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg406 <= $unsigned((wire400 ?
          forvar403[(3'h7):(3'h4)] : (wire396[(2'h2):(2'h2)] ?
              ("owwZ4XUYbSg9WstAd1PseP" ? {reg402} : "20nQpkyoF4C7f") : "")));
      reg407 <= (reg404 ?
          $signed($signed(wire400[(4'h8):(3'h5)])) : $unsigned(($unsigned($unsigned((8'ha0))) <<< {$signed(reg404),
              "Fm8ryxBd"})));
    end
  always
    @(posedge clk) begin
      reg408 <= $signed(reg407);
      for (forvar409 = (1'h0); (forvar409 < (1'h1)); forvar409 = (forvar409 + (1'h1)))
        begin
          reg410 <= (("RO9scn" ?
              forvar403[(3'h7):(1'h1)] : $unsigned((^$signed(wire397)))) < (({(reg408 ?
                          wire397 : wire396),
                      $signed(reg401)} ?
                  reg405[(1'h1):(1'h1)] : ((~^(7'h44)) * (~&forvar409))) ?
              {$unsigned($signed(reg402)),
                  ($unsigned(reg408) ?
                      (wire396 >= reg408) : $unsigned(wire399))} : reg402));
        end
      reg411 <= $signed(wire399);
      if (((+reg410[(2'h3):(2'h2)]) >= "2bHtrTZsSRY"))
        begin
          reg412 = ((((~(reg406 - wire398)) || reg406[(4'ha):(2'h3)]) ?
                  (($signed((8'haa)) ?
                      (reg406 || wire397) : "OL") > reg404[(3'h4):(1'h1)]) : reg410) ?
              (wire399[(4'h8):(3'h7)] < wire397) : {$unsigned({reg408,
                      $unsigned(reg404)})});
        end
      else
        begin
          reg412 <= "ZK75k23aoc";
        end
      reg413 = (&($signed((8'hb9)) ? reg407 : reg404[(3'h5):(3'h5)]));
    end
  always
    @(posedge clk) begin
      reg414 <= $signed(forvar409[(2'h2):(1'h0)]);
      for (forvar415 = (1'h0); (forvar415 < (1'h0)); forvar415 = (forvar415 + (1'h1)))
        begin
          reg416 <= {(reg410[(3'h5):(3'h4)] ?
                  $unsigned($unsigned((^wire400))) : wire397[(1'h0):(1'h0)])};
          reg417 = reg402[(4'h8):(2'h3)];
          reg418 = (reg416 <= reg412);
        end
      reg419 = (+forvar403[(1'h1):(1'h1)]);
      if ("N4dOVGhuiOQ")
        begin
          reg420 <= (~^(($unsigned("x") - wire397[(1'h1):(1'h0)]) >> reg410));
          reg421 <= wire399;
          for (forvar422 = (1'h0); (forvar422 < (1'h1)); forvar422 = (forvar422 + (1'h1)))
            begin
              reg423 <= "L7";
              for (forvar424 = (1'h0); (forvar424 < (2'h3)); forvar424 = (forvar424 + (1'h1)))
                begin
                  reg425 = reg401;
                  reg426 = ($unsigned("53FRdkPyhUTvIfI") ?
                      "lmKJm2g20e4qFtO8" : ("NMBduY1" ?
                          (&($signed(forvar415) <<< {reg405})) : reg402));
                  reg427 = ("Gw2gKkMFp1km1RulHzo" ?
                      "F9H31r39aZDPUzXkgppmV" : $signed({"FbKF16O4LG3P1CdynQ9o"}));
                  for (forvar428 = (1'h0); (forvar428 < (3'h4)); forvar428 = (forvar428 + (1'h1)))
                    begin
                      reg429 <= $unsigned(((reg402 < ({wire399,
                          reg412} + (^~reg408))) < (-{{reg413, reg425},
                          (~^forvar415)})));
                    end
                  reg430 = ((reg401[(2'h3):(2'h2)] ?
                          reg429 : ($unsigned(forvar428[(3'h5):(1'h0)]) ?
                              (forvar424 << $signed(reg413)) : reg413[(3'h7):(1'h1)])) ?
                      reg423[(2'h3):(1'h1)] : $unsigned(($unsigned((8'had)) && wire399)));
                end
            end
          reg431 <= $signed((-reg404[(4'h8):(3'h7)]));
          reg432 <= ($signed(($signed({reg406}) ?
              {reg418[(1'h0):(1'h0)],
                  (~|(8'ha3))} : $unsigned($unsigned((7'h41))))) ~^ {(^$unsigned("LaZ4F3YTIy2KJ"))});
        end
      else
        begin
          reg420 <= forvar403[(4'hc):(4'hc)];
          reg421 <= (8'hb4);
          reg422 <= "m";
        end
      reg433 = ({$unsigned((reg426 ? (+forvar428) : forvar424[(2'h3):(1'h1)])),
              reg411} ?
          $signed(reg430) : $unsigned((&reg414[(2'h3):(2'h2)])));
    end
  always
    @(posedge clk) begin
      reg434 = (8'hb7);
      reg435 = (^reg419);
      reg436 <= wire396;
      reg437 <= $signed((wire400[(3'h7):(2'h3)] ?
          (($signed(wire396) <= $unsigned((8'hb4))) ?
              (~reg426) : $unsigned((reg405 ? forvar403 : reg410))) : (("yJc" ?
                  ((8'hab) ? reg433 : reg410) : reg407[(3'h6):(3'h4)]) ?
              reg418 : reg404)));
    end
  assign wire438 = {reg408};
  always
    @(posedge clk) begin
      reg439 = "QY2O";
      for (forvar440 = (1'h0); (forvar440 < (2'h3)); forvar440 = (forvar440 + (1'h1)))
        begin
          reg441 <= (^(-($unsigned({(7'h40), reg406}) ?
              $unsigned((^~reg407)) : "74Ix")));
          reg442 = (~|"IicbyCClh2uiQWMvZ");
          reg443 = (wire396[(2'h2):(1'h0)] != reg404);
        end
      reg444 <= reg401;
    end
  always
    @(posedge clk) begin
      for (forvar445 = (1'h0); (forvar445 < (2'h2)); forvar445 = (forvar445 + (1'h1)))
        begin
          for (forvar446 = (1'h0); (forvar446 < (2'h2)); forvar446 = (forvar446 + (1'h1)))
            begin
              for (forvar447 = (1'h0); (forvar447 < (2'h3)); forvar447 = (forvar447 + (1'h1)))
                begin
                  reg448 <= "DPygaKhvh0GBIdl";
                  reg449 <= reg423[(1'h1):(1'h1)];
                  reg450 <= {{wire399,
                          ($signed(reg419[(3'h5):(3'h4)]) ?
                              forvar446[(2'h3):(2'h3)] : $signed({reg430,
                                  (8'ha6)}))},
                      (reg436 ?
                          (($signed(forvar409) ?
                                  $unsigned(forvar446) : $signed(forvar409)) ?
                              (+{reg414,
                                  reg422}) : $signed("")) : wire397[(2'h2):(1'h0)])};
                end
              reg451 = (-((7'h43) ?
                  ((!(^~reg444)) ?
                      ($signed((8'hbf)) ?
                          "1g0" : $signed(reg442)) : "7iBQ") : $signed(forvar447)));
            end
          reg452 = $unsigned(($signed("26KtK") ?
              (reg449[(2'h3):(1'h0)] ?
                  (~{reg416}) : $signed($unsigned(forvar440))) : $unsigned($signed((&reg421)))));
          reg453 <= (-(($unsigned("o") ? reg401[(4'h8):(1'h0)] : reg432) ?
              ((~&reg425) ?
                  "urrZWk0CeWEARelw" : $unsigned($signed((7'h42)))) : reg416));
          for (forvar454 = (1'h0); (forvar454 < (1'h0)); forvar454 = (forvar454 + (1'h1)))
            begin
              reg455 = reg412;
              reg456 <= "N";
              reg457 = $signed({reg442[(4'ha):(4'ha)], reg432});
              reg458 = wire399;
            end
        end
    end
  assign wire459 = $unsigned((reg429[(4'hc):(4'ha)] ^ {((reg420 * (7'h46)) & $unsigned(reg432)),
                       "T8fS"}));
  always
    @(posedge clk) begin
      reg460 <= $unsigned({{"scel", $unsigned((^~wire459))}, (8'ha1)});
    end
  module461 modinst729 (.wire466(reg449), .wire464(reg419), .clk(clk), .y(wire728), .wire465(reg425), .wire463(wire397), .wire462(reg448));
  always
    @(posedge clk) begin
      reg730 <= (^("rJko9DI" * (reg452 ? forvar403 : reg402[(2'h3):(1'h1)])));
      reg731 = wire728;
    end
  assign wire732 = $signed({($unsigned((|reg434)) | {(~reg436), "Eh66"})});
  always
    @(posedge clk) begin
      for (forvar733 = (1'h0); (forvar733 < (1'h0)); forvar733 = (forvar733 + (1'h1)))
        begin
          for (forvar734 = (1'h0); (forvar734 < (1'h1)); forvar734 = (forvar734 + (1'h1)))
            begin
              reg735 <= (("5w89" ?
                      "g9oKn9yG1uaSgik" : (forvar440[(3'h4):(1'h0)] - $signed((reg420 ?
                          reg448 : reg406)))) ?
                  reg420 : {(~((wire438 ?
                          reg419 : reg451) << reg443[(2'h3):(1'h1)]))});
              reg736 <= {$signed(reg444[(1'h0):(1'h0)]),
                  (~$signed(reg413[(4'h8):(3'h5)]))};
              reg737 <= "6E";
            end
          reg738 <= ((^~$unsigned(reg414[(3'h4):(1'h1)])) ?
              $unsigned($signed($unsigned("KgDbJSJM"))) : $unsigned(reg407));
          reg739 <= forvar440[(5'h10):(1'h0)];
        end
      reg740 <= "dql";
    end
  always
    @(posedge clk) begin
      reg741 <= {forvar733};
      reg742 <= $unsigned($signed(((~|(reg436 ?
          reg444 : reg738)) == $unsigned($unsigned(forvar447)))));
      reg743 = (+((reg422 || (|{(8'ha9)})) ?
          (+{(reg430 - reg458)}) : reg457[(4'h8):(3'h6)]));
      reg744 <= "IiK";
    end
  always
    @(posedge clk) begin
      reg745 = "IHsubyDGx";
    end
  always
    @(posedge clk) begin
      reg746 <= $signed((reg739[(3'h5):(2'h3)] <<< (reg444[(3'h7):(1'h0)] ?
          reg455 : (reg456[(4'h9):(3'h5)] ? $unsigned(reg425) : (7'h43)))));
      reg747 <= reg450;
      reg748 <= reg452[(1'h1):(1'h1)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module461
#( parameter param727 = ((+(((8'ha0) ? ((7'h40) | (8'hb6)) : (^~(8'hb8))) ~^ (((8'haa) ? (7'h44) : (7'h43)) | (8'ha6)))) >>> ((((-(8'ha5)) ? ((8'ha7) || (7'h43)) : (8'hba)) ? ((~^(8'hac)) < ((8'h9e) ? (8'ha3) : (7'h46))) : {((8'hbf) != (8'hab)), ((8'ha0) ? (8'hb0) : (8'hbd))}) ? (((&(8'hbf)) ^ ((7'h44) || (7'h41))) ? ((-(8'ha5)) ? ((7'h42) >>> (7'h42)) : ((7'h48) <<< (8'h9c))) : {(-(8'hbc))}) : {({(8'hb2)} ^ {(8'hb3), (8'hb6)})})) )
(y, clk, wire466, wire465, wire464, wire463, wire462);
  output wire [(32'h789):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire466;
  input wire [(5'h17):(1'h0)] wire465;
  input wire [(3'h6):(1'h0)] wire464;
  input wire signed [(4'he):(1'h0)] wire463;
  input wire signed [(2'h3):(1'h0)] wire462;
  reg signed [(4'ha):(1'h0)] reg726 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar725 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg723 = (1'h0);
  reg signed [(4'he):(1'h0)] reg722 = (1'h0);
  reg [(5'h14):(1'h0)] reg721 = (1'h0);
  reg [(5'h12):(1'h0)] forvar720 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire719;
  wire [(3'h6):(1'h0)] wire718;
  reg [(5'h12):(1'h0)] reg717 = (1'h0);
  reg [(5'h13):(1'h0)] reg716 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg715 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg714 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg713 = (1'h0);
  reg [(5'h11):(1'h0)] reg712 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar711 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg710 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg709 = (1'h0);
  reg [(3'h6):(1'h0)] reg708 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg707 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg706 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg705 = (1'h0);
  reg [(2'h3):(1'h0)] reg704 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar703 = (1'h0);
  reg signed [(4'he):(1'h0)] reg702 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg701 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg700 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar699 = (1'h0);
  reg [(4'hf):(1'h0)] forvar698 = (1'h0);
  reg [(5'h17):(1'h0)] reg697 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg696 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg695 = (1'h0);
  reg [(3'h4):(1'h0)] reg694 = (1'h0);
  reg [(3'h7):(1'h0)] reg693 = (1'h0);
  reg [(5'h13):(1'h0)] reg692 = (1'h0);
  reg [(5'h15):(1'h0)] reg691 = (1'h0);
  reg [(5'h11):(1'h0)] reg690 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg689 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg688 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg687 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar686 = (1'h0);
  reg [(2'h3):(1'h0)] forvar685 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg685 = (1'h0);
  reg [(4'hd):(1'h0)] reg684 = (1'h0);
  reg [(4'h9):(1'h0)] reg683 = (1'h0);
  reg [(4'hd):(1'h0)] reg682 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg681 = (1'h0);
  reg [(4'hb):(1'h0)] reg680 = (1'h0);
  reg [(3'h4):(1'h0)] reg679 = (1'h0);
  reg [(3'h4):(1'h0)] reg678 = (1'h0);
  wire [(3'h5):(1'h0)] wire677;
  reg [(4'ha):(1'h0)] reg676 = (1'h0);
  reg [(4'hf):(1'h0)] reg675 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg674 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar673 = (1'h0);
  reg [(4'he):(1'h0)] reg672 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg671 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg670 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg669 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg668 = (1'h0);
  reg [(5'h10):(1'h0)] forvar667 = (1'h0);
  reg [(4'hc):(1'h0)] reg666 = (1'h0);
  reg [(2'h2):(1'h0)] forvar665 = (1'h0);
  reg [(5'h11):(1'h0)] reg664 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg663 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar662 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg661 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg660 = (1'h0);
  reg [(2'h2):(1'h0)] forvar659 = (1'h0);
  reg [(4'h9):(1'h0)] reg658 = (1'h0);
  reg [(2'h2):(1'h0)] reg657 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar656 = (1'h0);
  reg [(5'h14):(1'h0)] reg655 = (1'h0);
  reg [(3'h6):(1'h0)] reg654 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar653 = (1'h0);
  reg signed [(4'he):(1'h0)] reg652 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg651 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar650 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar649 = (1'h0);
  reg [(4'hd):(1'h0)] reg648 = (1'h0);
  reg [(5'h14):(1'h0)] reg647 = (1'h0);
  reg [(4'hd):(1'h0)] reg646 = (1'h0);
  wire signed [(4'he):(1'h0)] wire545;
  reg signed [(4'he):(1'h0)] reg506 = (1'h0);
  reg [(3'h4):(1'h0)] reg505 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg504 = (1'h0);
  reg [(4'ha):(1'h0)] reg503 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg502 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar501 = (1'h0);
  reg [(4'he):(1'h0)] reg500 = (1'h0);
  reg [(3'h7):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar498 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar497 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg496 = (1'h0);
  reg [(4'he):(1'h0)] reg495 = (1'h0);
  reg [(5'h10):(1'h0)] reg494 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar493 = (1'h0);
  reg [(3'h4):(1'h0)] reg492 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg491 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg490 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg489 = (1'h0);
  reg [(5'h12):(1'h0)] reg488 = (1'h0);
  reg [(4'hd):(1'h0)] reg487 = (1'h0);
  reg [(5'h11):(1'h0)] reg486 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg485 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg484 = (1'h0);
  reg [(4'hf):(1'h0)] reg483 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg482 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg481 = (1'h0);
  reg [(3'h6):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar479 = (1'h0);
  reg [(5'h16):(1'h0)] reg478 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire477;
  reg [(2'h3):(1'h0)] reg476 = (1'h0);
  reg [(5'h17):(1'h0)] reg475 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg474 = (1'h0);
  reg [(4'hb):(1'h0)] reg473 = (1'h0);
  reg [(5'h12):(1'h0)] reg472 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg471 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg470 = (1'h0);
  reg [(5'h14):(1'h0)] forvar469 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar468 = (1'h0);
  reg [(3'h5):(1'h0)] reg467 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar547 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg548 = (1'h0);
  reg [(4'he):(1'h0)] forvar549 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg550 = (1'h0);
  reg [(5'h14):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg552 = (1'h0);
  reg [(5'h14):(1'h0)] reg553 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg554 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg555 = (1'h0);
  reg [(4'he):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg557 = (1'h0);
  reg signed [(4'he):(1'h0)] reg558 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar559 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg560 = (1'h0);
  reg [(3'h7):(1'h0)] forvar561 = (1'h0);
  reg [(4'hf):(1'h0)] reg562 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar563 = (1'h0);
  reg [(4'hd):(1'h0)] reg564 = (1'h0);
  reg [(4'hb):(1'h0)] reg565 = (1'h0);
  reg [(2'h3):(1'h0)] reg566 = (1'h0);
  reg [(3'h6):(1'h0)] forvar567 = (1'h0);
  reg [(5'h13):(1'h0)] reg568 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar569 = (1'h0);
  reg [(5'h10):(1'h0)] reg570 = (1'h0);
  reg signed [(4'he):(1'h0)] reg571 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg572 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire573;
  wire [(4'hd):(1'h0)] wire574;
  reg [(4'hb):(1'h0)] forvar575 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg576 = (1'h0);
  wire [(4'hd):(1'h0)] wire644;
  assign y = {reg726,
                 forvar725,
                 reg724,
                 reg723,
                 reg722,
                 reg721,
                 forvar720,
                 wire719,
                 wire718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 reg713,
                 reg712,
                 forvar711,
                 reg710,
                 reg709,
                 reg708,
                 reg707,
                 reg706,
                 reg705,
                 reg704,
                 forvar703,
                 reg702,
                 reg701,
                 reg700,
                 forvar699,
                 forvar698,
                 reg697,
                 reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 reg691,
                 reg690,
                 reg689,
                 reg688,
                 reg687,
                 forvar686,
                 forvar685,
                 reg685,
                 reg684,
                 reg683,
                 reg682,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 wire677,
                 reg676,
                 reg675,
                 reg674,
                 forvar673,
                 reg672,
                 reg671,
                 reg670,
                 reg669,
                 reg668,
                 forvar667,
                 reg666,
                 forvar665,
                 reg664,
                 reg663,
                 forvar662,
                 reg661,
                 reg660,
                 forvar659,
                 reg658,
                 reg657,
                 forvar656,
                 reg655,
                 reg654,
                 forvar653,
                 reg652,
                 reg651,
                 forvar650,
                 forvar649,
                 reg648,
                 reg647,
                 reg646,
                 wire545,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 forvar501,
                 reg500,
                 reg499,
                 forvar498,
                 forvar497,
                 reg496,
                 reg495,
                 reg494,
                 forvar493,
                 reg492,
                 reg491,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 forvar479,
                 reg478,
                 wire477,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 forvar469,
                 forvar468,
                 reg467,
                 forvar547,
                 reg548,
                 forvar549,
                 reg550,
                 reg551,
                 reg552,
                 reg553,
                 reg554,
                 reg555,
                 reg556,
                 reg557,
                 reg558,
                 forvar559,
                 reg560,
                 forvar561,
                 reg562,
                 forvar563,
                 reg564,
                 reg565,
                 reg566,
                 forvar567,
                 reg568,
                 forvar569,
                 reg570,
                 reg571,
                 reg572,
                 wire573,
                 wire574,
                 forvar575,
                 reg576,
                 wire644,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg467 = $signed({wire462, "iYpIgt9YyL9q"});
      for (forvar468 = (1'h0); (forvar468 < (2'h2)); forvar468 = (forvar468 + (1'h1)))
        begin
          for (forvar469 = (1'h0); (forvar469 < (1'h0)); forvar469 = (forvar469 + (1'h1)))
            begin
              reg470 <= $signed($unsigned(wire463[(4'h8):(2'h2)]));
            end
          reg471 <= ({(wire464 < ((wire463 << wire464) ?
                      reg467[(3'h4):(2'h2)] : wire463[(3'h7):(1'h0)]))} ?
              wire462 : ($signed((~forvar469)) || reg467));
        end
      reg472 <= "hKpk";
    end
  always
    @(posedge clk) begin
      reg473 <= (wire465[(2'h2):(1'h0)] || ($unsigned((forvar469 ?
              (~^forvar469) : {reg470, reg471})) ?
          "HcJDt" : (forvar469[(1'h1):(1'h1)] > (((8'ha4) ?
              reg467 : wire464) * $signed(wire465)))));
      reg474 <= reg473;
      reg475 <= (8'hab);
      if (reg470[(4'h9):(4'h9)])
        begin
          reg476 <= ((("h4ge4" ?
                  (reg470[(1'h1):(1'h0)] ?
                      wire463[(2'h3):(1'h1)] : (reg475 ?
                          reg470 : (8'hb8))) : $unsigned(reg467)) << wire465[(5'h12):(4'h8)]) ?
              ("GANmFD" ?
                  (reg473 ^~ $unsigned(reg474)) : (!($unsigned(wire463) * (reg467 >>> reg475)))) : "Ph5");
        end
      else
        begin
          reg476 <= reg470[(1'h1):(1'h0)];
        end
    end
  assign wire477 = $unsigned($unsigned(("9k35NPcWE5avsvwvN" ?
                       ($unsigned(forvar468) ?
                           (~&(8'haf)) : (8'hab)) : (8'hb3))));
  always
    @(posedge clk) begin
      reg478 <= $signed($signed((wire463 ? reg471[(2'h2):(1'h1)] : wire463)));
      for (forvar479 = (1'h0); (forvar479 < (3'h4)); forvar479 = (forvar479 + (1'h1)))
        begin
          reg480 = $unsigned({((&(wire466 <= wire462)) >= wire477), reg478});
          reg481 <= reg474[(1'h1):(1'h0)];
          reg482 <= "iwrcvmrg2ZW6eOdecRtE8p";
          reg483 <= ("9fTk8549Vcat9Y1gUCffA" ^ reg473[(2'h2):(1'h1)]);
          reg484 <= forvar468;
        end
      reg485 = reg481[(3'h6):(1'h1)];
      reg486 = {wire477, $unsigned("aHAmsLY2goH4Rvq8")};
    end
  always
    @(posedge clk) begin
      reg487 <= (+wire463[(4'h9):(1'h1)]);
      reg488 = reg471[(4'ha):(3'h5)];
    end
  always
    @(posedge clk) begin
      reg489 <= wire462;
      reg490 <= (~&(-"I"));
      reg491 <= ("m8X2" || reg475[(5'h15):(4'h9)]);
    end
  always
    @(posedge clk) begin
      reg492 <= (~&$unsigned($signed("41aHcgEypOA6EV2fYAizqt")));
    end
  always
    @(posedge clk) begin
      for (forvar493 = (1'h0); (forvar493 < (3'h4)); forvar493 = (forvar493 + (1'h1)))
        begin
          reg494 <= (("ykH8xa91Nh" ?
                  wire464[(1'h1):(1'h1)] : ("OwpR" | reg475)) ?
              {(reg486 && reg478[(2'h3):(1'h0)])} : $unsigned("GOmgKRwPoq"));
          reg495 <= (((~|"d") << $signed(reg478)) & ((^reg489[(1'h0):(1'h0)]) ?
              $signed($signed($signed(wire462))) : (($unsigned(reg494) ?
                      (wire466 - (8'hb8)) : (reg472 ? reg482 : forvar469)) ?
                  (8'hb5) : "")));
          reg496 = {$signed($unsigned($unsigned("1fVtWzBASzoW")))};
          for (forvar497 = (1'h0); (forvar497 < (2'h3)); forvar497 = (forvar497 + (1'h1)))
            begin
              for (forvar498 = (1'h0); (forvar498 < (1'h0)); forvar498 = (forvar498 + (1'h1)))
                begin
                  reg499 = $unsigned(reg485[(1'h0):(1'h0)]);
                  reg500 = (^~(!"YMQmH8rYYZ"));
                  for (forvar501 = (1'h0); (forvar501 < (3'h4)); forvar501 = (forvar501 + (1'h1)))
                    begin
                      reg502 = reg490;
                    end
                end
              reg503 <= $unsigned(($signed("S1fegOKe9KKG") - forvar469));
            end
        end
      reg504 = reg480[(3'h6):(3'h5)];
      reg505 <= (($signed(((reg476 ? reg502 : reg485) & (reg472 ?
              reg502 : (8'haf)))) * reg475) ?
          reg470 : $unsigned((^$unsigned("CEkhPKkKuLrcFJID"))));
      reg506 <= ($unsigned("bpmCeMHhQTDgaD") ?
          (&{{forvar497, forvar497[(4'ha):(3'h6)]}, reg489}) : reg472);
    end
  module507 modinst546 (wire545, clk, forvar498, wire466, reg471, forvar469, reg500);
  always
    @(posedge clk) begin
      for (forvar547 = (1'h0); (forvar547 < (2'h3)); forvar547 = (forvar547 + (1'h1)))
        begin
          reg548 <= ($unsigned($unsigned((wire463[(4'hd):(4'ha)] << reg475))) <= $signed(("LvGM" ?
              reg496 : (reg504 >> $signed(reg500)))));
          for (forvar549 = (1'h0); (forvar549 < (2'h3)); forvar549 = (forvar549 + (1'h1)))
            begin
              reg550 <= ($unsigned(($unsigned($signed((8'ha0))) + (^(-reg473)))) | forvar498);
              reg551 <= reg490[(3'h4):(2'h2)];
            end
        end
      reg552 <= (~&{reg476,
          (reg551[(2'h3):(2'h2)] || forvar501[(1'h0):(1'h0)])});
      reg553 <= ((reg473 ?
              (|((^(8'haa)) <= $signed(forvar501))) : "GktOibIcit1KxYzJ92x7") ?
          reg548 : wire466);
    end
  always
    @(posedge clk) begin
      reg554 <= ($signed($unsigned((~^{(7'h45), (7'h47)}))) ^ (8'ha9));
      if ("vVimEzXtZ5TT")
        begin
          reg555 <= ((wire463 | (reg492 && $unsigned({forvar493}))) < reg554[(4'h8):(3'h5)]);
          reg556 <= $signed($unsigned((^~($signed(reg483) ?
              (|(8'ha3)) : "AnC9YQLR7WPxWJOhSvYb40"))));
          reg557 <= $signed((reg478[(1'h0):(1'h0)] ?
              reg552[(4'h9):(3'h6)] : {(reg552 ? ((8'hac) | wire465) : reg470),
                  {$signed(wire464)}}));
          reg558 <= $signed(forvar498[(3'h5):(1'h0)]);
          for (forvar559 = (1'h0); (forvar559 < (1'h0)); forvar559 = (forvar559 + (1'h1)))
            begin
              reg560 <= (~"RIftVNF91lxDY9Gq");
              for (forvar561 = (1'h0); (forvar561 < (1'h0)); forvar561 = (forvar561 + (1'h1)))
                begin
                  reg562 <= (7'h41);
                  for (forvar563 = (1'h0); (forvar563 < (3'h4)); forvar563 = (forvar563 + (1'h1)))
                    begin
                      reg564 <= (&{(((^~reg494) <<< ((7'h44) ?
                                  (8'hb3) : reg500)) ?
                              (8'ha5) : ((forvar547 & (8'hb1)) ~^ "")),
                          (reg484[(2'h2):(2'h2)] ?
                              ($unsigned(reg552) ?
                                  reg553 : $signed(reg472)) : {$signed(reg560)})});
                      reg565 = $signed("toctSUVQYbHEuaZufQxv0");
                      reg566 = $signed($unsigned(forvar493));
                    end
                end
              for (forvar567 = (1'h0); (forvar567 < (2'h3)); forvar567 = (forvar567 + (1'h1)))
                begin
                  reg568 <= ($unsigned((reg554[(4'hd):(4'hc)] ?
                          reg556 : reg470)) ?
                      (|$signed({$signed(reg485)})) : (forvar498 ?
                          (forvar468[(4'h8):(3'h4)] ?
                              reg482[(4'hf):(2'h3)] : ("7F1EYJb" ?
                                  ((8'hae) ~^ reg551) : reg487[(3'h7):(3'h6)])) : "SUvziDChCsLzLTbr"));
                end
              for (forvar569 = (1'h0); (forvar569 < (3'h4)); forvar569 = (forvar569 + (1'h1)))
                begin
                  reg570 = $unsigned("YGJOH61DD5gH");
                  reg571 <= $unsigned(("R6eYBVIGMLzbKn2nw" ?
                      $unsigned((+(reg487 >>> (8'hb0)))) : (reg487[(4'h9):(1'h1)] + "ZEG2df")));
                end
              reg572 = reg484;
            end
        end
      else
        begin
          reg555 = ($unsigned((7'h42)) ?
              (forvar468[(2'h2):(2'h2)] | {reg564[(4'hb):(1'h1)]}) : "dlZiqDTaWg9nZGLog0bC");
          reg556 <= forvar547;
        end
    end
  assign wire573 = forvar549[(1'h0):(1'h0)];
  assign wire574 = $unsigned(forvar497[(2'h3):(1'h1)]);
  always
    @(posedge clk) begin
      for (forvar575 = (1'h0); (forvar575 < (2'h2)); forvar575 = (forvar575 + (1'h1)))
        begin
          reg576 = ($unsigned(reg565[(3'h5):(1'h1)]) ?
              (reg557 <<< wire463[(4'he):(3'h7)]) : forvar498[(4'h9):(1'h0)]);
        end
    end
  module577 modinst645 (.y(wire644), .clk(clk), .wire582(reg473), .wire581(reg470), .wire578(reg550), .wire580(reg491), .wire579(forvar493));
  always
    @(posedge clk) begin
      reg646 <= (reg489[(4'h9):(3'h6)] ~^ reg562[(3'h6):(1'h0)]);
      reg647 = "C5";
      reg648 <= reg486[(2'h3):(2'h2)];
    end
  always
    @(posedge clk) begin
      for (forvar649 = (1'h0); (forvar649 < (2'h3)); forvar649 = (forvar649 + (1'h1)))
        begin
          for (forvar650 = (1'h0); (forvar650 < (2'h2)); forvar650 = (forvar650 + (1'h1)))
            begin
              reg651 <= (((7'h43) & forvar649) | "CNSbE4ipLXFeS4");
              reg652 <= "";
              for (forvar653 = (1'h0); (forvar653 < (2'h2)); forvar653 = (forvar653 + (1'h1)))
                begin
                  reg654 <= (8'hac);
                end
              reg655 <= ({$unsigned(reg652[(2'h3):(1'h1)]),
                      $unsigned(((reg557 ?
                          reg562 : (8'ha1)) >> $unsigned(reg495)))} ?
                  "DkhSJE5oto" : {($unsigned(reg551[(3'h7):(1'h1)]) ?
                          $signed($unsigned(reg492)) : "EwXE7C1DOmIUt"),
                      reg560[(1'h0):(1'h0)]});
              for (forvar656 = (1'h0); (forvar656 < (1'h0)); forvar656 = (forvar656 + (1'h1)))
                begin
                  reg657 = reg565[(3'h7):(2'h3)];
                end
            end
          reg658 <= $signed($signed((|"gOzJAlGzLUOP3JKW")));
        end
      for (forvar659 = (1'h0); (forvar659 < (3'h4)); forvar659 = (forvar659 + (1'h1)))
        begin
          reg660 <= reg489[(4'h9):(2'h2)];
          reg661 <= {$signed(reg572), "2q"};
          for (forvar662 = (1'h0); (forvar662 < (1'h0)); forvar662 = (forvar662 + (1'h1)))
            begin
              reg663 <= {$unsigned((^reg504))};
              reg664 = $signed(reg478[(4'h8):(3'h7)]);
              for (forvar665 = (1'h0); (forvar665 < (1'h0)); forvar665 = (forvar665 + (1'h1)))
                begin
                  reg666 <= {$unsigned("4NC6kHK5Q")};
                  for (forvar667 = (1'h0); (forvar667 < (3'h4)); forvar667 = (forvar667 + (1'h1)))
                    begin
                      reg668 <= reg506;
                      reg669 <= reg485[(4'ha):(4'h9)];
                    end
                  reg670 <= (-((reg506 ?
                          $signed(reg485) : (-$unsigned(wire573))) ?
                      $unsigned($unsigned((reg487 ?
                          (8'haf) : wire574))) : $signed($unsigned(reg657[(2'h2):(2'h2)]))));
                  reg671 <= $unsigned(wire573);
                end
            end
          reg672 <= "vsUyoEzmU96sDgvZQIt";
          for (forvar673 = (1'h0); (forvar673 < (1'h0)); forvar673 = (forvar673 + (1'h1)))
            begin
              reg674 = $signed(reg492[(1'h0):(1'h0)]);
              reg675 = "ZE2p4tvfk4L";
              reg676 <= $unsigned($signed($unsigned("4d8qrXVb")));
            end
        end
    end
  assign wire677 = (&{($signed((reg565 ? forvar575 : forvar665)) ^~ (((8'ha2) ?
                           (8'had) : reg570) != "DYLtP0NSPdHkek"))});
  always
    @(posedge clk) begin
      reg678 <= {"NAr4fDKhl0kywiWU5vdb", $unsigned((^~(^~$unsigned(reg500))))};
      reg679 = reg486;
      reg680 <= $unsigned(reg568);
      reg681 <= reg504;
    end
  always
    @(posedge clk) begin
      reg682 <= $unsigned(reg664);
      reg683 = {$unsigned((reg483 != (reg565[(2'h3):(1'h1)] < (forvar667 + reg475))))};
      reg684 <= (~|(!((reg562[(4'hf):(2'h2)] ? {reg675} : {(8'ha6), reg668}) ?
          reg555[(1'h1):(1'h0)] : $unsigned(forvar665[(1'h1):(1'h0)]))));
      if ((^~$unsigned((wire477 != (^{wire644})))))
        begin
          reg685 = "N";
        end
      else
        begin
          for (forvar685 = (1'h0); (forvar685 < (1'h0)); forvar685 = (forvar685 + (1'h1)))
            begin
              for (forvar686 = (1'h0); (forvar686 < (1'h1)); forvar686 = (forvar686 + (1'h1)))
                begin
                  reg687 = reg499[(3'h6):(1'h0)];
                end
              reg688 <= reg505;
              reg689 <= "4Ryk";
              reg690 <= ("5" ?
                  $unsigned($signed($unsigned(reg485[(4'h8):(3'h5)]))) : $signed(($signed("gaap9y8guaaSlkZTq4Guwt") ?
                      reg558 : {"JgF4b"})));
            end
          reg691 = {wire573[(2'h3):(1'h0)], (|reg486[(2'h2):(1'h1)])};
          reg692 = ("oum2KFvD43QBS" ?
              "2GSRhIBgv1625SyY5w" : $signed($signed($signed("07LJgbE8OQlxpkbE"))));
          reg693 = (~"9QzNFWawxG5");
        end
      reg694 <= (forvar567 ?
          (|($unsigned($unsigned(forvar649)) < reg571)) : forvar468[(3'h7):(3'h7)]);
    end
  always
    @(posedge clk) begin
      reg695 <= ($signed("e4GCf") ? reg671 : (!{("U0" || $unsigned((8'hb9)))}));
      reg696 <= ("B9UKJBo9Evc4Z5yN5fTn1" ^ ($unsigned((|$unsigned(reg505))) >= $unsigned($unsigned(((8'hb5) ?
          reg672 : reg692)))));
      reg697 = $signed(reg679[(2'h2):(2'h2)]);
      for (forvar698 = (1'h0); (forvar698 < (1'h0)); forvar698 = (forvar698 + (1'h1)))
        begin
          for (forvar699 = (1'h0); (forvar699 < (2'h3)); forvar699 = (forvar699 + (1'h1)))
            begin
              if (reg478)
                begin
                  reg700 <= (~forvar650[(3'h6):(1'h1)]);
                  reg701 <= $signed((^$signed((reg499[(1'h0):(1'h0)] ?
                      reg564[(2'h3):(1'h0)] : $unsigned(reg647)))));
                  reg702 = {(^{((&(8'hbe)) ^ {(8'ha9), reg504}),
                          "gdU3rv6HUfc"})};
                  for (forvar703 = (1'h0); (forvar703 < (1'h1)); forvar703 = (forvar703 + (1'h1)))
                    begin
                      reg704 <= reg565[(2'h3):(1'h1)];
                      reg705 <= (~{$signed(((reg694 - reg702) ?
                              (reg487 ? reg475 : forvar549) : (~^(7'h41)))),
                          ($unsigned($signed(reg691)) ?
                              forvar498[(5'h13):(4'h9)] : $signed(reg491))});
                      reg706 <= (8'ha3);
                    end
                  reg707 <= (^$signed(reg689));
                end
              else
                begin
                  reg700 <= (((7'h42) ^~ "Dgma70gAuo") < "OTqOxe1qUpWC");
                end
              reg708 <= $signed("ag5SOMy16xMDMn");
              reg709 <= (^"w45DmRmMQH3zBApkRh");
              reg710 <= $unsigned({$signed($unsigned(""))});
              for (forvar711 = (1'h0); (forvar711 < (3'h4)); forvar711 = (forvar711 + (1'h1)))
                begin
                  if ({(reg661 ?
                          ($unsigned("Z9QArWhYfnoQVGOrYt") - forvar662[(4'ha):(4'h9)]) : forvar656),
                      wire573})
                    begin
                      reg712 = (7'h46);
                    end
                  else
                    begin
                      reg712 = (reg661[(3'h5):(2'h3)] ^ ((7'h41) <= (($signed((8'h9e)) - reg666) ?
                          {(reg472 <<< (8'hb1))} : (-reg706))));
                    end
                  reg713 <= reg712[(5'h11):(1'h0)];
                end
            end
          reg714 <= (~&reg660);
        end
    end
  always
    @(posedge clk) begin
      reg715 = (reg652[(3'h6):(3'h6)] > reg496);
      reg716 = ("HYnTIiRySC" ?
          "KAQ8K70GlElaQ8" : (reg646[(4'hd):(1'h0)] != (~|((reg669 ?
                  (8'h9d) : reg647) ?
              forvar685[(1'h1):(1'h1)] : "99sAvX"))));
      reg717 <= $signed("");
    end
  assign wire718 = (("6AA6xeX8u" ? "ZMkrG" : "lCc") ? forvar498 : "1s04F4A951");
  assign wire719 = (("ftKc6qNo" ?
                       ((((8'hbc) && reg476) & {forvar665,
                           (8'ha7)}) | (7'h43)) : $unsigned($signed((forvar703 ?
                           reg669 : wire464)))) ^~ "kAZJqZtdaJA19v");
  always
    @(posedge clk) begin
      for (forvar720 = (1'h0); (forvar720 < (1'h1)); forvar720 = (forvar720 + (1'h1)))
        begin
          reg721 <= $unsigned(({(7'h42)} * (~&"sUCDI7wravH9J")));
          reg722 <= $signed($unsigned($signed($signed($unsigned((8'hb7))))));
          reg723 = (&(((reg693[(2'h3):(2'h2)] ?
                  (reg664 > reg683) : ((8'ha4) != reg476)) ?
              (((7'h43) ?
                  (8'ha1) : reg557) & $unsigned(forvar667)) : ("ywd2HiSJCb" >= ((8'ha2) >>> (8'haa)))) >= (reg490[(1'h1):(1'h0)] ?
              (!(reg702 ? reg562 : forvar498)) : forvar569[(2'h3):(2'h3)])));
          reg724 = $unsigned(reg482[(4'ha):(4'h9)]);
        end
      for (forvar725 = (1'h0); (forvar725 < (1'h1)); forvar725 = (forvar725 + (1'h1)))
        begin
          reg726 <= $unsigned((|forvar662[(1'h0):(1'h0)]));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module577
#( parameter param642 = (^(~|({((7'h40) ? (8'hba) : (8'h9e)), (^~(8'ha6))} <<< (~^(~(8'hbd))))))
, parameter param643 = {(^(^((param642 ? (8'had) : param642) && (~&param642)))), ((~(~&(^param642))) ? (~(~|(~|param642))) : (-(~&(param642 >> param642))))} )
(y, clk, wire582, wire581, wire580, wire579, wire578);
  output wire [(32'h2e9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire582;
  input wire signed [(5'h16):(1'h0)] wire581;
  input wire signed [(4'hf):(1'h0)] wire580;
  input wire [(4'hc):(1'h0)] wire579;
  input wire signed [(4'h8):(1'h0)] wire578;
  reg signed [(5'h12):(1'h0)] reg641 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar640 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg639 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg638 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg637 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg636 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar635 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg634 = (1'h0);
  reg [(5'h10):(1'h0)] reg633 = (1'h0);
  reg [(3'h7):(1'h0)] reg632 = (1'h0);
  reg [(4'ha):(1'h0)] reg631 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg630 = (1'h0);
  reg [(3'h4):(1'h0)] reg629 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar628 = (1'h0);
  reg [(2'h3):(1'h0)] reg627 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg626 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg625 = (1'h0);
  reg [(5'h10):(1'h0)] reg624 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar623 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire622;
  reg signed [(4'hb):(1'h0)] reg621 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg620 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg619 = (1'h0);
  reg [(5'h10):(1'h0)] reg618 = (1'h0);
  reg [(3'h6):(1'h0)] reg617 = (1'h0);
  reg [(5'h17):(1'h0)] reg616 = (1'h0);
  reg [(5'h14):(1'h0)] reg615 = (1'h0);
  reg [(5'h13):(1'h0)] forvar614 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg613 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar612 = (1'h0);
  reg [(5'h14):(1'h0)] reg611 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg610 = (1'h0);
  reg [(5'h13):(1'h0)] reg609 = (1'h0);
  reg [(4'hc):(1'h0)] reg608 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg607 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar606 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg605 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg604 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg603 = (1'h0);
  reg [(3'h7):(1'h0)] reg602 = (1'h0);
  reg [(5'h16):(1'h0)] reg601 = (1'h0);
  reg [(5'h13):(1'h0)] forvar600 = (1'h0);
  reg [(2'h2):(1'h0)] reg599 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg598 = (1'h0);
  reg [(5'h10):(1'h0)] reg597 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg596 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg595 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg594 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg593 = (1'h0);
  reg [(5'h13):(1'h0)] reg592 = (1'h0);
  reg [(2'h3):(1'h0)] reg591 = (1'h0);
  reg [(3'h7):(1'h0)] forvar590 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg589 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg588 = (1'h0);
  reg [(4'h9):(1'h0)] reg587 = (1'h0);
  reg [(5'h14):(1'h0)] reg586 = (1'h0);
  reg [(3'h5):(1'h0)] forvar585 = (1'h0);
  reg [(5'h14):(1'h0)] forvar584 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg583 = (1'h0);
  assign y = {reg641,
                 forvar640,
                 reg639,
                 reg638,
                 reg637,
                 reg636,
                 forvar635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 reg630,
                 reg629,
                 forvar628,
                 reg627,
                 reg626,
                 reg625,
                 reg624,
                 forvar623,
                 wire622,
                 reg621,
                 reg620,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 reg615,
                 forvar614,
                 reg613,
                 forvar612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 forvar606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 forvar600,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 forvar590,
                 reg589,
                 reg588,
                 reg587,
                 reg586,
                 forvar585,
                 forvar584,
                 reg583,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg583 <= wire578;
      for (forvar584 = (1'h0); (forvar584 < (2'h3)); forvar584 = (forvar584 + (1'h1)))
        begin
          for (forvar585 = (1'h0); (forvar585 < (2'h3)); forvar585 = (forvar585 + (1'h1)))
            begin
              reg586 <= {{"Zr6rJzYxJl",
                      ((+(wire578 <<< wire582)) || ((forvar584 ?
                          (7'h41) : wire582) | (^~forvar584)))},
                  $unsigned(((~^$signed(wire581)) ?
                      wire579 : ((&wire578) ?
                          (+(8'h9e)) : (forvar584 ? wire579 : (8'hb1)))))};
            end
          if (wire581)
            begin
              reg587 = "g77aIIRg0sJKz4yA";
            end
          else
            begin
              reg587 = "ULDpvEma0";
              reg588 <= $unsigned($unsigned((8'ha5)));
              reg589 = (^~wire580[(4'hf):(3'h4)]);
              for (forvar590 = (1'h0); (forvar590 < (2'h2)); forvar590 = (forvar590 + (1'h1)))
                begin
                  reg591 <= "Keu2Aq9G8EaLsg";
                end
            end
          reg592 <= ($signed((+{(reg587 ~^ wire579)})) ^~ $unsigned(((reg588 || (reg587 >>> wire582)) > {"OEfom",
              $unsigned(forvar585)})));
          reg593 <= reg588;
          reg594 <= ({(({reg583, forvar585} + (^(8'h9f))) ?
                  "Ny" : $signed((wire579 > reg591))),
              (((+reg583) ?
                  (reg593 ?
                      reg593 : reg592) : "WVV0xBk2") - (-"a"))} & $signed(reg592));
        end
      reg595 = wire582;
    end
  always
    @(posedge clk) begin
      reg596 = reg583[(1'h0):(1'h0)];
      reg597 <= (&(^~((~|$signed(reg595)) ?
          wire578 : ($unsigned(reg586) ?
              (forvar590 < reg592) : (reg589 * (8'hb0))))));
      reg598 <= "b7QP0WBy7GT6smFDLzV";
    end
  always
    @(posedge clk) begin
      reg599 <= $signed(wire578[(2'h3):(1'h1)]);
      for (forvar600 = (1'h0); (forvar600 < (2'h3)); forvar600 = (forvar600 + (1'h1)))
        begin
          reg601 = (~&"YBx1hFhntd0u");
        end
      reg602 = $signed($signed({{reg601[(4'ha):(3'h7)]}}));
    end
  always
    @(posedge clk) begin
      reg603 <= reg586[(4'hf):(3'h4)];
      reg604 = (wire582[(2'h3):(1'h0)] + (+($signed("DXPU") < $unsigned(reg591))));
      reg605 = $signed($signed(((8'haa) ?
          $unsigned({wire582, wire581}) : wire582[(1'h1):(1'h1)])));
      for (forvar606 = (1'h0); (forvar606 < (1'h1)); forvar606 = (forvar606 + (1'h1)))
        begin
          reg607 <= (reg602[(2'h2):(1'h1)] ?
              reg597[(4'hd):(4'hc)] : (reg605 ?
                  reg604 : (($signed(wire581) <= "BhcaCnFPRih") ?
                      ("8sx5zT" ?
                          "BC16GBQk" : $signed(wire582)) : $unsigned($signed((8'haf))))));
          reg608 <= $unsigned(((reg588 ~^ ({forvar585,
                  forvar585} ^~ $unsigned((7'h47)))) ?
              ("s9NeQQ" ?
                  (forvar600 >= (~|wire581)) : $unsigned($signed(reg598))) : (!(|((8'hbd) ?
                  (8'ha7) : forvar606)))));
        end
    end
  always
    @(posedge clk) begin
      reg609 <= (8'ha0);
      reg610 <= (+(~(((reg604 ? (7'h44) : reg597) ?
              $unsigned((7'h44)) : (&forvar585)) ?
          $unsigned({reg604, reg609}) : "opLPIuHJAnLiNxhlfJD")));
      reg611 <= $unsigned((reg598 >>> "Q9Ypc7IXQ3Lyn"));
      for (forvar612 = (1'h0); (forvar612 < (1'h0)); forvar612 = (forvar612 + (1'h1)))
        begin
          reg613 <= wire578[(3'h4):(2'h2)];
          for (forvar614 = (1'h0); (forvar614 < (2'h3)); forvar614 = (forvar614 + (1'h1)))
            begin
              reg615 <= (|(reg599 ?
                  reg609[(4'he):(4'hb)] : $unsigned((8'ha7))));
              reg616 <= $unsigned(forvar590[(2'h3):(1'h0)]);
              reg617 = $unsigned(({"qZDQ3fquHchTGKu", (~$signed(reg609))} ?
                  reg603 : $signed("wvrw7FEDQcsm2mL")));
              reg618 <= reg587[(2'h3):(1'h1)];
            end
          reg619 <= $signed({(forvar585 ?
                  reg592 : {reg608, "IKq04P9SeJl71BEnPi"}),
              reg593});
          reg620 <= reg596[(2'h2):(2'h2)];
        end
      reg621 <= $signed((8'ha6));
    end
  assign wire622 = (~^(reg593[(4'hf):(4'ha)] >= reg615[(5'h11):(1'h0)]));
  always
    @(posedge clk) begin
      for (forvar623 = (1'h0); (forvar623 < (2'h3)); forvar623 = (forvar623 + (1'h1)))
        begin
          reg624 <= ((~&(forvar584 ^~ ((^~(8'hbd)) ?
              $signed(wire582) : (7'h46)))) < (((8'hb6) ?
                  $unsigned((~|forvar590)) : "pJEacm9i4GTL5mF") ?
              (reg621 ^~ (8'ha6)) : reg609));
          reg625 = reg596;
        end
      reg626 <= (~|reg604[(2'h3):(2'h3)]);
    end
  always
    @(posedge clk) begin
      reg627 <= "uRQ7f";
      for (forvar628 = (1'h0); (forvar628 < (1'h1)); forvar628 = (forvar628 + (1'h1)))
        begin
          reg629 = reg603[(3'h5):(1'h1)];
          reg630 <= (($unsigned("CzFOWqRkqpUy7o5Dy") ?
                  ($signed($signed(wire580)) || reg603) : $signed(((reg605 ?
                      (7'h44) : reg625) && (reg621 ? reg607 : reg611)))) ?
              $unsigned({($signed(reg625) ~^ "ydO6HHe1nXeUkInrHYwK")}) : wire579[(4'ha):(3'h6)]);
          reg631 = $signed(reg599);
          reg632 <= (8'ha7);
        end
    end
  always
    @(posedge clk) begin
      reg633 <= (wire578 + ((($unsigned(reg627) ?
                  (reg630 >> reg619) : (-reg621)) ?
              ((reg630 ? reg601 : reg615) ?
                  wire579[(4'h9):(4'h8)] : reg618[(4'hc):(4'h9)]) : (-reg599)) ?
          $unsigned(($unsigned(forvar623) >= $signed((8'hb5)))) : {{(wire578 ?
                      reg610 : (8'hb1))},
              ((reg625 == (8'ha1)) ? forvar590 : {reg611, reg629})}));
    end
  always
    @(posedge clk) begin
      reg634 <= ($signed(((8'ha2) > "9VygbQwr1")) * $unsigned((|$signed($unsigned(reg603)))));
      for (forvar635 = (1'h0); (forvar635 < (1'h1)); forvar635 = (forvar635 + (1'h1)))
        begin
          reg636 <= {reg615[(5'h13):(4'h9)], reg599};
          reg637 <= $unsigned(((-forvar600[(1'h0):(1'h0)]) ?
              (7'h46) : $unsigned(reg593[(3'h4):(1'h1)])));
          reg638 = (^~reg632);
        end
    end
  always
    @(posedge clk) begin
      reg639 = {$signed((reg632 == (&"gad17UYN2zxoM2UlbKEo")))};
      for (forvar640 = (1'h0); (forvar640 < (2'h3)); forvar640 = (forvar640 + (1'h1)))
        begin
          reg641 <= (-$unsigned(reg613[(4'hf):(4'hc)]));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module507
#( parameter param543 = (+(+(!((~^(7'h43)) ^ (~(7'h46))))))
, parameter param544 = (8'ha2) )
(y, clk, wire512, wire511, wire510, wire509, wire508);
  output wire [(32'h162):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire512;
  input wire [(5'h13):(1'h0)] wire511;
  input wire signed [(3'h7):(1'h0)] wire510;
  input wire [(3'h7):(1'h0)] wire509;
  input wire signed [(2'h2):(1'h0)] wire508;
  reg [(2'h3):(1'h0)] reg542 = (1'h0);
  reg [(4'hb):(1'h0)] reg541 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg540 = (1'h0);
  reg [(5'h14):(1'h0)] reg539 = (1'h0);
  reg [(2'h2):(1'h0)] reg538 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar537 = (1'h0);
  reg [(3'h5):(1'h0)] reg536 = (1'h0);
  reg [(5'h14):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg534 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg533 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg532 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg531 = (1'h0);
  reg [(3'h7):(1'h0)] reg530 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg529 = (1'h0);
  reg [(4'ha):(1'h0)] forvar528 = (1'h0);
  reg [(3'h5):(1'h0)] forvar527 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg526 = (1'h0);
  reg [(3'h7):(1'h0)] reg525 = (1'h0);
  reg [(5'h15):(1'h0)] reg524 = (1'h0);
  reg [(4'hf):(1'h0)] reg523 = (1'h0);
  reg [(4'hf):(1'h0)] reg522 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg521 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg520 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg519 = (1'h0);
  reg [(5'h11):(1'h0)] reg518 = (1'h0);
  reg [(5'h14):(1'h0)] reg517 = (1'h0);
  reg [(5'h11):(1'h0)] reg516 = (1'h0);
  reg [(4'hc):(1'h0)] reg515 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg514 = (1'h0);
  reg [(2'h2):(1'h0)] reg513 = (1'h0);
  assign y = {reg542,
                 reg541,
                 reg540,
                 reg539,
                 reg538,
                 forvar537,
                 reg536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 forvar528,
                 forvar527,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 reg517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg513 <= $signed(((+"o") ?
          $unsigned(({wire510, wire512} ?
              $unsigned(wire508) : wire511)) : (wire512[(1'h0):(1'h0)] ?
              $unsigned("m") : {((8'ha9) << (8'ha1))})));
      reg514 = $unsigned($unsigned((^wire508[(1'h1):(1'h0)])));
      reg515 <= wire511;
      reg516 <= reg513;
      reg517 <= (wire511[(5'h12):(4'hd)] >>> ($unsigned($unsigned((|reg515))) | wire509));
    end
  always
    @(posedge clk) begin
      reg518 <= reg516;
      reg519 <= ((~|$unsigned(((8'hb5) ?
              (reg516 ? (8'hb0) : reg517) : reg516[(4'he):(4'he)]))) ?
          $signed((wire509[(3'h4):(1'h1)] ^ $unsigned((!reg516)))) : (~&($signed({wire511,
                  wire512}) ?
              (wire510[(3'h6):(3'h4)] > $signed(wire512)) : reg513)));
    end
  always
    @(posedge clk) begin
      reg520 <= "hvo";
    end
  always
    @(posedge clk) begin
      reg521 <= {{$unsigned(($unsigned(reg517) ? "UEc6vfgSFQntOmwX6c" : "qt"))},
          (({(reg513 <= (8'hb1)), (!reg516)} ?
                  wire510[(2'h2):(1'h1)] : $unsigned("L5cywXhv2Qu")) ?
              $signed($signed((wire510 ? wire512 : reg516))) : (&wire512))};
      reg522 <= "4RBA8zrTVC9";
      reg523 = {{((-((7'h40) ? wire512 : wire512)) ?
                  $unsigned($signed(wire512)) : (~"ZXAmR7ryxGlIMKpq")),
              ((8'hb9) ? wire508[(2'h2):(1'h0)] : "NbNMYOUEb")},
          {$unsigned($unsigned($unsigned(wire508))),
              (((reg520 * wire509) && ((8'hb7) ? wire510 : reg513)) ?
                  ((reg521 <<< wire508) == "WUxcNcvuUd4TbHk6") : "rqth6xgGt9zZ3xPzh")}};
    end
  always
    @(posedge clk) begin
      reg524 <= (!"Vb1X69C");
      reg525 <= $unsigned($unsigned((8'ha7)));
    end
  always
    @(posedge clk) begin
      reg526 <= $unsigned($unsigned($signed((wire510 >>> (|reg519)))));
      for (forvar527 = (1'h0); (forvar527 < (3'h4)); forvar527 = (forvar527 + (1'h1)))
        begin
          for (forvar528 = (1'h0); (forvar528 < (1'h1)); forvar528 = (forvar528 + (1'h1)))
            begin
              reg529 <= ($signed(reg523[(4'he):(4'hd)]) ~^ "");
              reg530 <= {"xLXhfeIxSJ7Qr54WGp"};
              reg531 = (reg523 ?
                  ($signed($signed(reg514[(4'hc):(3'h7)])) ?
                      $signed(($signed(wire508) == $unsigned(reg526))) : reg530) : $signed(((~|$signed(reg520)) | $signed({reg518,
                      reg526}))));
            end
        end
      reg532 = $signed($unsigned(reg519[(3'h6):(3'h4)]));
      reg533 = {(!(("q8ZcNzAUKxck" ?
                  (wire511 ~^ reg515) : reg519[(1'h1):(1'h1)]) ?
              (~^wire511) : $unsigned(reg519[(2'h3):(1'h0)])))};
      reg534 <= (&($signed("2NY8S9XO5FN2D") ?
          (reg519 ?
              {{reg525}} : reg514[(3'h5):(2'h3)]) : reg521[(5'h16):(5'h15)]));
    end
  always
    @(posedge clk) begin
      reg535 = (7'h44);
      reg536 <= (|$unsigned(reg533[(3'h4):(1'h0)]));
      for (forvar537 = (1'h0); (forvar537 < (3'h4)); forvar537 = (forvar537 + (1'h1)))
        begin
          reg538 <= $signed(reg517);
          reg539 <= $unsigned((8'hbc));
        end
      reg540 = ($unsigned(wire508) <<< reg520[(3'h5):(2'h3)]);
    end
  always
    @(posedge clk) begin
      reg541 <= {$signed("rfDZ")};
      reg542 = "8MwZb2zm4NvfUevRx";
    end
endmodule