(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param1883 = (+(({((8'ha6) ^~ (8'had))} ? (((8'h9f) ^ (8'hb7)) + (~^(7'h41))) : ({(8'hb4)} & {(8'haa)})) ? (({(8'h9e), (7'h44)} == ((8'hb6) & (8'hac))) <= (8'hbc)) : (~|(((8'hb6) ? (8'hbf) : (8'hb2)) * (8'hb1))))) )
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h317):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire0;
  input wire signed [(5'h15):(1'h0)] wire1;
  input wire [(5'h12):(1'h0)] wire2;
  input wire signed [(5'h15):(1'h0)] wire3;
  input wire [(5'h15):(1'h0)] wire4;
  wire signed [(3'h7):(1'h0)] wire1882;
  reg [(4'hf):(1'h0)] reg1881 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1880 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1879 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1878 = (1'h0);
  reg [(3'h6):(1'h0)] reg1877 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1876 = (1'h0);
  reg [(4'ha):(1'h0)] reg1875 = (1'h0);
  reg [(5'h11):(1'h0)] reg1874 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1873 = (1'h0);
  reg [(3'h6):(1'h0)] reg1872 = (1'h0);
  reg [(3'h5):(1'h0)] reg1871 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1870 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1869 = (1'h0);
  reg [(2'h2):(1'h0)] reg1868 = (1'h0);
  reg [(4'he):(1'h0)] reg1867 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1866 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1865 = (1'h0);
  reg [(5'h15):(1'h0)] reg1864 = (1'h0);
  reg [(3'h5):(1'h0)] reg1863 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1862 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1861 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1860 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1859 = (1'h0);
  reg [(4'hf):(1'h0)] reg1858 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1857;
  wire signed [(3'h4):(1'h0)] wire1856;
  reg signed [(4'hf):(1'h0)] reg1855 = (1'h0);
  reg [(5'h15):(1'h0)] reg1854 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1853 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1852 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1851 = (1'h0);
  reg [(3'h6):(1'h0)] reg1850 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1849 = (1'h0);
  reg [(3'h5):(1'h0)] reg1848 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1847 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1846 = (1'h0);
  reg [(3'h6):(1'h0)] reg1845 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1844 = (1'h0);
  reg [(5'h10):(1'h0)] reg1843 = (1'h0);
  reg [(3'h5):(1'h0)] reg1842 = (1'h0);
  wire [(4'hb):(1'h0)] wire1841;
  wire signed [(2'h3):(1'h0)] wire1840;
  wire signed [(4'hc):(1'h0)] wire485;
  wire signed [(5'h14):(1'h0)] wire43;
  wire signed [(5'h11):(1'h0)] wire41;
  wire signed [(3'h7):(1'h0)] wire487;
  reg [(3'h6):(1'h0)] reg488 = (1'h0);
  wire [(3'h7):(1'h0)] wire489;
  wire [(4'hf):(1'h0)] wire490;
  reg [(4'hd):(1'h0)] reg491 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg492 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg493 = (1'h0);
  reg [(5'h13):(1'h0)] reg494 = (1'h0);
  reg [(4'he):(1'h0)] reg495 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg496 = (1'h0);
  reg [(4'hd):(1'h0)] reg497 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg498 = (1'h0);
  reg [(3'h6):(1'h0)] reg499 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg500 = (1'h0);
  reg [(5'h10):(1'h0)] reg501 = (1'h0);
  wire signed [(4'he):(1'h0)] wire502;
  wire signed [(5'h12):(1'h0)] wire503;
  reg signed [(3'h6):(1'h0)] reg504 = (1'h0);
  reg [(2'h2):(1'h0)] reg505 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg506 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg507 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg508 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg510 = (1'h0);
  reg signed [(4'he):(1'h0)] reg511 = (1'h0);
  reg [(4'h9):(1'h0)] reg512 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire513;
  wire [(5'h13):(1'h0)] wire1838;
  assign y = {wire1882,
                 reg1881,
                 reg1880,
                 reg1879,
                 reg1878,
                 reg1877,
                 reg1876,
                 reg1875,
                 reg1874,
                 reg1873,
                 reg1872,
                 reg1871,
                 reg1870,
                 reg1869,
                 reg1868,
                 reg1867,
                 reg1866,
                 reg1865,
                 reg1864,
                 reg1863,
                 reg1862,
                 reg1861,
                 reg1860,
                 reg1859,
                 reg1858,
                 wire1857,
                 wire1856,
                 reg1855,
                 reg1854,
                 reg1853,
                 reg1852,
                 reg1851,
                 reg1850,
                 reg1849,
                 reg1848,
                 reg1847,
                 reg1846,
                 reg1845,
                 reg1844,
                 reg1843,
                 reg1842,
                 wire1841,
                 wire1840,
                 wire485,
                 wire43,
                 wire41,
                 wire487,
                 reg488,
                 wire489,
                 wire490,
                 reg491,
                 reg492,
                 reg493,
                 reg494,
                 reg495,
                 reg496,
                 reg497,
                 reg498,
                 reg499,
                 reg500,
                 reg501,
                 wire502,
                 wire503,
                 reg504,
                 reg505,
                 reg506,
                 reg507,
                 reg508,
                 reg509,
                 reg510,
                 reg511,
                 reg512,
                 wire513,
                 wire1838,
                 (1'h0)};
  module5 modinst42 (.wire8(wire4), .wire10(wire0), .wire9(wire2), .wire6(wire1), .y(wire41), .wire7(wire3), .clk(clk));
  assign wire43 = wire4;
  module44 modinst486 (.y(wire485), .wire47(wire0), .clk(clk), .wire48(wire43), .wire45(wire41), .wire49(wire4), .wire46(wire2));
  assign wire487 = ((wire1 ?
                       wire43 : (+(^~$unsigned(wire2)))) != $signed({((wire485 * wire2) <= (8'hbd))}));
  always
    @(posedge clk) begin
      reg488 <= ($unsigned((&($unsigned((8'ha9)) >> $signed(wire487)))) ^~ wire41);
    end
  assign wire489 = ((~|{$unsigned(wire487)}) >> ($unsigned(wire2[(4'h8):(1'h1)]) ?
                       ({(^(8'hb5))} ?
                           wire487[(2'h2):(2'h2)] : $unsigned((wire41 ?
                               (8'h9d) : wire4))) : wire3));
  assign wire490 = $signed(wire487[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      if (((8'hb3) ?
          {(!$signed($unsigned(wire487)))} : (wire0[(2'h2):(1'h0)] || $unsigned($unsigned(wire4)))))
        begin
          if (($unsigned((&(^~$unsigned(wire490)))) ?
              wire1 : ((8'hb7) < wire3)))
            begin
              reg491 <= $unsigned(wire490[(4'h9):(2'h3)]);
              reg492 <= $signed($signed(((~^(wire487 ? wire2 : wire2)) ?
                  ((wire1 ?
                      wire2 : wire489) - (!wire490)) : ((|wire2) == $unsigned(wire485)))));
              reg493 <= $signed(wire4);
              reg494 <= ((wire489 ?
                  (+((wire3 ? reg491 : wire4) ?
                      (wire43 ^ reg493) : (-wire489))) : wire0[(4'hb):(2'h3)]) + wire4);
            end
          else
            begin
              reg491 <= ((wire0[(5'h15):(3'h6)] ? $signed(reg492) : {wire1}) ?
                  ({$unsigned((~&wire485))} ^~ {(wire485[(3'h7):(3'h5)] && (reg494 >= wire43)),
                      $unsigned((reg488 ? wire490 : wire485))}) : (8'haa));
              reg492 <= ((8'hb9) ?
                  (8'hbb) : $signed(($unsigned((wire487 ? wire4 : wire4)) ?
                      ((&wire490) <<< (reg494 ? wire1 : wire487)) : {{(8'hb6)},
                          reg492[(1'h0):(1'h0)]})));
              reg493 <= $unsigned((+wire3));
            end
        end
      else
        begin
          if ($unsigned(wire3[(2'h2):(1'h1)]))
            begin
              reg491 <= {(($signed((wire0 ? wire43 : wire43)) ?
                          (wire2 == $unsigned(wire490)) : $signed((wire490 != wire487))) ?
                      ((~&(wire485 ? wire3 : reg488)) ?
                          (+(wire4 ?
                              wire4 : wire1)) : wire4) : $unsigned(reg492[(1'h1):(1'h0)]))};
              reg492 <= {((^~wire487[(1'h1):(1'h0)]) && ((^~$unsigned(wire2)) ?
                      reg488[(3'h6):(1'h1)] : $unsigned(wire0))),
                  (8'ha3)};
              reg493 <= wire487;
            end
          else
            begin
              reg491 <= ($signed($unsigned((^{wire487}))) ?
                  reg494[(4'h9):(2'h3)] : $unsigned(($signed($unsigned(reg488)) | (+(wire3 ?
                      wire1 : (8'ha3))))));
              reg492 <= wire2;
              reg493 <= (~^($signed(($unsigned(wire489) ?
                      $signed(reg491) : (~&(8'hbb)))) ?
                  wire41[(4'hd):(1'h1)] : $signed((~(wire490 <= wire0)))));
            end
          if (({($unsigned(wire3) ?
                      wire485[(4'h9):(1'h0)] : $unsigned(((8'hb9) == reg491)))} ?
              $signed(wire3) : $unsigned($unsigned((wire43 || wire3)))))
            begin
              reg494 <= $unsigned(($unsigned({(8'hbd), {reg494}}) ?
                  wire4 : (wire490[(4'ha):(4'h9)] >> wire2)));
            end
          else
            begin
              reg494 <= $signed(((wire3[(1'h1):(1'h1)] ^ $unsigned((&wire3))) ?
                  (~|$signed((reg488 | reg493))) : ($unsigned($signed(wire41)) ?
                      {wire0, {wire1, wire43}} : wire4[(1'h1):(1'h0)])));
              reg495 <= ({$signed(wire41[(5'h11):(2'h3)]),
                  (reg494 ?
                      $unsigned((wire489 ?
                          reg491 : wire43)) : $signed($unsigned(wire485)))} > (~^$signed($signed($signed(wire0)))));
              reg496 <= (8'h9d);
              reg497 <= (^$unsigned(reg494));
              reg498 <= ($unsigned((~^{(wire4 ?
                      reg488 : wire1)})) || ((~^($signed(wire3) & {wire3,
                      wire43})) ?
                  wire489 : $signed($unsigned(wire3[(5'h11):(2'h2)]))));
            end
          reg499 <= $unsigned($unsigned((($signed((7'h42)) || (|(8'ha3))) > ((wire41 ?
                  reg496 : reg493) ?
              (wire485 & reg491) : $signed(reg494)))));
        end
      reg500 <= $signed(reg499[(2'h2):(1'h1)]);
      reg501 <= $signed($signed($signed(($signed(reg495) ?
          {reg488, wire0} : wire41))));
    end
  assign wire502 = wire490;
  assign wire503 = wire485[(3'h4):(3'h4)];
  always
    @(posedge clk) begin
      if ($signed($unsigned(($unsigned($signed(reg497)) & (~^$unsigned(reg498))))))
        begin
          reg504 <= $unsigned(((8'haa) && {($signed(reg492) ?
                  wire43 : (|reg498))}));
          if ($unsigned($signed($signed((wire487[(2'h3):(2'h3)] ^~ (wire43 - reg493))))))
            begin
              reg505 <= {(~&((reg488 ~^ (~^reg496)) ?
                      ((+wire41) ?
                          (wire0 && reg500) : (^~reg497)) : $signed($signed(wire487)))),
                  reg491[(3'h6):(2'h3)]};
              reg506 <= (^~wire2);
              reg507 <= (+((!reg488[(2'h3):(1'h0)]) >> ((wire2 - {reg499}) << ($signed(reg494) ?
                  wire489[(3'h6):(2'h2)] : (reg488 ? wire1 : (8'had))))));
              reg508 <= $unsigned((~^reg505));
            end
          else
            begin
              reg505 <= $unsigned(reg501[(3'h4):(1'h1)]);
              reg506 <= reg495;
              reg507 <= (reg500 <= reg498);
            end
          reg509 <= (8'h9d);
          reg510 <= (((reg500 != wire489[(3'h7):(1'h0)]) ~^ wire4[(2'h3):(2'h3)]) || (($unsigned($signed(reg488)) ^ ((wire502 > reg507) ?
              $unsigned(wire489) : (~^wire2))) & $unsigned(reg508[(2'h3):(1'h0)])));
          reg511 <= (reg508[(2'h3):(2'h2)] >>> {reg507[(1'h0):(1'h0)], reg494});
        end
      else
        begin
          reg504 <= ($unsigned((reg509 ?
                  $signed(wire41[(4'he):(4'h9)]) : (8'hb7))) ?
              reg510 : reg499);
        end
      reg512 <= $signed($signed($signed(reg498)));
    end
  assign wire513 = reg512[(1'h0):(1'h0)];
  module514 modinst1839 (wire1838, clk, wire503, reg510, reg492, reg501, reg498);
  assign wire1840 = {wire513,
                        (~|{reg499, {((8'hb3) ? reg496 : wire503), {reg495}}})};
  assign wire1841 = $unsigned($signed(wire487[(3'h7):(3'h7)]));
  always
    @(posedge clk) begin
      reg1842 <= ((((wire485[(1'h1):(1'h0)] ?
                      wire0 : (reg504 ? reg494 : wire43)) ?
                  reg507[(2'h2):(2'h2)] : $signed($unsigned(reg505))) ?
              (reg501[(4'h8):(1'h0)] >> reg501) : $signed(wire513)) ?
          $signed((+{$signed(reg512)})) : $unsigned({$unsigned(((8'h9f) >>> wire503)),
              ((wire3 ? (8'h9e) : wire41) ? (~|reg493) : $unsigned((8'hac)))}));
      if ((^~$signed(wire0[(5'h10):(5'h10)])))
        begin
          reg1843 <= $signed((&($signed($signed(reg511)) == ((reg504 ^ wire1841) << reg498[(4'ha):(3'h5)]))));
          if (reg1842[(2'h3):(2'h3)])
            begin
              reg1844 <= wire1[(1'h1):(1'h1)];
              reg1845 <= ($signed((&(((8'hac) ? wire1 : wire489) ?
                      $unsigned(wire487) : reg498))) ?
                  $signed($signed(reg509[(4'ha):(2'h2)])) : wire513[(2'h2):(1'h1)]);
              reg1846 <= (|reg511);
              reg1847 <= wire1838[(5'h11):(2'h2)];
              reg1848 <= (reg509[(4'hd):(4'h9)] << $signed($unsigned(reg488)));
            end
          else
            begin
              reg1844 <= ($signed({(8'hb9),
                      ((wire1838 ~^ reg1846) ^ $unsigned(reg512))}) ?
                  $unsigned(reg509) : (~&$unsigned($signed($unsigned(reg1843)))));
              reg1845 <= $signed((&(8'hae)));
            end
          if ($unsigned(($unsigned($signed((wire490 ?
              reg511 : (8'h9e)))) != (({reg491} ?
              reg500[(1'h0):(1'h0)] : (reg512 + reg1842)) ~^ (^(8'ha2))))))
            begin
              reg1849 <= {reg1845};
              reg1850 <= (8'hb6);
              reg1851 <= ((+(~&((~reg1842) ?
                  (+wire503) : (^(7'h44))))) ^~ ($signed((^~$unsigned(reg488))) >>> $unsigned($unsigned($unsigned((7'h42))))));
            end
          else
            begin
              reg1849 <= ($unsigned((+reg492)) ?
                  (wire2 | (|(reg1847 ?
                      (reg501 && reg512) : reg507))) : (^$unsigned((~&(wire1 ?
                      reg511 : wire41)))));
              reg1850 <= ($signed((reg507 ? {$unsigned(wire489)} : reg1843)) ?
                  (^($unsigned($signed((8'h9f))) ?
                      wire43[(4'h8):(3'h5)] : reg496)) : wire2[(5'h12):(4'hd)]);
              reg1851 <= (^(reg491 == (-$signed((wire3 == reg504)))));
              reg1852 <= $unsigned(reg496[(4'hd):(4'ha)]);
            end
          reg1853 <= $unsigned(wire485[(4'h8):(4'h8)]);
        end
      else
        begin
          if (reg505)
            begin
              reg1843 <= $unsigned(reg500[(2'h3):(1'h1)]);
              reg1844 <= $signed(($signed(wire1838) <<< $unsigned(($signed(wire2) >= $signed(reg1853)))));
              reg1845 <= reg492;
              reg1846 <= (~^(((wire1841 && (~(8'ha5))) >> ($unsigned(wire513) ?
                  reg1850[(2'h3):(1'h1)] : $unsigned(reg1844))) + (+(^~wire1))));
              reg1847 <= $unsigned(wire490);
            end
          else
            begin
              reg1843 <= (wire1840 >= {(~|($signed((7'h43)) <= $unsigned(reg1853)))});
              reg1844 <= reg1853;
              reg1845 <= $unsigned($unsigned({((~reg1845) ?
                      (reg494 ? reg1848 : wire513) : reg504[(3'h4):(3'h4)]),
                  (wire502[(3'h5):(3'h5)] >= reg1851[(2'h3):(2'h2)])}));
              reg1846 <= (((~^(((8'ha4) * wire502) ?
                          (reg498 <<< reg500) : (8'hbe))) ?
                      wire4 : (&((reg508 ? wire485 : reg1842) ?
                          {reg500, wire1841} : $signed(wire487)))) ?
                  reg496 : ({reg506[(3'h7):(3'h5)]} ?
                      (reg1853[(2'h3):(1'h1)] ?
                          $unsigned($signed(wire487)) : (wire0 >>> wire502)) : (($signed(reg1852) || (reg499 == wire4)) ?
                          $signed((+(8'hb4))) : (~&reg497[(4'h9):(3'h6)]))));
              reg1847 <= $signed($signed($signed($signed(reg497))));
            end
          reg1848 <= (+$signed((^~(^~reg1846[(1'h0):(1'h0)]))));
          reg1849 <= ((($signed((reg495 ? wire489 : reg509)) <<< ((-wire485) ?
                  $signed(reg1849) : (8'hb9))) <= (reg1846 >>> $signed(reg512[(2'h3):(1'h0)]))) ?
              (wire4[(3'h7):(1'h0)] & $signed((wire4 ?
                  {reg501,
                      reg1850} : (8'ha0)))) : $unsigned((((wire4 <<< wire1838) * (-wire43)) >= reg1846[(1'h0):(1'h0)])));
          reg1850 <= (~^$unsigned((wire485 ?
              reg496 : $signed($signed(reg509)))));
        end
      reg1854 <= reg498[(2'h2):(1'h1)];
      reg1855 <= $unsigned(reg1847[(2'h2):(2'h2)]);
    end
  assign wire1856 = {$unsigned($unsigned($unsigned((|reg1847))))};
  assign wire1857 = $signed((-wire1838[(4'ha):(1'h0)]));
  always
    @(posedge clk) begin
      reg1858 <= reg500[(2'h2):(2'h2)];
      reg1859 <= $unsigned({({wire2[(2'h3):(2'h2)]} > ((|reg1850) > (reg491 ?
              reg499 : reg1854))),
          wire513[(2'h2):(1'h0)]});
      if ($signed((~{reg1851[(3'h5):(1'h0)]})))
        begin
          reg1860 <= {($signed(reg491[(2'h2):(1'h1)]) ~^ (~&$signed((~|reg1848))))};
          reg1861 <= ((|(8'ha5)) ?
              ($unsigned(reg1855[(4'he):(4'hb)]) ?
                  (8'h9c) : (&(reg1848 ?
                      {reg501,
                          wire1838} : (reg493 != wire1856)))) : {(-(~^$signed(reg1854))),
                  ($signed((reg1854 ~^ wire1856)) != (&(&wire2)))});
          if ($unsigned({reg500,
              {$signed(wire43[(1'h1):(1'h1)]), $unsigned({wire3, (8'h9e)})}}))
            begin
              reg1862 <= ((wire502 <<< $signed($unsigned($unsigned(wire1838)))) ?
                  ($unsigned($signed((wire513 | reg1860))) ?
                      $unsigned(reg488) : $unsigned($signed(reg1853[(3'h5):(2'h3)]))) : (^~(^$unsigned((reg1853 <= (8'h9e))))));
              reg1863 <= wire1841[(4'h8):(3'h4)];
            end
          else
            begin
              reg1862 <= {(+reg1860),
                  (~({(reg1847 ~^ reg1844)} == $signed(wire2)))};
              reg1863 <= (~&$unsigned(((8'ha6) ?
                  reg1861 : (-(reg493 ? wire4 : reg510)))));
              reg1864 <= {reg501[(4'ha):(4'h9)]};
              reg1865 <= ((-wire1840) != $unsigned(((reg499[(3'h5):(1'h1)] ?
                      (~reg1847) : (&reg1852)) ?
                  $unsigned((reg512 >>> reg501)) : (-(~reg1852)))));
            end
          reg1866 <= reg1847[(2'h2):(2'h2)];
        end
      else
        begin
          if ((^~(8'haa)))
            begin
              reg1860 <= reg1847;
              reg1861 <= reg1855[(4'h9):(3'h7)];
              reg1862 <= $unsigned((&{$unsigned((reg1851 << wire513)),
                  {$unsigned(reg1860)}}));
              reg1863 <= $unsigned($unsigned((reg1854 != $signed((^reg495)))));
              reg1864 <= $unsigned(wire1841);
            end
          else
            begin
              reg1860 <= (((|reg497) >>> ((reg1865 >> (wire43 <<< (8'h9e))) == (|(~(7'h43))))) ?
                  (($unsigned((wire41 ?
                      reg1850 : reg1851)) ^~ $unsigned(reg504)) ^~ (!reg1862)) : ($signed({wire503,
                      (reg1843 ? (8'hbf) : reg510)}) | (~^$signed({reg499}))));
            end
          if ((8'hb5))
            begin
              reg1865 <= $unsigned((^$signed($unsigned(reg504[(2'h2):(1'h1)]))));
              reg1866 <= {$unsigned($signed($signed({wire0})))};
              reg1867 <= $signed($unsigned($signed($unsigned(reg509))));
            end
          else
            begin
              reg1865 <= $unsigned(($unsigned($signed((^~reg512))) ?
                  ($signed((reg494 >> reg496)) & ($unsigned((8'ha5)) ?
                      (&reg509) : (reg492 ^ reg1866))) : (wire3[(4'hb):(4'ha)] ?
                      $signed($unsigned(wire1856)) : $unsigned($signed(reg488)))));
              reg1866 <= $signed($signed(((8'ha9) ?
                  (reg511[(2'h3):(1'h0)] ?
                      reg492 : (wire485 ?
                          (8'h9c) : reg1862)) : $signed(reg492))));
              reg1867 <= (reg505 ?
                  reg1854 : ((~|$unsigned(reg1855[(3'h7):(3'h5)])) | (($signed(reg1843) + wire3[(3'h6):(2'h2)]) ?
                      (-(~reg1842)) : {reg1862[(3'h4):(1'h0)],
                          reg1859[(3'h7):(3'h4)]})));
              reg1868 <= wire1838;
              reg1869 <= (reg497 ?
                  ($unsigned((~$unsigned(reg511))) ?
                      ($signed({reg1845, reg1850}) ?
                          $signed(wire41[(3'h5):(2'h2)]) : $unsigned(reg1863)) : $unsigned($unsigned($signed((7'h42))))) : $unsigned($signed($unsigned((reg491 == reg1867)))));
            end
          reg1870 <= {((!wire1838) ?
                  ($unsigned((reg1865 ? reg1867 : reg512)) ?
                      reg511[(1'h1):(1'h1)] : (|$unsigned(reg493))) : ($signed((8'hb1)) ?
                      (~|(8'hb9)) : reg508))};
        end
      if (((8'h9d) ?
          $unsigned(reg1855[(4'hf):(4'he)]) : ((($unsigned(reg1853) ?
                  {reg498} : reg1865[(3'h5):(1'h1)]) ?
              (7'h41) : reg500) & (^($unsigned(reg496) == $signed(reg1863))))))
        begin
          reg1871 <= (reg1845 ?
              wire487 : $unsigned(($signed({reg1859, reg1850}) ?
                  ($signed((8'hab)) == {reg1853}) : (-reg1861[(4'hc):(4'hc)]))));
          if (reg1860[(3'h7):(1'h1)])
            begin
              reg1872 <= $unsigned((!reg1869));
              reg1873 <= ({(8'ha9),
                  $signed($signed((+reg497)))} * (reg1871[(1'h1):(1'h0)] ?
                  (reg501[(1'h1):(1'h1)] ?
                      reg1858 : wire503[(1'h0):(1'h0)]) : (|$unsigned((reg1865 ?
                      wire513 : reg1860)))));
              reg1874 <= (-(-(+($signed(reg1858) == $unsigned(reg496)))));
              reg1875 <= reg1868;
            end
          else
            begin
              reg1872 <= ($signed(reg507[(1'h1):(1'h0)]) && (-(((reg508 ?
                  wire1 : reg1864) || $signed(wire1856)) ~^ $unsigned(wire503[(4'h9):(2'h3)]))));
            end
          reg1876 <= reg508[(1'h1):(1'h0)];
          if (reg1845[(3'h4):(1'h1)])
            begin
              reg1877 <= ((wire489[(2'h3):(1'h1)] ?
                  ((reg496[(4'h9):(2'h2)] ?
                      (reg1844 < reg1871) : (reg1842 >> reg492)) | reg496[(3'h5):(3'h4)]) : $unsigned($unsigned(reg1858))) > (({(8'hb4)} ?
                  reg1844 : (8'ha1)) ~^ {(8'hbb), reg1862[(4'hb):(4'ha)]}));
              reg1878 <= (~&(&reg501));
              reg1879 <= $signed(reg1855[(1'h0):(1'h0)]);
              reg1880 <= ($signed((|$unsigned((wire43 ?
                  reg1850 : reg1874)))) * {$unsigned((!reg1872))});
            end
          else
            begin
              reg1877 <= ((((~&(8'hb7)) ?
                  $unsigned((reg507 ~^ wire485)) : reg492) ^ (~&(|{wire490,
                  reg508}))) || {(reg1849 ?
                      $signed((-(8'hbb))) : (-$signed(reg509))),
                  $signed((^{(8'hb5)}))});
            end
          reg1881 <= ($signed((({reg1863} | $signed(reg1860)) ?
                  (&reg1875) : (8'hac))) ?
              reg1865 : (|(~wire1840[(2'h2):(2'h2)])));
        end
      else
        begin
          reg1871 <= $signed($signed(reg1866));
          if (wire1856)
            begin
              reg1872 <= ((~reg496) ~^ (reg498 >= (!((~|reg1858) ?
                  wire1838[(5'h11):(3'h6)] : (~|wire489)))));
              reg1873 <= reg493[(4'hb):(2'h3)];
            end
          else
            begin
              reg1872 <= {reg1855};
              reg1873 <= {(8'hb5),
                  {(^({reg491} || wire2[(4'hb):(4'h8)])),
                      $unsigned((reg1867 ?
                          $unsigned((8'hbc)) : reg500[(2'h2):(1'h0)]))}};
            end
          reg1874 <= ($signed((~(^~reg1876[(1'h1):(1'h0)]))) <= reg1859[(4'hc):(2'h2)]);
        end
    end
  assign wire1882 = (reg500[(1'h1):(1'h1)] <= (($unsigned((8'ha1)) > $signed((reg1871 ?
                            reg488 : reg1845))) ?
                        {{(+(8'ha8))}, reg1850} : $unsigned(wire485)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module514  (y, clk, wire515, wire516, wire517, wire518, wire519);
  output wire [(32'h1e9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire515;
  input wire [(5'h10):(1'h0)] wire516;
  input wire [(4'hc):(1'h0)] wire517;
  input wire signed [(5'h10):(1'h0)] wire518;
  input wire [(4'h8):(1'h0)] wire519;
  wire [(5'h15):(1'h0)] wire1836;
  wire [(3'h4):(1'h0)] wire520;
  reg [(4'ha):(1'h0)] reg521 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg522 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg523 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg524 = (1'h0);
  reg [(3'h4):(1'h0)] reg525 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg526 = (1'h0);
  reg [(2'h3):(1'h0)] reg527 = (1'h0);
  reg [(3'h6):(1'h0)] reg528 = (1'h0);
  reg [(5'h13):(1'h0)] reg529 = (1'h0);
  reg [(4'ha):(1'h0)] reg530 = (1'h0);
  reg [(5'h15):(1'h0)] reg531 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg532 = (1'h0);
  wire [(4'hf):(1'h0)] wire533;
  wire signed [(5'h15):(1'h0)] wire534;
  reg signed [(3'h6):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg536 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg537 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire538;
  wire signed [(5'h13):(1'h0)] wire539;
  wire [(4'hf):(1'h0)] wire540;
  wire signed [(5'h12):(1'h0)] wire541;
  wire signed [(4'h8):(1'h0)] wire542;
  wire [(5'h14):(1'h0)] wire543;
  wire signed [(4'ha):(1'h0)] wire544;
  reg signed [(4'hd):(1'h0)] reg545 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg546 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg547 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg548 = (1'h0);
  reg [(2'h3):(1'h0)] reg549 = (1'h0);
  reg [(3'h4):(1'h0)] reg550 = (1'h0);
  reg [(3'h7):(1'h0)] reg551 = (1'h0);
  reg [(4'h8):(1'h0)] reg552 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire553;
  wire [(4'hd):(1'h0)] wire554;
  wire signed [(5'h13):(1'h0)] wire1834;
  assign y = {wire1836,
                 wire520,
                 reg521,
                 reg522,
                 reg523,
                 reg524,
                 reg525,
                 reg526,
                 reg527,
                 reg528,
                 reg529,
                 reg530,
                 reg531,
                 reg532,
                 wire533,
                 wire534,
                 reg535,
                 reg536,
                 reg537,
                 wire538,
                 wire539,
                 wire540,
                 wire541,
                 wire542,
                 wire543,
                 wire544,
                 reg545,
                 reg546,
                 reg547,
                 reg548,
                 reg549,
                 reg550,
                 reg551,
                 reg552,
                 wire553,
                 wire554,
                 wire1834,
                 (1'h0)};
  assign wire520 = $unsigned(($signed((wire516[(4'h9):(2'h2)] << (wire519 ?
                       wire518 : wire517))) >= wire517));
  always
    @(posedge clk) begin
      reg521 <= $unsigned({$signed(wire517),
          ((&((8'hb4) < wire516)) >= wire516)});
      reg522 <= ((+{$signed(((8'hbc) ? wire519 : wire516)),
          (8'ha4)}) || wire516[(2'h2):(1'h0)]);
      if ((8'haa))
        begin
          reg523 <= wire520[(3'h4):(2'h2)];
          reg524 <= (8'h9d);
          reg525 <= {(8'ha7),
              $signed(((wire520 ? $unsigned(reg521) : {wire520}) ?
                  (((8'haa) <= (8'hbe)) > (~&(8'hb8))) : wire520))};
          reg526 <= reg525;
          reg527 <= (~&(&(8'h9c)));
        end
      else
        begin
          reg523 <= $unsigned((~|reg525[(1'h1):(1'h0)]));
          reg524 <= reg522[(3'h6):(3'h4)];
          reg525 <= wire519;
          if ($unsigned((+{$signed(reg525)})))
            begin
              reg526 <= {wire520[(2'h2):(1'h1)]};
              reg527 <= $unsigned($unsigned(((&$unsigned(reg525)) >= ((wire517 ?
                  wire519 : (7'h43)) ^~ (+wire518)))));
            end
          else
            begin
              reg526 <= ($signed(wire518[(1'h1):(1'h1)]) >> reg523[(5'h10):(2'h3)]);
              reg527 <= $unsigned(wire516);
              reg528 <= wire515[(4'ha):(2'h3)];
              reg529 <= (wire516[(4'ha):(2'h3)] ?
                  ($unsigned(wire520) ?
                      (((~^reg524) != (wire519 ? wire516 : wire515)) ?
                          reg525 : reg527[(1'h1):(1'h0)]) : {$unsigned($unsigned(reg525)),
                          wire516[(2'h3):(2'h3)]}) : wire518[(1'h1):(1'h1)]);
            end
          reg530 <= $signed($unsigned($unsigned($signed($unsigned((8'hb1))))));
        end
      reg531 <= $signed({$signed({(8'ha6)}), reg527});
      reg532 <= $unsigned((($signed($signed(reg524)) | ((-reg526) ?
              (wire515 * reg522) : wire520[(2'h2):(1'h0)])) ?
          reg527 : reg523));
    end
  assign wire533 = reg521;
  assign wire534 = ((8'hb0) < reg529[(3'h4):(1'h0)]);
  always
    @(posedge clk) begin
      if (reg522)
        begin
          if (wire517[(4'h8):(3'h5)])
            begin
              reg535 <= wire533;
              reg536 <= $signed(reg523[(4'he):(4'hc)]);
            end
          else
            begin
              reg535 <= $signed($unsigned(reg523[(4'h9):(2'h3)]));
            end
          reg537 <= $unsigned((|(reg531 << {(reg531 ? wire518 : wire519),
              wire519})));
        end
      else
        begin
          reg535 <= $signed($unsigned(((~^$unsigned((8'ha9))) < $signed((reg528 <= reg526)))));
        end
    end
  assign wire538 = $unsigned($signed($signed(wire520[(3'h4):(2'h2)])));
  assign wire539 = (~wire517);
  assign wire540 = ($signed((7'h41)) ?
                       (~|(-($signed(reg530) | $signed((8'ha5))))) : $unsigned(reg532[(5'h10):(3'h7)]));
  assign wire541 = $unsigned((($signed((wire518 ? reg532 : reg524)) ?
                           ($signed((8'hb4)) >>> wire539[(2'h3):(2'h2)]) : wire520) ?
                       wire519 : {(wire515[(3'h5):(3'h4)] ?
                               wire517 : $unsigned(reg535)),
                           ((wire518 ? reg529 : wire539) + (-reg527))}));
  assign wire542 = (^~(reg529[(3'h7):(3'h4)] || $signed(reg531[(4'hb):(2'h3)])));
  assign wire543 = (^reg524[(3'h6):(3'h5)]);
  assign wire544 = ($signed((|$unsigned($unsigned(wire539)))) ?
                       $unsigned(((~|reg528) ?
                           reg529 : $signed(reg524[(3'h4):(2'h2)]))) : ($signed(({wire540} ?
                               (~&reg522) : (wire519 ? reg521 : wire516))) ?
                           $unsigned(wire543[(1'h1):(1'h1)]) : (8'hb4)));
  always
    @(posedge clk) begin
      reg545 <= wire541;
      if (((reg522[(4'ha):(4'h9)] != reg537[(1'h1):(1'h0)]) ?
          $signed(((+reg525) ?
              ($unsigned(wire533) && reg535[(1'h0):(1'h0)]) : {(wire517 ?
                      wire539 : wire533)})) : ($unsigned($unsigned((reg535 & reg523))) ?
              $signed($signed($signed(wire517))) : $signed(($signed(reg531) ~^ $unsigned(reg545))))))
        begin
          reg546 <= $signed(reg521[(2'h2):(2'h2)]);
        end
      else
        begin
          if (wire541)
            begin
              reg546 <= ((wire519[(3'h5):(1'h0)] ?
                      (8'hbc) : ((~&$unsigned(reg530)) ?
                          (((8'h9f) ? wire534 : reg521) ?
                              (reg524 ?
                                  reg532 : reg531) : (~|wire541)) : $unsigned($unsigned(wire533)))) ?
                  ($unsigned((|(reg545 ? reg530 : wire516))) ?
                      $signed((+wire542)) : (wire538 >> reg527[(1'h0):(1'h0)])) : (!(8'ha4)));
              reg547 <= wire518[(2'h3):(1'h0)];
            end
          else
            begin
              reg546 <= ({wire542[(1'h0):(1'h0)]} ?
                  ({(reg527[(1'h0):(1'h0)] ? ((8'ha2) && wire539) : wire538)} ?
                      (&((reg532 >>> reg536) ?
                          (^reg537) : wire516[(4'h8):(2'h3)])) : $unsigned((~^reg546))) : $signed(reg536[(3'h6):(3'h4)]));
              reg547 <= (wire543 >>> $signed($unsigned($signed(((7'h43) & wire543)))));
            end
          reg548 <= ((reg545 + wire533) >> reg537);
          reg549 <= (~|(((8'ha6) ?
              $signed(wire517[(4'ha):(3'h7)]) : $signed($signed(wire534))) >>> $signed(wire539[(1'h1):(1'h1)])));
          reg550 <= $signed((!reg547[(2'h3):(1'h0)]));
        end
      reg551 <= (~|wire544[(4'ha):(3'h6)]);
      reg552 <= $signed(reg526);
    end
  assign wire553 = reg545;
  assign wire554 = $unsigned(reg532);
  module555 modinst1835 (wire1834, clk, reg545, wire541, reg531, reg547, wire543);
  module950 modinst1837 (.wire954(wire544), .wire952(wire543), .y(wire1836), .wire953(reg537), .clk(clk), .wire951(wire518));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module44
#( parameter param484 = {((~|({(8'ha8)} & {(8'hb3)})) ^ ((((8'h9c) ? (8'hb0) : (8'hbc)) ? {(8'ha0), (7'h42)} : ((7'h42) ? (8'hb5) : (8'ha3))) ? (((8'hb5) ? (8'hab) : (8'hb5)) < (&(7'h43))) : (((7'h40) - (8'ha5)) ? ((8'hab) > (8'hbd)) : (~^(8'ha8)))))} )
(y, clk, wire45, wire46, wire47, wire48, wire49);
  output wire [(32'h8a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire45;
  input wire signed [(5'h12):(1'h0)] wire46;
  input wire signed [(5'h15):(1'h0)] wire47;
  input wire [(5'h14):(1'h0)] wire48;
  input wire [(5'h15):(1'h0)] wire49;
  wire [(2'h3):(1'h0)] wire483;
  wire [(4'hc):(1'h0)] wire482;
  wire [(3'h7):(1'h0)] wire481;
  wire [(5'h14):(1'h0)] wire480;
  wire [(4'hc):(1'h0)] wire479;
  wire signed [(5'h14):(1'h0)] wire478;
  wire [(5'h15):(1'h0)] wire477;
  wire [(5'h12):(1'h0)] wire476;
  wire signed [(4'ha):(1'h0)] wire475;
  wire [(4'he):(1'h0)] wire473;
  assign y = {wire483,
                 wire482,
                 wire481,
                 wire480,
                 wire479,
                 wire478,
                 wire477,
                 wire476,
                 wire475,
                 wire473,
                 (1'h0)};
  module50 modinst474 (.wire51(wire45), .wire53(wire47), .y(wire473), .clk(clk), .wire54(wire46), .wire55(wire48), .wire52(wire49));
  assign wire475 = $signed({({$unsigned((8'hb9))} && ($signed((7'h42)) ?
                           $signed(wire47) : (^wire47)))});
  assign wire476 = wire475[(1'h1):(1'h0)];
  assign wire477 = (!$signed((7'h41)));
  assign wire478 = wire473[(4'hd):(3'h4)];
  assign wire479 = wire48;
  assign wire480 = wire47[(5'h13):(2'h2)];
  assign wire481 = ((wire476 + ($signed(wire479[(2'h2):(1'h0)]) & (-(wire45 ?
                       wire473 : wire48)))) * $unsigned($unsigned(wire475[(4'h8):(2'h3)])));
  assign wire482 = wire47;
  assign wire483 = (^~(wire479[(4'hc):(3'h5)] & $unsigned((!wire475))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module5  (y, clk, wire10, wire9, wire8, wire7, wire6);
  output wire [(32'h185):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire10;
  input wire [(4'ha):(1'h0)] wire9;
  input wire signed [(4'hd):(1'h0)] wire8;
  input wire signed [(4'he):(1'h0)] wire7;
  input wire [(5'h10):(1'h0)] wire6;
  wire [(5'h11):(1'h0)] wire40;
  reg [(4'he):(1'h0)] reg39 = (1'h0);
  reg [(5'h14):(1'h0)] reg38 = (1'h0);
  reg [(4'ha):(1'h0)] reg37 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg35 = (1'h0);
  reg [(4'hf):(1'h0)] reg34 = (1'h0);
  wire [(4'hf):(1'h0)] wire33;
  wire signed [(5'h14):(1'h0)] wire32;
  wire signed [(4'hd):(1'h0)] wire31;
  wire signed [(4'ha):(1'h0)] wire30;
  wire signed [(4'hd):(1'h0)] wire29;
  reg [(5'h12):(1'h0)] reg28 = (1'h0);
  reg [(4'hb):(1'h0)] reg27 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg26 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg24 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg23 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg22 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg21 = (1'h0);
  reg [(3'h7):(1'h0)] reg20 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg19 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg18 = (1'h0);
  reg [(4'h9):(1'h0)] reg17 = (1'h0);
  reg [(4'hd):(1'h0)] reg16 = (1'h0);
  reg [(5'h12):(1'h0)] reg15 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg14 = (1'h0);
  reg [(3'h4):(1'h0)] reg13 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg12 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire11;
  assign y = {wire40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 wire33,
                 wire32,
                 wire31,
                 wire30,
                 wire29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 wire11,
                 (1'h0)};
  assign wire11 = wire6;
  always
    @(posedge clk) begin
      reg12 <= (wire7[(1'h0):(1'h0)] && wire9);
    end
  always
    @(posedge clk) begin
      if (($signed(wire7[(3'h6):(3'h5)]) & $unsigned($unsigned(reg12[(2'h3):(1'h0)]))))
        begin
          reg13 <= (($unsigned(((wire11 ? wire8 : (8'hbd)) ?
                  wire10[(5'h10):(3'h4)] : (7'h40))) ?
              $unsigned($signed(wire6[(5'h10):(3'h6)])) : (!{((8'ha5) | wire9)})) <<< (wire9 & (~(8'ha0))));
          reg14 <= wire8;
          reg15 <= wire10;
          if ($unsigned($signed(wire7[(4'hd):(3'h4)])))
            begin
              reg16 <= (^~(wire7 || wire11));
              reg17 <= $signed(({(8'ha1), reg16} ?
                  $unsigned((reg14 >> reg16)) : wire10));
              reg18 <= (~^(!(8'ha3)));
              reg19 <= ($unsigned((reg15[(4'hd):(3'h7)] ~^ $signed((~|wire9)))) ^~ (&$signed(reg18)));
              reg20 <= ({wire11,
                  wire10} * $unsigned($unsigned($unsigned((reg15 * wire9)))));
            end
          else
            begin
              reg16 <= ((reg13[(2'h2):(1'h0)] ?
                      wire10 : (+((reg16 || reg19) ?
                          wire9[(1'h0):(1'h0)] : (8'hae)))) ?
                  (reg18 != (~|((^~wire6) ?
                      ((7'h43) >> wire9) : $unsigned(wire6)))) : $unsigned((8'hab)));
              reg17 <= reg16;
              reg18 <= $signed({($signed((wire8 <<< reg16)) >>> ((~|reg12) <= $signed((8'ha9)))),
                  ($signed(reg20) ^ wire9)});
              reg19 <= (((((wire8 <<< reg16) ?
                      reg17 : {reg17, (8'h9d)}) > wire7) * reg14) ?
                  (wire6 ^ $signed(($unsigned(wire8) >= (7'h43)))) : ($signed((^(wire9 ?
                          wire9 : reg20))) ?
                      (wire6[(4'he):(3'h7)] ?
                          {(^~wire11)} : $signed({reg14, reg17})) : {wire6}));
              reg20 <= (wire10 ?
                  ((!wire6[(2'h2):(1'h1)]) + ((reg20[(1'h0):(1'h0)] ?
                          ((8'h9d) ? wire10 : wire6) : wire10) ?
                      wire6 : reg17[(1'h0):(1'h0)])) : ((~|((wire9 ?
                          reg13 : reg18) ^ $unsigned(reg16))) ?
                      (-reg18[(3'h7):(3'h6)]) : (-$unsigned(wire6))));
            end
        end
      else
        begin
          if (((+((^reg16[(2'h2):(1'h1)]) ? {(+reg12)} : $signed((8'hb2)))) ?
              $unsigned({reg19[(2'h2):(2'h2)],
                  {$signed(reg13), $signed(reg20)}}) : {(8'h9f),
                  wire6[(2'h3):(2'h3)]}))
            begin
              reg13 <= {reg13[(2'h2):(2'h2)]};
              reg14 <= (^~reg16[(2'h2):(1'h0)]);
              reg15 <= (+(~|reg19));
              reg16 <= ($unsigned(reg14) ?
                  $signed(wire8) : $unsigned($signed($signed((reg14 ?
                      reg13 : wire9)))));
              reg17 <= $signed($unsigned(reg18[(3'h4):(1'h0)]));
            end
          else
            begin
              reg13 <= reg17[(1'h0):(1'h0)];
            end
          reg18 <= ({(+(&reg19)),
              $signed((~&wire9[(2'h2):(2'h2)]))} && {(((reg17 ? reg17 : reg12) ?
                  ((8'ha5) > wire9) : $signed((8'hac))) >> reg19)});
        end
      reg21 <= wire11[(2'h3):(2'h2)];
      reg22 <= $signed(wire9[(4'h8):(3'h7)]);
    end
  always
    @(posedge clk) begin
      reg23 <= wire9[(3'h6):(1'h1)];
      if ($unsigned($unsigned(({(reg13 ? wire9 : reg13),
          reg22} * reg18[(4'h8):(4'h8)]))))
        begin
          if (reg22[(3'h5):(2'h2)])
            begin
              reg24 <= $unsigned((+reg18[(2'h2):(1'h0)]));
            end
          else
            begin
              reg24 <= reg15;
            end
          reg25 <= (8'ha5);
          reg26 <= (~^$signed(reg14[(2'h2):(1'h1)]));
          reg27 <= ({$unsigned(((reg24 >> reg13) == (!wire7))), reg19} ?
              wire10 : reg17);
          reg28 <= ((~^{((wire7 ? wire9 : reg27) ? (!reg25) : (~^reg27)),
              reg21[(4'h9):(4'h8)]}) >> {$signed(((reg22 ? reg18 : reg15) ?
                  $unsigned(reg27) : $unsigned(wire11))),
              $unsigned((wire9[(3'h4):(1'h1)] ?
                  $signed(reg25) : $signed(reg12)))});
        end
      else
        begin
          reg24 <= (wire7[(1'h0):(1'h0)] && wire11);
        end
    end
  assign wire29 = $unsigned({(!((^reg28) * reg14[(1'h1):(1'h0)]))});
  assign wire30 = ((($unsigned($unsigned(reg22)) ?
                          reg13[(3'h4):(2'h3)] : (8'ha8)) ?
                      $unsigned(({reg24} ?
                          reg18[(3'h4):(2'h3)] : (~|reg15))) : reg21) < wire11[(3'h4):(1'h0)]);
  assign wire31 = (~^(^~$signed(wire29[(1'h1):(1'h0)])));
  assign wire32 = $unsigned(((~|$unsigned((reg18 || wire31))) != $unsigned({$unsigned(reg28)})));
  assign wire33 = ({(+{$unsigned(reg18), (|reg13)})} ?
                      ({$signed(((8'hb9) == wire32))} ?
                          (wire8 ?
                              (~^(reg17 ^ reg14)) : (!(^reg22))) : ((reg21[(1'h0):(1'h0)] ?
                                  {(8'hbb), wire8} : (&wire7)) ?
                              (~^{reg22, reg13}) : (reg23 ?
                                  (reg28 ?
                                      wire6 : wire6) : reg26))) : (($signed({wire9}) <= (8'ha2)) ?
                          reg19 : $signed($unsigned($unsigned(wire10)))));
  always
    @(posedge clk) begin
      reg34 <= $unsigned($unsigned({reg23[(2'h2):(1'h1)], wire31}));
      if (wire32[(4'ha):(1'h0)])
        begin
          reg35 <= (+$unsigned($unsigned((~|((8'ha2) ? wire11 : reg25)))));
          reg36 <= (&wire29);
          reg37 <= reg17[(3'h5):(2'h3)];
        end
      else
        begin
          reg35 <= (~&$signed(reg24[(3'h7):(2'h3)]));
          reg36 <= (8'ha5);
          reg37 <= {($unsigned({(8'haa)}) >> (reg19[(4'h9):(2'h2)] && ((reg20 != reg36) ?
                  (~^reg28) : (&wire7))))};
        end
      reg38 <= (+$signed(wire9));
      reg39 <= reg25;
    end
  assign wire40 = reg19[(2'h3):(1'h1)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module50
#( parameter param471 = ((|((((8'hb7) ? (8'hb7) : (8'hb4)) | (&(8'h9d))) ? ({(8'haa), (8'hb8)} ? ((8'had) ? (8'hae) : (8'h9f)) : {(8'hbc), (8'hb5)}) : ((~&(8'h9e)) ? (8'h9c) : (&(7'h42))))) ? (((-{(8'hb4)}) <= (((8'ha8) <= (8'haa)) ^~ ((8'hb7) ? (7'h40) : (8'hae)))) ? ({(&(8'hb8))} ~^ ((~(8'hb0)) ^~ (8'ha8))) : (&(8'ha4))) : (({(-(7'h43)), (|(8'ha0))} >>> (((8'hab) != (8'h9e)) ~^ ((8'had) != (8'ha7)))) ? (^(+((8'haa) ~^ (8'ha4)))) : ((((8'ha6) > (8'h9c)) * (^~(8'had))) >= ((8'hb8) + ((8'ha7) - (8'hb9))))))
, parameter param472 = (~((+param471) - param471)) )
(y, clk, wire51, wire52, wire53, wire54, wire55);
  output wire [(32'h165):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire51;
  input wire signed [(5'h15):(1'h0)] wire52;
  input wire signed [(5'h15):(1'h0)] wire53;
  input wire signed [(5'h12):(1'h0)] wire54;
  input wire [(5'h14):(1'h0)] wire55;
  reg [(4'h9):(1'h0)] reg470 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg469 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg468 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg467 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg466 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire465;
  wire signed [(4'hc):(1'h0)] wire464;
  wire [(3'h7):(1'h0)] wire463;
  wire [(4'h8):(1'h0)] wire461;
  wire signed [(5'h10):(1'h0)] wire103;
  wire [(5'h10):(1'h0)] wire102;
  wire signed [(5'h12):(1'h0)] wire101;
  wire signed [(4'h8):(1'h0)] wire100;
  wire [(5'h13):(1'h0)] wire99;
  wire [(4'h9):(1'h0)] wire98;
  wire [(4'hb):(1'h0)] wire97;
  wire [(4'ha):(1'h0)] wire96;
  reg [(2'h3):(1'h0)] reg95 = (1'h0);
  reg [(4'he):(1'h0)] reg94 = (1'h0);
  reg [(2'h3):(1'h0)] reg93 = (1'h0);
  reg signed [(4'he):(1'h0)] reg92 = (1'h0);
  reg [(5'h10):(1'h0)] reg91 = (1'h0);
  reg [(3'h5):(1'h0)] reg90 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire89;
  wire [(5'h12):(1'h0)] wire88;
  wire signed [(3'h5):(1'h0)] wire87;
  wire [(3'h7):(1'h0)] wire86;
  wire [(4'he):(1'h0)] wire56;
  wire [(4'he):(1'h0)] wire57;
  wire [(3'h7):(1'h0)] wire58;
  wire [(5'h10):(1'h0)] wire84;
  assign y = {reg470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 wire465,
                 wire464,
                 wire463,
                 wire461,
                 wire103,
                 wire102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 wire97,
                 wire96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 wire89,
                 wire88,
                 wire87,
                 wire86,
                 wire56,
                 wire57,
                 wire58,
                 wire84,
                 (1'h0)};
  assign wire56 = ($signed((wire51[(3'h5):(1'h1)] >>> (~^wire54[(2'h2):(2'h2)]))) >>> (~(&$unsigned($unsigned(wire55)))));
  assign wire57 = wire54;
  assign wire58 = (-{{wire51,
                          (wire51 ? $signed(wire53) : wire57[(4'he):(2'h2)])}});
  module59 modinst85 (.clk(clk), .y(wire84), .wire61(wire54), .wire60(wire55), .wire63(wire56), .wire64(wire51), .wire62(wire53));
  assign wire86 = (wire58[(3'h6):(3'h4)] && ($unsigned(wire53) ^~ $signed(wire53[(5'h12):(2'h2)])));
  assign wire87 = wire56[(4'h9):(2'h3)];
  assign wire88 = wire87[(1'h1):(1'h1)];
  assign wire89 = wire87[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg90 <= $signed((wire86 ?
          wire58[(1'h1):(1'h0)] : $signed({{wire52, wire88}})));
      reg91 <= wire52;
      reg92 <= ($unsigned($signed($signed({reg90, wire86}))) >= wire88);
      reg93 <= $unsigned($signed((8'ha3)));
      if (({$signed($unsigned(reg93))} ?
          (+reg91) : $signed((wire52[(4'he):(1'h0)] ^~ wire58))))
        begin
          reg94 <= (~wire56[(1'h1):(1'h1)]);
          reg95 <= $signed(((+wire56[(3'h5):(2'h2)]) < $unsigned(($unsigned(wire88) & reg90[(2'h2):(1'h1)]))));
        end
      else
        begin
          reg94 <= wire56;
        end
    end
  assign wire96 = {reg91};
  assign wire97 = $unsigned(((((reg90 <<< wire51) >> $signed(wire53)) >> ($unsigned((8'hab)) ?
                      $unsigned(reg90) : $unsigned(wire84))) != wire58[(3'h7):(2'h3)]));
  assign wire98 = ($signed((((reg91 ? wire97 : wire97) >= $signed(wire54)) ?
                          (reg92[(2'h2):(1'h1)] ^ wire57[(4'hd):(4'hc)]) : {wire53,
                              reg90[(2'h2):(1'h1)]})) ?
                      $signed($signed(wire87[(1'h0):(1'h0)])) : (^~(~|(reg94 ?
                          (wire56 ? wire96 : wire56) : (wire58 ?
                              wire53 : (8'ha3))))));
  assign wire99 = wire53[(4'h9):(3'h5)];
  assign wire100 = ({(((wire55 ? wire53 : reg94) ?
                                   (wire99 ?
                                       reg95 : wire87) : $unsigned(wire87)) ?
                               {(wire99 || wire98)} : $signed((+wire51))),
                           (({wire96} ? (wire52 <= wire53) : $signed(wire96)) ?
                               wire56 : ($signed((8'ha6)) <= $signed(wire54)))} ?
                       wire88[(4'ha):(4'h9)] : $signed((reg95[(2'h2):(2'h2)] ?
                           (~reg93[(1'h1):(1'h1)]) : wire89)));
  assign wire101 = reg93;
  assign wire102 = wire96[(3'h5):(1'h0)];
  assign wire103 = $unsigned(((((8'ha4) ? (!wire99) : reg92[(3'h4):(3'h4)]) ?
                           reg93[(1'h0):(1'h0)] : wire57[(3'h7):(2'h2)]) ?
                       ((reg90 <= $unsigned((8'hb6))) ?
                           wire97[(4'h8):(1'h0)] : wire53[(4'he):(4'hc)]) : (~&wire102[(4'he):(2'h2)])));
  module104 modinst462 (.wire108(wire51), .wire106(wire101), .y(wire461), .wire105(wire99), .clk(clk), .wire107(wire52));
  assign wire463 = wire87;
  assign wire464 = (|wire99[(3'h7):(3'h4)]);
  assign wire465 = ((($signed(wire52[(1'h0):(1'h0)]) | $unsigned((wire58 || wire103))) ?
                       ((!wire100) ?
                           $unsigned(reg91[(4'hf):(4'h8)]) : (8'ha8)) : wire463) * (($signed($unsigned(wire57)) ?
                           (wire84[(2'h2):(1'h1)] ?
                               (wire102 == wire464) : reg90) : $unsigned(((8'ha0) ?
                               (8'h9d) : wire89))) ?
                       (~^((^reg91) ? {wire99, (8'hb1)} : wire56)) : wire84));
  always
    @(posedge clk) begin
      reg466 <= ($signed(wire97[(3'h4):(2'h3)]) ?
          wire97[(2'h2):(1'h0)] : $unsigned($signed(($signed(wire103) ?
              (wire55 ? wire97 : wire461) : $unsigned(wire103)))));
      if ($unsigned($signed($signed(((reg92 ?
          reg95 : reg93) ^~ $signed(wire461))))))
        begin
          if ((wire464 ? (-{$unsigned((&wire86))}) : wire102[(4'hc):(2'h3)]))
            begin
              reg467 <= ($unsigned($unsigned({$signed(reg93), (&wire96)})) ?
                  wire88[(3'h4):(2'h3)] : wire54);
              reg468 <= $signed(($signed({{(8'ha1)}}) >> (|(!((8'h9d) ?
                  reg91 : (8'ha8))))));
              reg469 <= $unsigned((-reg92));
              reg470 <= wire97[(4'h9):(1'h1)];
            end
          else
            begin
              reg467 <= $signed(wire53);
            end
        end
      else
        begin
          reg467 <= $signed(wire53[(1'h0):(1'h0)]);
          reg468 <= $unsigned({$unsigned(reg93)});
          reg469 <= wire53;
          reg470 <= ((wire86 ?
              (((^reg94) >= (wire463 ?
                  wire463 : reg468)) ~^ wire53) : (reg470[(2'h2):(1'h1)] ?
                  (8'hab) : wire57[(3'h7):(3'h6)])) << {$unsigned($signed(wire87[(1'h1):(1'h1)]))});
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module104
#( parameter param460 = ((~^(^(((8'ha8) < (8'hbd)) ? (|(8'ha6)) : ((7'h43) ? (8'h9e) : (7'h40))))) ? (({((8'hb4) ? (7'h43) : (8'hbc))} ? ((!(7'h44)) ? {(8'had)} : (8'ha0)) : ({(7'h44)} >>> ((8'hbe) ? (8'h9f) : (8'ha7)))) ? {(((8'h9d) ? (7'h40) : (8'hba)) ? (7'h44) : (8'h9d))} : (~(8'ha4))) : ((-(^~((8'ha9) ? (8'hbb) : (7'h41)))) ? ((^~{(8'hb2), (8'ha5)}) ? (|((8'hb8) ^~ (8'hb9))) : ({(7'h43)} >>> ((8'hb9) ? (8'hbd) : (8'ha5)))) : ((~(~&(8'hbe))) ? ((8'hba) ? ((8'hbf) ? (8'ha7) : (8'hb2)) : ((8'hbf) != (7'h43))) : (((8'ha6) | (8'hba)) <<< ((8'hbd) * (8'ha9)))))) )
(y, clk, wire105, wire106, wire107, wire108);
  output wire [(32'h434):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire105;
  input wire [(2'h3):(1'h0)] wire106;
  input wire [(5'h13):(1'h0)] wire107;
  input wire signed [(3'h7):(1'h0)] wire108;
  wire signed [(4'hb):(1'h0)] wire458;
  wire [(5'h14):(1'h0)] wire271;
  wire signed [(5'h10):(1'h0)] wire270;
  wire signed [(4'hf):(1'h0)] wire269;
  reg [(5'h14):(1'h0)] reg109 = (1'h0);
  reg [(3'h5):(1'h0)] reg110 = (1'h0);
  reg [(3'h4):(1'h0)] reg111 = (1'h0);
  reg [(4'hf):(1'h0)] reg112 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg113 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg114 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg115 = (1'h0);
  reg [(4'h8):(1'h0)] reg116 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg117 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg118 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg119 = (1'h0);
  reg [(2'h2):(1'h0)] reg120 = (1'h0);
  reg [(4'hf):(1'h0)] reg121 = (1'h0);
  reg [(4'h8):(1'h0)] reg122 = (1'h0);
  reg [(5'h11):(1'h0)] reg123 = (1'h0);
  reg [(4'hb):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg125 = (1'h0);
  reg [(3'h7):(1'h0)] reg126 = (1'h0);
  reg [(5'h13):(1'h0)] reg127 = (1'h0);
  wire [(5'h10):(1'h0)] wire128;
  wire signed [(4'ha):(1'h0)] wire129;
  reg [(4'hb):(1'h0)] reg130 = (1'h0);
  reg [(5'h12):(1'h0)] reg131 = (1'h0);
  reg [(4'hc):(1'h0)] reg132 = (1'h0);
  reg [(2'h2):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg135 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg136 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg137 = (1'h0);
  reg [(4'h8):(1'h0)] reg138 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg139 = (1'h0);
  reg signed [(4'he):(1'h0)] reg140 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg142 = (1'h0);
  wire [(4'he):(1'h0)] wire143;
  reg [(4'hb):(1'h0)] reg144 = (1'h0);
  reg [(5'h10):(1'h0)] reg145 = (1'h0);
  reg [(3'h4):(1'h0)] reg146 = (1'h0);
  reg [(5'h14):(1'h0)] reg147 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg148 = (1'h0);
  reg [(4'he):(1'h0)] reg149 = (1'h0);
  reg [(5'h14):(1'h0)] reg150 = (1'h0);
  reg [(4'hf):(1'h0)] reg151 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg152 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg154 = (1'h0);
  reg [(5'h10):(1'h0)] reg155 = (1'h0);
  reg [(4'he):(1'h0)] reg156 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire157;
  reg signed [(2'h3):(1'h0)] reg158 = (1'h0);
  reg [(5'h15):(1'h0)] reg159 = (1'h0);
  reg [(5'h15):(1'h0)] reg160 = (1'h0);
  reg [(5'h13):(1'h0)] reg161 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg162 = (1'h0);
  reg [(4'he):(1'h0)] reg163 = (1'h0);
  reg [(5'h13):(1'h0)] reg164 = (1'h0);
  reg [(5'h13):(1'h0)] reg165 = (1'h0);
  reg [(4'h9):(1'h0)] reg166 = (1'h0);
  reg [(4'he):(1'h0)] reg167 = (1'h0);
  reg [(3'h7):(1'h0)] reg168 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg169 = (1'h0);
  reg [(5'h13):(1'h0)] reg170 = (1'h0);
  reg [(5'h11):(1'h0)] reg171 = (1'h0);
  wire [(2'h2):(1'h0)] wire172;
  wire [(4'he):(1'h0)] wire173;
  wire signed [(4'ha):(1'h0)] wire174;
  wire [(5'h12):(1'h0)] wire175;
  wire [(4'ha):(1'h0)] wire176;
  reg [(4'h8):(1'h0)] reg177 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg178 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg179 = (1'h0);
  reg [(5'h13):(1'h0)] reg180 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg182 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg183 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg184 = (1'h0);
  reg [(5'h15):(1'h0)] reg185 = (1'h0);
  reg [(3'h4):(1'h0)] reg186 = (1'h0);
  reg [(2'h2):(1'h0)] reg187 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg188 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire267;
  assign y = {wire458,
                 wire271,
                 wire270,
                 wire269,
                 reg109,
                 reg110,
                 reg111,
                 reg112,
                 reg113,
                 reg114,
                 reg115,
                 reg116,
                 reg117,
                 reg118,
                 reg119,
                 reg120,
                 reg121,
                 reg122,
                 reg123,
                 reg124,
                 reg125,
                 reg126,
                 reg127,
                 wire128,
                 wire129,
                 reg130,
                 reg131,
                 reg132,
                 reg133,
                 reg134,
                 reg135,
                 reg136,
                 reg137,
                 reg138,
                 reg139,
                 reg140,
                 reg141,
                 reg142,
                 wire143,
                 reg144,
                 reg145,
                 reg146,
                 reg147,
                 reg148,
                 reg149,
                 reg150,
                 reg151,
                 reg152,
                 reg153,
                 reg154,
                 reg155,
                 reg156,
                 wire157,
                 reg158,
                 reg159,
                 reg160,
                 reg161,
                 reg162,
                 reg163,
                 reg164,
                 reg165,
                 reg166,
                 reg167,
                 reg168,
                 reg169,
                 reg170,
                 reg171,
                 wire172,
                 wire173,
                 wire174,
                 wire175,
                 wire176,
                 reg177,
                 reg178,
                 reg179,
                 reg180,
                 reg181,
                 reg182,
                 reg183,
                 reg184,
                 reg185,
                 reg186,
                 reg187,
                 reg188,
                 wire267,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg109 <= {{$unsigned({wire108[(1'h0):(1'h0)], wire107}),
              wire106[(2'h2):(2'h2)]}};
      if (wire106[(2'h2):(1'h1)])
        begin
          if ($unsigned(wire108[(2'h2):(1'h1)]))
            begin
              reg110 <= wire108[(2'h2):(2'h2)];
              reg111 <= ($signed($unsigned((reg110 + (~^reg110)))) ?
                  {(-{reg110[(2'h3):(2'h2)]})} : $signed((&{{wire105},
                      {wire108, wire105}})));
              reg112 <= ({wire107,
                  $signed($unsigned(((8'hbe) * reg110)))} > $unsigned($unsigned($unsigned(((8'ha6) << reg109)))));
            end
          else
            begin
              reg110 <= $signed({$signed($signed({reg109}))});
            end
          if ($unsigned(reg111))
            begin
              reg113 <= $signed($signed($unsigned(((reg111 ? reg111 : (8'hb9)) ?
                  $signed(reg110) : reg110))));
              reg114 <= $unsigned(((reg110 >>> $unsigned((^wire106))) ^ $unsigned(((wire105 <= reg109) >> wire107))));
            end
          else
            begin
              reg113 <= ($signed({((wire108 ? reg112 : reg111) ^ wire105)}) ?
                  ($unsigned(reg114[(1'h0):(1'h0)]) ?
                      ($unsigned($unsigned(wire106)) ?
                          wire106[(1'h1):(1'h0)] : (-$signed(wire108))) : $signed((8'hbb))) : (^reg112));
              reg114 <= (-(&reg110));
            end
          if (wire105)
            begin
              reg115 <= $unsigned($signed({$unsigned((+reg113)),
                  (wire106[(1'h0):(1'h0)] ?
                      (wire106 ? reg113 : reg112) : (reg111 ?
                          wire106 : reg111))}));
              reg116 <= reg115;
              reg117 <= wire106[(1'h0):(1'h0)];
              reg118 <= ((8'ha2) ?
                  $signed($unsigned({$unsigned(reg113)})) : (wire106 != $unsigned(reg111[(3'h4):(2'h2)])));
              reg119 <= $unsigned(reg115);
            end
          else
            begin
              reg115 <= $signed((8'hb3));
            end
          reg120 <= (reg116[(2'h3):(1'h1)] ?
              $unsigned(reg113) : $unsigned($signed((wire107[(1'h1):(1'h0)] ?
                  $signed(reg111) : (reg119 >>> reg119)))));
          if (wire105)
            begin
              reg121 <= reg111[(3'h4):(1'h0)];
              reg122 <= (&reg115[(1'h1):(1'h1)]);
              reg123 <= ((!$unsigned($unsigned((7'h44)))) ? (8'hab) : reg110);
              reg124 <= (({((^reg117) <= reg111[(2'h2):(1'h0)])} ?
                  (((-reg112) ?
                      {reg110} : (~reg110)) >= $signed((reg116 || (8'hb5)))) : ((^~(reg121 > wire108)) & $unsigned(reg112))) + (8'hbb));
              reg125 <= ($unsigned($signed($unsigned($unsigned((8'hb6))))) + {(reg122[(1'h0):(1'h0)] ?
                      reg112[(4'hc):(3'h4)] : {$unsigned(reg114),
                          reg124[(4'h8):(3'h5)]}),
                  reg112[(4'hf):(4'he)]});
            end
          else
            begin
              reg121 <= reg121;
              reg122 <= (!(reg113[(2'h3):(2'h2)] ?
                  (~((reg125 ? reg109 : wire105) >= (wire107 ?
                      reg125 : reg121))) : reg110[(1'h1):(1'h0)]));
              reg123 <= (reg111 ?
                  (&reg123) : {(-((reg124 << reg115) ?
                          {reg113, (8'hbf)} : {(8'ha3), reg111}))});
              reg124 <= {reg116};
            end
        end
      else
        begin
          if (reg121[(1'h0):(1'h0)])
            begin
              reg110 <= {{$signed(($unsigned((8'ha0)) * $unsigned(reg114)))},
                  reg124[(4'h8):(3'h4)]};
              reg111 <= $signed(wire105[(4'hb):(1'h1)]);
            end
          else
            begin
              reg110 <= $unsigned((8'hac));
              reg111 <= (reg115 ?
                  ((^~((reg125 ? reg123 : (8'h9c)) <<< (8'hb4))) ?
                      (8'hbd) : $signed((8'had))) : ($unsigned(reg121[(1'h0):(1'h0)]) != (8'hb1)));
              reg112 <= $signed(reg110);
              reg113 <= $signed($signed({({reg117} ?
                      reg117[(4'h9):(4'h9)] : reg122)}));
              reg114 <= $signed($unsigned(((~^(wire106 ?
                  reg116 : wire106)) != $unsigned($signed(wire106)))));
            end
        end
      reg126 <= wire107[(1'h0):(1'h0)];
      reg127 <= (&$unsigned($unsigned(((wire105 * reg126) ?
          wire105 : reg123))));
    end
  assign wire128 = (|($signed($signed(reg119[(3'h4):(1'h0)])) & (wire105[(3'h7):(1'h0)] ?
                       $unsigned((reg123 << wire106)) : $signed($signed(reg124)))));
  assign wire129 = (reg113 ?
                       $signed((((!reg114) ^ (|wire107)) != reg120)) : reg125);
  always
    @(posedge clk) begin
      if ({((~|$signed((reg112 | reg114))) ?
              wire106[(1'h0):(1'h0)] : wire105[(3'h5):(1'h0)])})
        begin
          if ((($unsigned(reg110[(1'h0):(1'h0)]) > ((!(^(8'hbd))) ?
                  $signed($unsigned(reg122)) : {reg117, $signed(wire108)})) ?
              {(({wire108} ? (8'ha8) : (~^reg122)) ?
                      ((wire106 ?
                          (8'ha9) : wire128) * ((7'h41) || wire108)) : ((wire128 ?
                          reg110 : reg111) ^ wire108[(1'h0):(1'h0)]))} : $signed(reg111)))
            begin
              reg130 <= {(!$signed({(~^reg117)}))};
              reg131 <= $unsigned(($signed((~&{reg110,
                  wire105})) - {$signed($unsigned(reg130))}));
              reg132 <= (~^(^~reg121));
              reg133 <= {$unsigned(wire128[(4'h9):(2'h2)])};
            end
          else
            begin
              reg130 <= ({$signed($unsigned(reg113[(3'h5):(2'h2)]))} > reg115[(3'h4):(2'h2)]);
            end
          if (($unsigned(($signed({reg120}) ?
                  $signed($signed(reg110)) : wire108[(3'h6):(1'h0)])) ?
              (reg125[(3'h7):(3'h6)] ?
                  reg126 : reg121[(3'h5):(1'h1)]) : ({$unsigned(reg109),
                      $signed(reg130)} ?
                  (^~reg120) : $signed({((8'h9c) ? reg119 : reg119)}))))
            begin
              reg134 <= $signed(reg125[(1'h1):(1'h1)]);
              reg135 <= {(8'ha5),
                  (((reg120 ?
                      reg119 : reg122[(1'h0):(1'h0)]) ^~ reg114) <<< (~^((wire106 <= reg131) ?
                      (reg134 ? reg115 : reg132) : reg109)))};
            end
          else
            begin
              reg134 <= $unsigned($signed(reg121[(4'hb):(3'h5)]));
            end
          reg136 <= reg123[(4'hf):(2'h2)];
        end
      else
        begin
          if (($signed(reg124[(4'ha):(1'h1)]) >> (((reg110[(3'h4):(1'h0)] + $signed(reg112)) ?
              ({reg135} ?
                  (wire128 ?
                      reg126 : reg111) : $unsigned(reg133)) : $unsigned($unsigned(reg132))) << reg113)))
            begin
              reg130 <= (reg117 <= ((reg123 ?
                      $signed((+reg127)) : $unsigned($signed(reg121))) ?
                  ($unsigned($unsigned((8'hb9))) ?
                      ($unsigned(wire128) ?
                          $unsigned(reg112) : $unsigned((8'hb3))) : ($signed((8'ha7)) <= $unsigned(reg112))) : {(~&$unsigned(reg134))}));
              reg131 <= (+({(wire128[(3'h4):(2'h2)] ?
                          ((8'hb1) ? reg109 : reg136) : (8'hb7)),
                      reg119} ?
                  wire107[(2'h3):(2'h2)] : reg127));
            end
          else
            begin
              reg130 <= (((|reg118) ?
                  reg118[(3'h5):(2'h3)] : $unsigned(((!reg136) ?
                      $unsigned((8'hba)) : (&reg123)))) >> $signed({(^~(wire129 && reg134))}));
              reg131 <= (reg112 ~^ (!reg111));
              reg132 <= reg124;
            end
          if ($signed(((({reg132, wire105} ?
                  (+(8'ha7)) : $unsigned(reg123)) >>> reg133[(1'h1):(1'h0)]) ?
              $unsigned($unsigned((reg113 ? reg132 : (8'hba)))) : reg116)))
            begin
              reg133 <= reg118;
            end
          else
            begin
              reg133 <= {$unsigned((8'hbd)), wire128};
              reg134 <= (!$unsigned({reg133[(1'h0):(1'h0)]}));
              reg135 <= ($signed($signed(($unsigned(reg109) <<< reg118[(4'h8):(3'h6)]))) ?
                  $unsigned(((reg135 * wire108[(3'h5):(2'h3)]) >> $signed((8'h9d)))) : (reg135[(3'h6):(2'h3)] == $unsigned($signed(((8'ha5) * (8'hae))))));
              reg136 <= (($unsigned($unsigned($unsigned(reg135))) >>> reg130) + $signed(((-reg122) ?
                  $unsigned(reg119) : wire108[(3'h6):(3'h4)])));
            end
          reg137 <= (reg110[(3'h4):(1'h1)] || $unsigned((((&reg112) <<< {reg114}) == (((7'h44) || reg127) >= (~&reg113)))));
          reg138 <= reg114[(1'h1):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned(((8'hab) ~^ wire108)))
        begin
          reg139 <= reg121[(1'h1):(1'h1)];
          reg140 <= {reg130[(4'ha):(1'h1)]};
          reg141 <= {((wire128[(4'hc):(1'h0)] && (&(&wire128))) ?
                  reg120[(1'h1):(1'h1)] : $signed(({wire106} ~^ reg127)))};
          reg142 <= {$unsigned((((reg138 >>> reg117) + (reg139 <<< (8'ha2))) == $unsigned($signed((8'ha2)))))};
        end
      else
        begin
          reg139 <= ($unsigned(reg123) != $signed($unsigned($signed({reg141}))));
          reg140 <= reg130;
          reg141 <= {wire106, reg134};
        end
    end
  assign wire143 = $unsigned((($unsigned((&reg115)) ?
                       ((reg141 ? wire107 : wire128) ?
                           reg119 : (wire108 ?
                               reg139 : reg136)) : ($unsigned(reg141) & (~&reg109))) && ((((7'h41) ?
                               reg133 : (8'ha1)) ?
                           (~^reg132) : $unsigned(reg118)) ?
                       reg133[(1'h1):(1'h1)] : $signed($unsigned(reg140)))));
  always
    @(posedge clk) begin
      if (reg138[(1'h1):(1'h0)])
        begin
          reg144 <= reg110[(3'h5):(1'h1)];
          reg145 <= reg114;
          reg146 <= $unsigned(((($signed(reg112) ~^ (reg145 ?
              (8'ha2) : reg119)) > $unsigned((-reg111))) < $signed(reg136)));
        end
      else
        begin
          reg144 <= $signed((wire107 ?
              $unsigned((8'hae)) : reg127[(2'h2):(2'h2)]));
          if ($signed($unsigned({(+{(8'h9e)})})))
            begin
              reg145 <= $unsigned($unsigned(((|reg119[(2'h2):(1'h1)]) | ((~reg125) || (7'h40)))));
              reg146 <= (~^($unsigned((~reg124)) || {$unsigned((reg144 <<< reg137))}));
            end
          else
            begin
              reg145 <= (&reg118);
              reg146 <= $signed((reg138 ?
                  ($signed(reg135) ?
                      $unsigned((^reg127)) : reg138[(4'h8):(2'h2)]) : (^reg134)));
              reg147 <= $signed((^~reg138[(2'h3):(2'h2)]));
              reg148 <= ($signed($signed((-reg137))) >>> (~$signed(reg147)));
              reg149 <= (^~$unsigned((reg118 >> $unsigned((reg146 ?
                  reg138 : reg146)))));
            end
          reg150 <= (($signed(({reg147, (8'hb5)} ?
                  (reg144 ? reg149 : reg126) : reg126[(2'h2):(1'h1)])) ?
              {((reg148 - reg146) ?
                      (reg127 ^~ reg146) : (reg112 ?
                          reg149 : reg109))} : $signed($signed((reg121 && reg138)))) >= $unsigned({$signed((~&reg141)),
              $signed((^wire106))}));
        end
      reg151 <= reg130[(4'hb):(3'h6)];
      reg152 <= $signed(($unsigned(reg151) - (wire106[(1'h0):(1'h0)] << ((8'haf) << (~^wire128)))));
      if ((!reg144))
        begin
          reg153 <= $signed(reg127[(3'h7):(1'h0)]);
        end
      else
        begin
          reg153 <= ((wire105 <= $signed(($signed(wire107) ?
                  reg116 : (reg151 ? reg115 : reg118)))) ?
              (reg149[(4'h9):(1'h0)] ?
                  reg125[(4'ha):(2'h2)] : (8'ha8)) : ((((reg118 ~^ reg121) ?
                      (reg115 ? reg109 : reg142) : (reg118 && reg115)) ?
                  {$signed(wire105),
                      (reg123 && wire107)} : ((^reg115) & reg122)) | reg149[(3'h7):(2'h2)]));
          reg154 <= ((~$unsigned($unsigned(reg139[(1'h0):(1'h0)]))) ?
              reg140 : (wire143[(4'hb):(4'h9)] ?
                  reg151 : ($unsigned(wire105) ?
                      $signed((wire128 <= reg146)) : {((8'h9c) ?
                              wire143 : reg150)})));
          reg155 <= ($unsigned((&(reg154 ?
              $unsigned(reg114) : reg126))) * ($signed($unsigned($unsigned((8'hb1)))) ?
              ((&reg115[(2'h2):(1'h0)]) ?
                  {(reg135 ? reg144 : reg125)} : {(wire143 ? (8'h9f) : (7'h43)),
                      $unsigned(reg146)}) : {($signed(reg141) ^ (wire108 ?
                      reg133 : (8'hb7))),
                  ($unsigned(reg135) ? reg112 : wire106[(1'h1):(1'h1)])}));
        end
      reg156 <= ((-(8'ha7)) + $unsigned((reg114 ?
          ($signed(wire106) < (wire107 ~^ reg110)) : $unsigned($unsigned(reg135)))));
    end
  assign wire157 = reg142;
  always
    @(posedge clk) begin
      if ({((~^((|(8'hbc)) ? (~^reg141) : $unsigned(reg144))) >= ((!{reg127}) ?
              reg146[(2'h2):(1'h1)] : reg115))})
        begin
          reg158 <= reg121;
          reg159 <= $unsigned((reg111 ?
              ({((7'h41) << (7'h44)), (~wire157)} ?
                  $signed(reg135) : reg152[(2'h2):(1'h0)]) : reg155));
          reg160 <= (($unsigned((!(7'h42))) >>> ((~|$unsigned(reg116)) ?
              reg130 : (8'hb4))) >= $unsigned(reg133));
          reg161 <= wire107;
        end
      else
        begin
          reg158 <= reg113;
          if ((~&{wire143, (8'hba)}))
            begin
              reg159 <= reg159[(5'h14):(1'h1)];
              reg160 <= $unsigned((8'ha7));
              reg161 <= (reg134[(1'h1):(1'h1)] ?
                  ((|wire107) <= ((reg152 > (wire128 ? reg154 : reg123)) ?
                      $signed((wire129 ? reg116 : reg121)) : (^~(reg131 ?
                          reg130 : (8'ha8))))) : reg156);
              reg162 <= $signed($signed(reg160[(2'h3):(2'h2)]));
            end
          else
            begin
              reg159 <= reg139;
              reg160 <= (+reg125[(1'h0):(1'h0)]);
              reg161 <= reg153[(1'h1):(1'h1)];
            end
          if (wire157[(1'h0):(1'h0)])
            begin
              reg163 <= reg122[(1'h0):(1'h0)];
              reg164 <= $unsigned({{(~(reg161 >> reg112))}});
            end
          else
            begin
              reg163 <= $unsigned($unsigned((((reg146 == reg149) == reg145) < ((reg137 && reg152) >> reg156))));
              reg164 <= (((((wire129 && reg159) ? reg149 : wire107) ?
                      ((+wire129) <<< {reg158}) : reg116[(2'h2):(2'h2)]) ?
                  reg109 : (((reg124 ~^ reg119) | $signed(reg142)) ?
                      $unsigned(((8'ha0) ?
                          (8'hba) : (8'h9d))) : (~reg124))) >> (!(($unsigned(reg114) - (~|(7'h40))) >> {$unsigned(wire157)})));
              reg165 <= $signed($signed($unsigned((~|(8'hb0)))));
              reg166 <= (!reg118);
            end
          reg167 <= {(8'ha9),
              (({(&reg113)} ?
                      (wire129 ?
                          $signed(reg159) : {reg115, wire128}) : ((7'h40) ?
                          (|reg150) : $unsigned(wire157))) ?
                  {((+reg137) ?
                          reg130 : reg122[(3'h5):(2'h2)])} : (((&reg123) == {(8'ha6)}) > reg111))};
          if (reg159)
            begin
              reg168 <= reg150[(5'h12):(4'ha)];
              reg169 <= reg119;
              reg170 <= ((8'haf) ?
                  {{$signed($signed(reg146)),
                          ($signed((8'ha9)) ?
                              ((8'hbf) ? wire128 : reg167) : (wire143 ?
                                  reg167 : reg123))}} : {(($unsigned(reg130) >= (-reg132)) == $unsigned($signed(reg148))),
                      $signed((reg113 ?
                          (reg119 ? (8'hbc) : (8'hb0)) : $unsigned((8'h9d))))});
              reg171 <= ($signed($signed(((~reg152) ?
                  ((8'hac) ?
                      reg132 : (8'hab)) : $unsigned((8'ha9))))) >>> (+reg119));
            end
          else
            begin
              reg168 <= (wire129[(3'h4):(2'h2)] ?
                  (-$unsigned($signed($unsigned(reg126)))) : (($signed($signed(reg123)) ~^ (^~(8'h9f))) > $signed(($unsigned(reg171) && wire129))));
              reg169 <= reg155;
              reg170 <= ((~&(8'ha4)) ?
                  $unsigned($signed(reg122)) : {(+(8'hb8))});
              reg171 <= wire157;
            end
        end
    end
  assign wire172 = (~&reg150);
  assign wire173 = ((+reg154) ?
                       {({$signed(reg167)} ?
                               $unsigned((reg111 * (8'had))) : $signed(reg171[(1'h0):(1'h0)]))} : $signed(reg170));
  assign wire174 = reg155[(4'hf):(4'hd)];
  assign wire175 = $unsigned(reg118[(5'h14):(3'h5)]);
  assign wire176 = ((8'hbc) ~^ {{reg152[(2'h2):(2'h2)]},
                       reg142[(5'h14):(4'h9)]});
  always
    @(posedge clk) begin
      reg177 <= (~^$unsigned((8'hb6)));
      if (($signed((~|{wire106[(2'h3):(2'h2)],
          $signed((8'hab))})) <= (&reg141)))
        begin
          reg178 <= (($signed(((7'h42) ? reg136 : (8'hb1))) ?
              ($unsigned($unsigned(reg150)) + reg164) : {$unsigned(reg155),
                  ($signed(wire176) ?
                      reg149[(3'h4):(3'h4)] : $unsigned(reg120))}) != (+$unsigned({$signed((8'hb3))})));
          reg179 <= $signed(($signed($unsigned((reg177 < (8'hbb)))) ?
              reg131 : (wire105[(4'he):(4'he)] & $signed((!reg137)))));
          reg180 <= $unsigned($signed(($unsigned((reg123 <<< wire105)) >> $signed(reg170[(5'h11):(4'h9)]))));
          if ($signed($unsigned((~|((reg145 <<< reg153) != (reg120 ?
              reg116 : reg126))))))
            begin
              reg181 <= (&(!($signed(reg149[(3'h6):(2'h2)]) ?
                  (!(~reg180)) : reg132)));
              reg182 <= ($unsigned({$unsigned((~^(8'hb3)))}) ?
                  $unsigned(reg179) : $signed(((reg136 >= $signed(reg134)) ?
                      $signed((+reg135)) : ((reg155 ? reg151 : reg162) ?
                          (reg159 & (8'hb2)) : (reg120 ? reg131 : (8'h9e))))));
              reg183 <= $signed((&(reg142 ?
                  reg121[(3'h7):(3'h6)] : $unsigned($unsigned(wire176)))));
            end
          else
            begin
              reg181 <= ($unsigned({reg179, (8'hb6)}) ?
                  $signed(reg126[(3'h7):(3'h7)]) : $signed((7'h44)));
              reg182 <= $signed(($unsigned((~&(wire108 ? wire172 : reg132))) ?
                  (^~(~|reg153[(1'h1):(1'h1)])) : reg124));
            end
          if ($signed((8'had)))
            begin
              reg184 <= $unsigned($signed(reg150));
              reg185 <= reg130;
              reg186 <= ((($unsigned(((7'h42) ?
                          reg122 : reg182)) >= $unsigned(wire173)) ?
                      (reg159[(5'h14):(3'h7)] & (reg140[(4'h9):(4'h8)] ?
                          wire175 : reg117)) : $unsigned(reg158[(2'h3):(2'h2)])) ?
                  $unsigned($unsigned(($signed(reg109) != (reg146 ^ reg127)))) : ($signed(reg170) < $signed(reg130)));
              reg187 <= $unsigned(reg161[(4'he):(1'h1)]);
            end
          else
            begin
              reg184 <= ($unsigned($unsigned((8'hbc))) >>> (-(reg166[(2'h3):(2'h3)] != ((wire157 + wire105) <= (~(7'h44))))));
            end
        end
      else
        begin
          if (reg138[(4'h8):(3'h5)])
            begin
              reg178 <= (reg168[(3'h7):(3'h5)] >>> {$signed(((reg169 <= reg155) ?
                      (reg155 >> reg169) : (reg151 * reg110))),
                  $unsigned($signed((|reg156)))});
              reg179 <= ((~|$unsigned($signed((~|reg124)))) ?
                  (($signed((7'h41)) ?
                      (reg168 ~^ (|reg133)) : (reg147 ?
                          {reg141,
                              reg178} : $unsigned(reg135))) == (|reg181[(2'h3):(2'h2)])) : (reg116 <= wire143[(4'ha):(3'h4)]));
              reg180 <= $unsigned(($signed(reg145[(3'h6):(2'h2)]) ?
                  ($signed((~&reg122)) << (+(reg169 >> reg166))) : (-(~^(!wire106)))));
              reg181 <= (^({(reg130 <<< reg115),
                  ((-reg154) << reg110)} | $signed($unsigned(wire105[(5'h12):(3'h4)]))));
            end
          else
            begin
              reg178 <= ({($signed(((7'h44) >= (8'ha0))) > $signed(reg153[(2'h2):(1'h0)]))} >> {$unsigned((reg113 + (reg121 ?
                      reg138 : reg183)))});
              reg179 <= reg171[(4'hb):(2'h3)];
            end
          if (((~reg154[(2'h3):(1'h1)]) ? $unsigned(reg122) : {reg109}))
            begin
              reg182 <= reg155[(3'h5):(3'h5)];
              reg183 <= wire175;
              reg184 <= reg144[(2'h3):(1'h1)];
            end
          else
            begin
              reg182 <= $unsigned(((+(reg151 ?
                  $signed(reg127) : $signed(reg132))) - ($unsigned($unsigned(reg142)) && reg187)));
              reg183 <= $signed(wire106[(1'h0):(1'h0)]);
            end
          reg185 <= ($unsigned($unsigned((((8'ha5) ?
                  (8'had) : reg121) >> (wire143 ? reg132 : reg163)))) ?
              reg136 : $unsigned(reg118[(5'h13):(2'h2)]));
          if ((((+($signed(wire107) > reg147[(3'h5):(3'h5)])) ?
                  (reg137 ^ ($signed(wire128) < (reg177 >>> reg166))) : $signed($signed((reg109 <= reg124)))) ?
              (^$unsigned($unsigned(reg142[(4'hd):(1'h1)]))) : reg183[(3'h4):(3'h4)]))
            begin
              reg186 <= ((~(reg153[(5'h11):(1'h1)] ? reg167 : wire108)) ?
                  ($unsigned($unsigned($unsigned(reg162))) != $unsigned($signed($unsigned(reg170)))) : reg184[(3'h6):(2'h3)]);
            end
          else
            begin
              reg186 <= $signed(reg149);
            end
          reg187 <= $signed(reg162);
        end
      reg188 <= ({reg137[(2'h3):(2'h3)],
              $signed(({reg118} ? reg135[(4'h8):(1'h1)] : reg118))} ?
          $signed($signed(reg112)) : (wire173[(2'h3):(1'h1)] << $unsigned(reg130[(4'h9):(4'h9)])));
    end
  module189 modinst268 (wire267, clk, wire107, reg182, reg165, reg162, reg181);
  assign wire269 = ({$signed(((reg159 - wire174) ?
                               reg177[(3'h4):(3'h4)] : reg154))} ?
                       reg166 : (|({reg121[(1'h0):(1'h0)],
                               (reg137 ? wire143 : (8'hbe))} ?
                           reg119[(4'h9):(3'h6)] : (&$signed(reg184)))));
  assign wire270 = reg186;
  assign wire271 = $signed(($unsigned(((-(8'ha6)) <= (~wire143))) ?
                       (|reg166[(2'h2):(2'h2)]) : reg117));
  module272 modinst459 (wire458, clk, reg167, wire157, wire107, reg166);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module59
#(parameter param82 = (^~(8'ha4)), parameter param83 = param82)
(y, clk, wire64, wire63, wire62, wire61, wire60);
  output wire [(32'hb1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire64;
  input wire signed [(4'he):(1'h0)] wire63;
  input wire signed [(5'h15):(1'h0)] wire62;
  input wire signed [(5'h12):(1'h0)] wire61;
  input wire signed [(5'h14):(1'h0)] wire60;
  wire [(5'h12):(1'h0)] wire81;
  wire signed [(3'h5):(1'h0)] wire80;
  reg [(5'h12):(1'h0)] reg79 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg78 = (1'h0);
  reg [(2'h3):(1'h0)] reg77 = (1'h0);
  reg [(4'hc):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg75 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg72 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg70 = (1'h0);
  reg [(3'h6):(1'h0)] reg69 = (1'h0);
  reg [(2'h2):(1'h0)] reg68 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg67 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire66;
  wire signed [(2'h3):(1'h0)] wire65;
  assign y = {wire81,
                 wire80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 wire66,
                 wire65,
                 (1'h0)};
  assign wire65 = wire64;
  assign wire66 = ($signed((8'hbe)) ?
                      {(wire61[(4'h8):(2'h2)] ?
                              wire61 : (^~$unsigned((8'ha0)))),
                          $signed(wire63[(4'he):(4'hc)])} : ((wire61 >> (!(~&(8'hb1)))) ?
                          $unsigned((wire65[(1'h1):(1'h0)] ?
                              $signed(wire64) : wire61[(3'h6):(3'h5)])) : (({wire63,
                                  wire64} ?
                              wire63 : wire62[(4'hf):(1'h1)]) >= $unsigned((+wire65)))));
  always
    @(posedge clk) begin
      if ((((^~($signed(wire65) <= $signed(wire60))) != $unsigned($unsigned(wire61))) ?
          wire64[(2'h3):(2'h3)] : $unsigned(wire61)))
        begin
          if (($signed(wire65) ?
              $unsigned(wire62) : (~|(($unsigned((8'hbd)) + wire64) ?
                  {(~^wire65), $unsigned(wire62)} : (&(wire64 >= (8'ha9)))))))
            begin
              reg67 <= wire65[(2'h3):(2'h3)];
            end
          else
            begin
              reg67 <= (-$unsigned($signed(((wire63 <= wire61) ?
                  {wire62, (8'hb5)} : (+wire64)))));
              reg68 <= (((~|$unsigned((^wire60))) ?
                  ($signed(wire66) != $unsigned($signed(wire60))) : (^$signed(wire66))) < (~&$signed(wire64)));
              reg69 <= $unsigned((|$unsigned($unsigned((~&(8'hb2))))));
              reg70 <= (wire62 ?
                  wire64[(3'h4):(2'h2)] : ($signed($unsigned(wire64[(3'h7):(3'h4)])) == $unsigned($signed($unsigned((8'ha5))))));
              reg71 <= $unsigned({(~$unsigned(((8'hb7) ? wire63 : wire62))),
                  ({((8'haf) >>> wire64)} ?
                      (+(reg68 ? wire61 : reg69)) : ((^~reg69) ?
                          (8'hae) : wire65))});
            end
          reg72 <= {reg69[(3'h4):(1'h0)],
              (({$unsigned(reg68)} <= ($unsigned(wire66) ?
                      (reg70 & (8'hb5)) : $signed(reg67))) ?
                  $unsigned(((reg69 ? reg69 : reg71) ?
                      {wire60} : $unsigned(reg69))) : (($unsigned((8'hba)) ?
                          (^wire61) : wire61) ?
                      $unsigned($unsigned((8'hba))) : ($unsigned(wire62) ?
                          (~&(7'h41)) : wire61)))};
          reg73 <= (wire63[(1'h0):(1'h0)] ?
              $signed(wire62) : (wire60[(5'h14):(2'h2)] >= $signed(reg68)));
          if (wire66[(2'h2):(1'h1)])
            begin
              reg74 <= wire62[(5'h13):(4'hf)];
            end
          else
            begin
              reg74 <= reg68[(1'h1):(1'h0)];
              reg75 <= reg69;
              reg76 <= $signed((reg69[(3'h4):(3'h4)] > ($unsigned(wire60[(4'h9):(3'h6)]) ?
                  $signed(wire63) : (~|wire63))));
              reg77 <= $signed(reg75);
            end
          reg78 <= $unsigned($signed(wire65[(2'h3):(1'h1)]));
        end
      else
        begin
          if (reg67[(3'h4):(2'h3)])
            begin
              reg67 <= (^~(($unsigned($signed(reg75)) ?
                  ({(8'ha0)} + (reg77 < wire61)) : (reg72[(3'h4):(2'h2)] ^ ((8'hb3) >= reg78))) <= reg68));
              reg68 <= reg76[(1'h1):(1'h0)];
              reg69 <= $unsigned((|(!$unsigned((reg68 ? reg71 : reg78)))));
              reg70 <= $signed($signed((((reg70 ?
                      wire63 : reg73) | (reg73 > (8'hb9))) ?
                  ($unsigned(wire60) && (reg73 <<< reg68)) : (|reg68[(1'h1):(1'h1)]))));
              reg71 <= wire65[(2'h3):(1'h1)];
            end
          else
            begin
              reg67 <= (reg75 == wire66);
            end
        end
      reg79 <= (wire61 ?
          (-((((8'h9c) < reg67) && (~&reg73)) ?
              (~&reg75[(3'h4):(2'h2)]) : ($signed(reg76) ?
                  wire63[(3'h6):(1'h0)] : wire60[(2'h3):(1'h0)]))) : reg69);
    end
  assign wire80 = (~&(~^((!$unsigned(reg74)) || (^$signed(reg74)))));
  assign wire81 = $unsigned((wire80 ?
                      (reg77 - wire64[(2'h3):(1'h1)]) : {$unsigned(reg72),
                          (reg79[(1'h1):(1'h0)] * wire65[(2'h2):(1'h0)])}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module272  (y, clk, wire276, wire275, wire274, wire273);
  output wire [(32'h27c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire276;
  input wire signed [(5'h11):(1'h0)] wire275;
  input wire signed [(5'h13):(1'h0)] wire274;
  input wire [(4'h9):(1'h0)] wire273;
  wire signed [(5'h14):(1'h0)] wire397;
  wire signed [(4'ha):(1'h0)] wire328;
  wire signed [(3'h6):(1'h0)] wire303;
  wire signed [(2'h2):(1'h0)] wire302;
  wire [(5'h11):(1'h0)] wire301;
  wire signed [(4'he):(1'h0)] wire300;
  wire signed [(4'he):(1'h0)] wire299;
  wire signed [(3'h5):(1'h0)] wire298;
  wire signed [(4'ha):(1'h0)] wire297;
  wire signed [(2'h2):(1'h0)] wire296;
  reg signed [(3'h4):(1'h0)] reg295 = (1'h0);
  reg [(3'h6):(1'h0)] reg294 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg293 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg292 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg291 = (1'h0);
  reg [(5'h12):(1'h0)] reg290 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg289 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg288 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg286 = (1'h0);
  reg [(5'h12):(1'h0)] reg285 = (1'h0);
  reg [(5'h14):(1'h0)] reg284 = (1'h0);
  reg [(5'h15):(1'h0)] reg283 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg282 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg281 = (1'h0);
  reg [(5'h11):(1'h0)] reg280 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg279 = (1'h0);
  reg [(5'h11):(1'h0)] reg278 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire277;
  wire signed [(5'h15):(1'h0)] wire399;
  wire signed [(3'h7):(1'h0)] wire400;
  reg [(4'hf):(1'h0)] reg401 = (1'h0);
  wire [(5'h14):(1'h0)] wire402;
  reg [(4'he):(1'h0)] reg403 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire404;
  reg signed [(4'he):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg406 = (1'h0);
  reg [(3'h6):(1'h0)] reg407 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg408 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg409 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg410 = (1'h0);
  reg [(3'h7):(1'h0)] reg411 = (1'h0);
  reg [(5'h11):(1'h0)] reg412 = (1'h0);
  reg [(4'h8):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg414 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg415 = (1'h0);
  reg [(4'hc):(1'h0)] reg416 = (1'h0);
  reg [(5'h14):(1'h0)] reg417 = (1'h0);
  wire [(5'h13):(1'h0)] wire456;
  assign y = {wire397,
                 wire328,
                 wire303,
                 wire302,
                 wire301,
                 wire300,
                 wire299,
                 wire298,
                 wire297,
                 wire296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 wire277,
                 wire399,
                 wire400,
                 reg401,
                 wire402,
                 reg403,
                 wire404,
                 reg405,
                 reg406,
                 reg407,
                 reg408,
                 reg409,
                 reg410,
                 reg411,
                 reg412,
                 reg413,
                 reg414,
                 reg415,
                 reg416,
                 reg417,
                 wire456,
                 (1'h0)};
  assign wire277 = wire273;
  always
    @(posedge clk) begin
      reg278 <= ($signed(wire274) ?
          $unsigned(wire276[(3'h5):(2'h2)]) : $signed(wire275));
      if ((((|(-$unsigned(wire276))) ?
          wire276 : $unsigned(wire274[(3'h5):(3'h4)])) & $unsigned((((~&reg278) ~^ (wire275 ?
              wire275 : reg278)) ?
          (+reg278[(4'hf):(3'h6)]) : wire276[(1'h0):(1'h0)]))))
        begin
          reg279 <= wire274[(4'hf):(3'h6)];
          reg280 <= reg279;
        end
      else
        begin
          reg279 <= {wire276[(1'h0):(1'h0)]};
        end
      reg281 <= {(!wire276)};
      reg282 <= $signed(reg280[(4'he):(4'hb)]);
      if ($unsigned(reg279))
        begin
          reg283 <= wire273;
          reg284 <= (8'h9e);
          reg285 <= (8'hb8);
          if (wire277[(5'h15):(4'he)])
            begin
              reg286 <= {(8'hb3), {$unsigned(($signed(reg283) ~^ (+wire273)))}};
              reg287 <= $signed(wire275);
              reg288 <= (reg282 & $unsigned(($unsigned(reg284[(4'h8):(3'h5)]) & reg279)));
              reg289 <= $signed(((((reg285 ^~ reg281) <<< $signed(wire276)) && (|reg287[(1'h0):(1'h0)])) ?
                  $unsigned((|$unsigned(wire274))) : reg280[(1'h0):(1'h0)]));
            end
          else
            begin
              reg286 <= reg285[(2'h3):(2'h3)];
            end
          reg290 <= ((~|(8'had)) ?
              reg279[(3'h4):(1'h0)] : wire277[(5'h11):(4'hf)]);
        end
      else
        begin
          if (reg286)
            begin
              reg283 <= reg283;
            end
          else
            begin
              reg283 <= $unsigned({$unsigned($unsigned(reg282))});
            end
          if ((~&wire273[(2'h2):(1'h0)]))
            begin
              reg284 <= $signed($unsigned(wire276));
              reg285 <= reg282[(4'h9):(1'h0)];
              reg286 <= ((8'ha3) ? reg279[(1'h1):(1'h1)] : reg279);
              reg287 <= {(7'h41),
                  ($unsigned(($unsigned(reg278) ?
                      $signed(wire274) : (reg290 ?
                          reg280 : reg282))) * reg286[(4'ha):(2'h3)])};
            end
          else
            begin
              reg284 <= $signed((^$signed((-((8'hbd) <<< (8'h9f))))));
              reg285 <= $signed(((((~(8'hba)) ?
                      (reg283 > reg290) : (reg288 ^~ reg279)) ?
                  $unsigned((reg282 * reg280)) : ($signed(reg287) == ((7'h44) < (7'h41)))) < (~^{(^~reg280),
                  $unsigned(reg279)})));
              reg286 <= (((reg286[(4'h8):(1'h1)] ?
                          $signed((~reg285)) : $signed((wire274 * wire277))) ?
                      $signed((reg283[(4'hb):(3'h6)] ?
                          reg286[(1'h1):(1'h0)] : reg283)) : ($signed({reg278}) < reg278[(1'h1):(1'h1)])) ?
                  (&$unsigned($signed((~reg288)))) : $unsigned(((-reg287) ?
                      $signed($unsigned(reg280)) : $signed((~|wire273)))));
              reg287 <= (((reg284 ? ((reg280 < reg288) >>> reg280) : reg279) ?
                  $signed(((wire277 ? reg281 : reg287) ?
                      $signed(reg287) : reg286)) : (+$unsigned((reg285 ?
                      reg285 : wire276)))) > (-(7'h40)));
              reg288 <= (^$unsigned((((reg285 ? (8'hbd) : wire275) == ((8'hae) ?
                      wire276 : wire277)) ?
                  (^$unsigned(reg285)) : ($signed((8'haf)) ?
                      reg286[(5'h12):(2'h2)] : $signed(reg279)))));
            end
          reg289 <= ((+$signed(((wire273 ? reg286 : reg283) ?
              wire275[(3'h7):(2'h3)] : {reg290}))) >= reg286[(1'h1):(1'h1)]);
          if ($signed(reg279[(2'h2):(1'h0)]))
            begin
              reg290 <= (((~^wire276) != {((reg282 ?
                          reg279 : (7'h42)) * (reg290 == (8'ha5))),
                      $signed(((8'haf) >>> wire275))}) ?
                  $signed({($unsigned((8'ha8)) ?
                          (reg286 <= reg282) : (reg285 == reg284)),
                      $signed((wire277 >= reg282))}) : (8'hb7));
              reg291 <= $unsigned($unsigned(wire277));
              reg292 <= (!((8'haa) ?
                  (reg282 ?
                      ((-reg285) ?
                          {(8'hbb),
                              (8'hae)} : $unsigned(wire277)) : {$unsigned(wire275)}) : (~&$signed({reg291}))));
              reg293 <= (reg288[(3'h4):(1'h0)] != ({$unsigned(reg284)} << $unsigned($signed($unsigned(reg285)))));
              reg294 <= (($signed((~&$signed(reg282))) ?
                      {{{reg288}}} : (~reg279[(5'h11):(4'hf)])) ?
                  reg288[(1'h0):(1'h0)] : wire273);
            end
          else
            begin
              reg290 <= (8'hb6);
            end
          reg295 <= ((^(reg289 ?
                  ((reg283 << reg286) ? (~&(8'ha6)) : (~|reg294)) : reg278)) ?
              $unsigned(((reg280[(4'h8):(3'h7)] >= (reg280 ?
                  wire277 : wire275)) | $signed($unsigned(reg287)))) : (($unsigned(((8'hbc) || reg283)) << reg288[(3'h5):(1'h0)]) ?
                  $signed($signed((~&reg293))) : $signed({$unsigned(reg280),
                      (^(7'h41))})));
        end
    end
  assign wire296 = (wire273 ? wire276 : $unsigned(wire274));
  assign wire297 = ($unsigned((&$unsigned((reg284 - wire273)))) ?
                       (-(((reg280 ^~ reg282) ?
                           ((8'had) ?
                               (8'hb1) : reg285) : $signed((8'ha3))) << (wire276 ?
                           (wire276 ?
                               (8'haa) : wire273) : (^~reg294)))) : $unsigned((8'h9e)));
  assign wire298 = (($signed(((|reg292) ?
                       (wire274 ?
                           reg290 : reg286) : (reg289 - reg284))) || ($unsigned(wire277) ?
                       (~^(reg283 << (8'ha9))) : reg281)) >>> reg283);
  assign wire299 = {reg289[(3'h5):(2'h2)],
                       (reg289[(3'h7):(1'h1)] | $unsigned(({reg283, wire296} ?
                           reg286[(1'h1):(1'h1)] : $signed(wire298))))};
  assign wire300 = reg289[(3'h7):(2'h3)];
  assign wire301 = reg284;
  assign wire302 = reg290[(3'h5):(1'h1)];
  assign wire303 = reg281;
  module304 modinst329 (.wire307(wire274), .y(wire328), .wire306(reg283), .wire305(reg279), .wire308(reg288), .clk(clk));
  module330 modinst398 (.clk(clk), .wire332(reg288), .wire331(wire276), .wire335(reg281), .y(wire397), .wire334(reg280), .wire333(reg287));
  assign wire399 = (8'hba);
  assign wire400 = reg293[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg401 <= $unsigned($unsigned((8'ha0)));
    end
  assign wire402 = {(+{(((8'haa) ? reg278 : (8'h9f)) * $signed((8'hb7)))}),
                       reg293[(2'h3):(1'h1)]};
  always
    @(posedge clk) begin
      reg403 <= (8'hb6);
    end
  assign wire404 = wire303[(2'h3):(2'h3)];
  always
    @(posedge clk) begin
      if ($unsigned((({(reg281 ? reg286 : wire276)} == (8'hbe)) ?
          $unsigned(reg283) : $unsigned(({wire397,
              (7'h40)} << $unsigned(reg287))))))
        begin
          if ($signed(reg286[(4'hb):(2'h3)]))
            begin
              reg405 <= $signed((!(($signed(reg286) ?
                  reg280 : wire274[(3'h7):(3'h5)]) >= ({reg289} ?
                  reg283[(4'hd):(4'hd)] : $signed((8'h9f))))));
              reg406 <= {reg294};
              reg407 <= {(~&$unsigned(reg289)), (&reg280)};
              reg408 <= $unsigned($unsigned($unsigned((&reg293))));
              reg409 <= $signed((~^reg288));
            end
          else
            begin
              reg405 <= (wire299 ^~ $unsigned((8'ha7)));
              reg406 <= (+reg401[(2'h3):(2'h2)]);
            end
          if (($unsigned($signed($unsigned($unsigned((8'ha5))))) < {(^$unsigned(reg279)),
              $signed((!wire399))}))
            begin
              reg410 <= $signed(reg285);
              reg411 <= $unsigned($unsigned(((~^((8'hb5) > reg291)) != ({reg407,
                      reg290} ?
                  $signed((8'hbd)) : $unsigned(reg291)))));
            end
          else
            begin
              reg410 <= ((~^wire300[(4'h9):(1'h0)]) ? reg407 : wire301);
              reg411 <= $unsigned((&wire273[(3'h5):(1'h1)]));
            end
        end
      else
        begin
          reg405 <= wire397;
          reg406 <= wire296;
          if ($signed((((reg289 >> (8'hb9)) ^ $signed({wire296})) ?
              {(~&wire301)} : reg411[(2'h2):(1'h1)])))
            begin
              reg407 <= {$signed(($signed((+wire298)) ?
                      $signed(reg291) : {{reg409}, (reg410 * reg293)})),
                  (reg403 || reg287)};
              reg408 <= wire300[(1'h0):(1'h0)];
              reg409 <= wire397;
            end
          else
            begin
              reg407 <= wire300[(3'h5):(1'h0)];
              reg408 <= $unsigned(((($unsigned(reg295) << $unsigned(reg284)) ?
                  $signed(wire301) : reg295[(1'h0):(1'h0)]) * ((^(~wire402)) < $unsigned((reg286 ?
                  wire397 : reg278)))));
              reg409 <= $signed(wire296);
            end
        end
      reg412 <= ((reg408 | $signed(reg292[(3'h5):(1'h1)])) != {($unsigned($signed(reg286)) ?
              wire277 : reg411),
          $unsigned((~{wire301, reg291}))});
      if (reg278[(3'h6):(2'h2)])
        begin
          reg413 <= $signed((wire328 ?
              wire328 : (reg412[(4'hd):(3'h5)] ?
                  (reg410[(4'h9):(4'h8)] ?
                      $unsigned(wire276) : (!wire404)) : {reg278,
                      $signed(reg293)})));
          reg414 <= (8'h9f);
          if (((wire276[(3'h5):(3'h5)] != $unsigned(wire300[(3'h7):(3'h6)])) ?
              ((!((reg407 <<< (8'hb2)) < {(8'ha5), reg286})) ?
                  {{(~^reg281), $unsigned(reg407)}} : ($signed((reg281 ?
                          reg295 : reg282)) ?
                      (~&(8'hb7)) : (wire399 | (wire397 ?
                          (8'haf) : reg403)))) : ($signed((+(wire296 ?
                      wire273 : reg414))) ?
                  $unsigned(reg284[(4'hf):(4'hb)]) : ((~|(&wire328)) ?
                      reg283[(3'h4):(3'h4)] : $signed($signed(reg282))))))
            begin
              reg415 <= (|((($signed(wire303) ?
                      (reg283 ?
                          wire299 : reg282) : reg286[(4'hf):(3'h6)]) >> $signed($signed(reg412))) ?
                  {$signed({(8'hb3), reg403}),
                      {(reg406 ? (8'haa) : reg408)}} : (~$signed({wire328}))));
              reg416 <= ($unsigned(({wire328} ?
                      (+reg285) : $unsigned((reg401 ? reg288 : wire399)))) ?
                  ($unsigned($unsigned(reg413)) < (!(~&$unsigned(reg401)))) : $signed(wire296));
              reg417 <= ($signed($unsigned(reg416[(3'h6):(1'h1)])) ?
                  (reg406[(1'h1):(1'h0)] != ((reg290 + (wire277 <<< reg278)) << wire276[(4'hb):(1'h0)])) : reg412);
            end
          else
            begin
              reg415 <= (-reg291);
            end
        end
      else
        begin
          reg413 <= $unsigned(reg408);
        end
    end
  module418 modinst457 (wire456, clk, wire275, wire402, reg414, reg293, reg285);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module189
#( parameter param266 = (({(((8'had) ? (7'h41) : (8'hbd)) | (-(8'ha6)))} <<< (!((!(8'h9c)) ? (+(7'h40)) : ((8'hae) ? (8'hbd) : (8'h9c))))) ? ((((8'hac) & ((8'hb0) ? (8'ha5) : (8'hbd))) ? (8'ha3) : (&((8'ha8) ? (8'had) : (8'hab)))) ^ {(((8'hae) && (7'h42)) + {(8'hab), (8'hb6)}), ((~|(8'ha1)) >>> ((8'hb6) ? (8'ha4) : (8'hbe)))}) : (~^({{(8'ha1), (8'ha4)}} + (8'hb1)))) )
(y, clk, wire194, wire193, wire192, wire191, wire190);
  output wire [(32'h2e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire194;
  input wire [(4'ha):(1'h0)] wire193;
  input wire signed [(4'hd):(1'h0)] wire192;
  input wire [(4'hc):(1'h0)] wire191;
  input wire signed [(3'h7):(1'h0)] wire190;
  wire signed [(5'h12):(1'h0)] wire265;
  wire signed [(4'ha):(1'h0)] wire264;
  wire [(4'hb):(1'h0)] wire263;
  wire signed [(3'h6):(1'h0)] wire261;
  assign y = {wire265, wire264, wire263, wire261, (1'h0)};
  module195 modinst262 (wire261, clk, wire194, wire193, wire192, wire191);
  assign wire263 = (wire194 ?
                       $signed(wire194[(3'h5):(1'h1)]) : (wire193[(4'h8):(3'h7)] >>> (^~((wire194 ?
                               wire192 : (7'h42)) ?
                           $signed(wire194) : $signed(wire193)))));
  assign wire264 = ($unsigned($unsigned({wire192})) ?
                       (wire190 && (^$unsigned($unsigned(wire192)))) : $signed(wire193[(3'h6):(3'h6)]));
  assign wire265 = wire193;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module195
#( parameter param259 = (-((({(8'ha1)} <= ((8'hb4) ? (8'ha9) : (8'ha3))) ? ({(7'h43)} <<< (~|(7'h44))) : ({(8'ha4), (7'h41)} ? (^~(8'hae)) : ((8'ha6) != (8'ha9)))) ? ((((8'h9d) && (8'hb4)) << ((8'h9e) <<< (7'h41))) ? (((8'h9d) == (8'hab)) * ((7'h42) ? (8'hb0) : (8'hb4))) : (((8'h9d) == (8'hbc)) ? ((7'h44) ? (8'hac) : (7'h40)) : ((8'hbc) ? (8'h9e) : (8'ha5)))) : (^~(((8'ha5) ? (8'hae) : (8'hbc)) ? (-(8'hb6)) : ((8'hac) ? (8'hb7) : (8'hb7))))))
, parameter param260 = (-((8'ha8) ? (&(&(&param259))) : (((param259 ? param259 : (8'hbd)) ? (param259 ? param259 : param259) : (param259 ? param259 : param259)) ^ {(param259 ? param259 : param259)}))) )
(y, clk, wire199, wire198, wire197, wire196);
  output wire [(32'h2c2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire199;
  input wire [(2'h3):(1'h0)] wire198;
  input wire [(4'hd):(1'h0)] wire197;
  input wire signed [(3'h5):(1'h0)] wire196;
  wire [(4'ha):(1'h0)] wire258;
  wire signed [(2'h3):(1'h0)] wire257;
  wire [(3'h6):(1'h0)] wire256;
  wire [(4'h9):(1'h0)] wire255;
  wire [(2'h2):(1'h0)] wire254;
  wire signed [(5'h13):(1'h0)] wire253;
  reg signed [(4'h8):(1'h0)] reg252 = (1'h0);
  reg [(3'h6):(1'h0)] reg251 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg250 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg249 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg248 = (1'h0);
  reg [(3'h5):(1'h0)] reg247 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg246 = (1'h0);
  reg signed [(4'he):(1'h0)] reg245 = (1'h0);
  reg [(4'hf):(1'h0)] reg244 = (1'h0);
  reg [(4'he):(1'h0)] reg243 = (1'h0);
  reg signed [(4'he):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg241 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg240 = (1'h0);
  reg [(5'h11):(1'h0)] reg239 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg237 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg236 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg234 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg233 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg232 = (1'h0);
  reg [(4'h8):(1'h0)] reg231 = (1'h0);
  reg signed [(4'he):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg229 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg228 = (1'h0);
  reg [(3'h7):(1'h0)] reg227 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg226 = (1'h0);
  reg [(4'hb):(1'h0)] reg225 = (1'h0);
  wire [(5'h15):(1'h0)] wire224;
  wire signed [(3'h7):(1'h0)] wire223;
  reg signed [(5'h12):(1'h0)] reg222 = (1'h0);
  reg [(5'h12):(1'h0)] reg221 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg220 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg219 = (1'h0);
  reg [(5'h13):(1'h0)] reg218 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg217 = (1'h0);
  reg [(5'h15):(1'h0)] reg216 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg214 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg213 = (1'h0);
  wire [(5'h11):(1'h0)] wire212;
  wire signed [(4'hf):(1'h0)] wire211;
  wire [(5'h10):(1'h0)] wire210;
  wire [(3'h4):(1'h0)] wire209;
  wire signed [(5'h13):(1'h0)] wire208;
  wire signed [(3'h7):(1'h0)] wire207;
  wire signed [(4'hf):(1'h0)] wire206;
  wire signed [(3'h4):(1'h0)] wire205;
  wire [(4'h8):(1'h0)] wire204;
  wire signed [(5'h12):(1'h0)] wire203;
  wire signed [(5'h12):(1'h0)] wire202;
  wire [(3'h4):(1'h0)] wire201;
  wire [(5'h15):(1'h0)] wire200;
  assign y = {wire258,
                 wire257,
                 wire256,
                 wire255,
                 wire254,
                 wire253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 wire224,
                 wire223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 wire212,
                 wire211,
                 wire210,
                 wire209,
                 wire208,
                 wire207,
                 wire206,
                 wire205,
                 wire204,
                 wire203,
                 wire202,
                 wire201,
                 wire200,
                 (1'h0)};
  assign wire200 = wire196;
  assign wire201 = (8'hbc);
  assign wire202 = wire200[(4'he):(3'h6)];
  assign wire203 = ($unsigned($signed(wire198)) <<< ($unsigned(wire202) & wire196[(2'h3):(1'h1)]));
  assign wire204 = {$signed($unsigned(wire203[(5'h11):(4'h8)]))};
  assign wire205 = wire202[(3'h4):(1'h0)];
  assign wire206 = wire203[(2'h2):(1'h0)];
  assign wire207 = wire197[(4'hd):(4'h8)];
  assign wire208 = $signed({(|((!wire205) != $unsigned(wire199))),
                       (~&($signed(wire199) && $signed(wire201)))});
  assign wire209 = wire206[(3'h6):(1'h0)];
  assign wire210 = wire203[(4'hc):(1'h0)];
  assign wire211 = wire206;
  assign wire212 = $signed((wire211[(3'h6):(2'h2)] <= (-wire209)));
  always
    @(posedge clk) begin
      reg213 <= (|($signed((|wire196[(1'h0):(1'h0)])) + $unsigned(wire200[(3'h4):(1'h0)])));
      reg214 <= (($unsigned($signed((~&(8'hb4)))) << ((~&wire197[(4'hc):(3'h6)]) + $unsigned((wire205 + wire205)))) ?
          (wire210[(2'h3):(2'h2)] ?
              $unsigned(wire212[(4'he):(3'h6)]) : (&$unsigned((&wire199)))) : $unsigned($unsigned(wire202[(4'h9):(2'h2)])));
      if ({(8'hb2),
          ((!(reg213 ~^ $signed(wire205))) <<< (&(wire200 ^~ wire204[(3'h4):(1'h0)])))})
        begin
          if ($unsigned($signed($signed($signed((~^wire196))))))
            begin
              reg215 <= $unsigned($unsigned($signed($unsigned((wire202 ?
                  wire212 : (8'ha0))))));
              reg216 <= ((8'hb6) ?
                  $signed($signed($signed((wire207 ?
                      wire210 : wire204)))) : {(~&({wire199,
                          reg213} ~^ wire206)),
                      $signed(reg214)});
            end
          else
            begin
              reg215 <= $signed(($unsigned((reg214[(1'h0):(1'h0)] > (~^(8'hb7)))) ?
                  ({wire207, $unsigned(reg213)} ?
                      wire208 : (wire199 > reg215)) : $unsigned(wire201)));
              reg216 <= wire212[(3'h7):(1'h0)];
              reg217 <= (wire205[(2'h2):(1'h1)] && (wire198[(1'h0):(1'h0)] != reg213[(3'h4):(3'h4)]));
              reg218 <= (reg216[(2'h3):(2'h3)] && $unsigned({((reg217 >>> (8'ha4)) == (wire198 ?
                      wire199 : (8'hb9)))}));
              reg219 <= (wire210[(2'h2):(2'h2)] ?
                  $unsigned({(^{wire206})}) : reg217);
            end
        end
      else
        begin
          if ($signed(wire203))
            begin
              reg215 <= (-wire199[(2'h2):(1'h0)]);
            end
          else
            begin
              reg215 <= $signed($unsigned({$unsigned($signed(wire208)),
                  {{wire205, (8'h9e)}, wire207[(1'h0):(1'h0)]}}));
              reg216 <= reg215;
              reg217 <= $signed({reg219[(2'h2):(1'h1)],
                  wire199[(2'h3):(1'h0)]});
            end
          if ($signed((~|reg219[(2'h3):(1'h1)])))
            begin
              reg218 <= (~^($signed(((+wire201) || ((8'hbf) <<< reg218))) << $unsigned($signed((reg214 | (8'ha3))))));
              reg219 <= {(^~(wire197[(4'hd):(4'h8)] << $signed(wire203)))};
              reg220 <= (wire204[(3'h4):(2'h2)] ? $unsigned(reg217) : wire208);
              reg221 <= wire200[(5'h13):(4'hc)];
            end
          else
            begin
              reg218 <= wire207;
              reg219 <= $unsigned($unsigned((wire205[(3'h4):(1'h1)] ?
                  (^(wire200 && wire199)) : $unsigned(wire197))));
              reg220 <= (^~$unsigned((~(wire210[(1'h0):(1'h0)] ^ (reg218 & (8'ha7))))));
              reg221 <= (($unsigned(wire205) >= wire203) ?
                  reg220[(1'h1):(1'h0)] : wire206[(2'h3):(1'h1)]);
              reg222 <= (|$signed($signed({$unsigned((8'ha9))})));
            end
        end
    end
  assign wire223 = wire212;
  assign wire224 = $unsigned((wire203[(3'h4):(1'h0)] >>> ((wire204 && $signed(wire205)) ?
                       ((!reg222) ?
                           (reg221 >> wire207) : {wire223}) : $unsigned({wire196,
                           (7'h43)}))));
  always
    @(posedge clk) begin
      reg225 <= $unsigned(reg217);
      if (wire204[(2'h2):(2'h2)])
        begin
          if ({$signed(reg214)})
            begin
              reg226 <= (wire201 ?
                  wire204[(3'h6):(1'h0)] : $signed($unsigned($unsigned(wire223))));
            end
          else
            begin
              reg226 <= (~{(-(reg213 ? wire212[(5'h11):(4'hb)] : (+reg215))),
                  $signed(reg213[(2'h2):(2'h2)])});
              reg227 <= {$unsigned({reg219,
                      ((wire202 ? (8'hb4) : reg226) ?
                          (~^wire199) : $signed(reg215))}),
                  wire211};
            end
          reg228 <= ((+((wire201 ? reg222[(3'h7):(1'h1)] : reg225) ?
                  {$unsigned((8'h9e)), (wire199 < wire202)} : ((^wire206) ?
                      (~|(7'h42)) : wire200[(5'h13):(1'h1)]))) ?
              $unsigned((!$signed((wire208 ?
                  reg217 : wire202)))) : $signed($unsigned(((~^wire199) ?
                  reg221[(4'hf):(3'h6)] : $signed(reg218)))));
          if ((reg227[(3'h4):(3'h4)] ~^ (((|{wire208, wire207}) ?
                  {$unsigned(reg227), reg222[(2'h3):(1'h0)]} : {(reg213 ?
                          (8'hba) : wire210)}) ?
              wire203[(4'hc):(4'ha)] : reg213[(3'h6):(1'h0)])))
            begin
              reg229 <= reg222[(5'h12):(4'hf)];
            end
          else
            begin
              reg229 <= $signed((reg217[(3'h5):(1'h1)] ?
                  reg219 : {$signed($signed(wire210)), reg226}));
              reg230 <= wire205[(2'h3):(1'h1)];
              reg231 <= $signed((-reg218));
            end
          if ($signed($unsigned((|$unsigned((-(8'hbd)))))))
            begin
              reg232 <= $unsigned((~^(~|wire211)));
            end
          else
            begin
              reg232 <= ({(&$signed(reg220)), reg213} <= wire212);
              reg233 <= $unsigned(({$signed({(7'h43), wire224})} ?
                  (8'hbc) : ($unsigned((^wire197)) ?
                      ((reg231 >> reg219) || (reg217 >>> wire206)) : ((wire208 ^ wire224) != (reg216 ?
                          (8'ha6) : wire201)))));
              reg234 <= $unsigned(({reg216,
                  $unsigned({wire208})} << (((wire207 ^~ reg228) ^~ {wire198,
                      wire206}) ?
                  (wire208 & (wire203 >>> wire197)) : wire200)));
              reg235 <= $signed(($unsigned((&wire198)) ?
                  reg220 : $unsigned(($unsigned((8'hba)) ?
                      $signed(reg219) : (~|wire196)))));
            end
          if ((($signed(wire209) ?
              ((wire201 ?
                  reg227[(3'h7):(3'h6)] : (|wire198)) != reg233[(3'h4):(1'h1)]) : wire199) >= $signed(({(^wire209)} ?
              ($unsigned((8'ha5)) || (~|reg226)) : (reg217[(1'h0):(1'h0)] ?
                  {(8'hb7), reg232} : wire198[(1'h0):(1'h0)])))))
            begin
              reg236 <= reg229[(5'h10):(4'hc)];
              reg237 <= (|((wire207[(2'h3):(2'h3)] | (-(^~(8'ha9)))) ?
                  wire210 : wire204[(3'h4):(2'h2)]));
              reg238 <= {($unsigned($signed($signed(reg231))) ^~ $unsigned((^$unsigned(wire203)))),
                  ((reg232[(2'h3):(2'h3)] * reg220[(4'hf):(4'hd)]) ?
                      {(8'h9c)} : reg220[(4'hb):(4'hb)])};
              reg239 <= wire210[(2'h3):(1'h0)];
            end
          else
            begin
              reg236 <= $unsigned($unsigned($unsigned($unsigned(reg213[(4'h8):(2'h3)]))));
            end
        end
      else
        begin
          if (wire212[(2'h3):(1'h0)])
            begin
              reg226 <= reg222[(4'h8):(3'h5)];
              reg227 <= (8'h9d);
              reg228 <= $signed((~|$unsigned((!$unsigned(reg237)))));
              reg229 <= {reg227[(2'h3):(1'h1)]};
              reg230 <= $unsigned(reg226);
            end
          else
            begin
              reg226 <= (wire197 + (|{wire199[(2'h2):(2'h2)],
                  {(!wire199), (wire208 || reg229)}}));
            end
          if ((^~(+(~|wire207))))
            begin
              reg231 <= (reg221[(4'h8):(2'h3)] ?
                  wire199 : ((({(8'h9c), wire200} > ((8'hb1) ?
                          wire208 : wire212)) ?
                      (wire205[(3'h4):(3'h4)] << wire201[(1'h0):(1'h0)]) : reg233) + reg231));
              reg232 <= (!$signed((-reg237)));
              reg233 <= reg233[(3'h5):(3'h5)];
            end
          else
            begin
              reg231 <= $signed(({$signed(wire208), $signed((!reg234))} ?
                  wire209[(1'h1):(1'h1)] : ((reg215[(1'h0):(1'h0)] ~^ $unsigned(wire208)) ?
                      ($signed(reg218) & $signed(wire201)) : $signed({wire199}))));
              reg232 <= {$signed(($signed(reg226) | wire211[(2'h3):(1'h0)])),
                  (wire205 >= {{$unsigned(reg216)},
                      $unsigned($unsigned(wire203))})};
              reg233 <= ($signed({wire199,
                  $unsigned((reg222 ?
                      wire202 : wire203))}) <<< $unsigned($unsigned((reg215[(3'h6):(3'h5)] ?
                  wire224 : $signed(wire203)))));
              reg234 <= ($unsigned((reg220[(2'h3):(1'h0)] ?
                  $unsigned(wire199) : wire197[(4'ha):(3'h4)])) || (+{$signed(wire209)}));
              reg235 <= ({(|(~^(wire201 <= wire196))),
                  $unsigned(reg218[(3'h7):(3'h4)])} ^~ wire203);
            end
          reg236 <= ((reg234[(3'h6):(3'h5)] == $unsigned(wire223)) && reg216[(4'he):(3'h5)]);
        end
      if (($signed({reg232,
          (((8'hb3) <= (8'hbc)) * $signed(wire200))}) != (reg217 && $signed((&reg233)))))
        begin
          if ({wire200})
            begin
              reg240 <= $unsigned(wire223[(3'h6):(1'h1)]);
            end
          else
            begin
              reg240 <= (reg218[(4'ha):(4'h9)] ?
                  $signed((reg214 < wire200[(1'h0):(1'h0)])) : wire223[(3'h6):(3'h4)]);
              reg241 <= {$signed((^~reg225[(3'h4):(2'h3)]))};
            end
          if ((&(($signed($signed(wire198)) ?
              $signed((!reg214)) : reg225[(4'h8):(1'h1)]) != ((~&(reg239 ~^ (8'haa))) ?
              ((reg227 ^ reg238) | $signed((7'h41))) : ($unsigned(reg220) ?
                  wire202[(4'hd):(3'h6)] : ((7'h44) & reg217))))))
            begin
              reg242 <= $signed($signed(wire210[(1'h1):(1'h1)]));
              reg243 <= $unsigned($unsigned($unsigned((~&(-reg217)))));
              reg244 <= $signed((&wire207));
            end
          else
            begin
              reg242 <= (wire207[(3'h7):(3'h6)] || $signed(wire204[(4'h8):(3'h7)]));
              reg243 <= (reg237[(4'hd):(2'h3)] + (8'hbe));
              reg244 <= {reg221};
              reg245 <= (|reg239);
              reg246 <= reg229[(2'h2):(1'h1)];
            end
          if (($unsigned({($signed(reg241) && $unsigned(reg218))}) ?
              reg233 : {{((^reg225) ? {(8'hb8)} : reg225),
                      ((reg242 ? reg215 : reg246) | (reg220 ?
                          reg214 : (8'hbd)))},
                  reg243}))
            begin
              reg247 <= ($unsigned(($signed((wire200 ?
                  reg213 : reg241)) && {(reg237 ?
                      wire196 : reg246)})) <= (^reg222));
              reg248 <= $signed(reg228[(1'h0):(1'h0)]);
              reg249 <= ($unsigned({((~|reg228) | $unsigned((8'hb9))),
                  reg222[(1'h0):(1'h0)]}) <= reg221);
            end
          else
            begin
              reg247 <= ($signed(($signed((reg234 ?
                  wire212 : wire207)) ^ $unsigned(reg248[(5'h10):(1'h1)]))) << $signed($unsigned({(~|reg247),
                  $signed(wire207)})));
            end
          reg250 <= (reg241[(3'h4):(1'h0)] & $unsigned($signed(($unsigned(wire199) < (-reg233)))));
          reg251 <= wire203[(3'h5):(3'h5)];
        end
      else
        begin
          if ($unsigned($unsigned((8'ha9))))
            begin
              reg240 <= ($signed($unsigned((reg214 ?
                      reg243[(3'h7):(3'h5)] : {reg222}))) ?
                  ((({reg229, reg250} ?
                          ((8'hbe) ? reg217 : (8'hab)) : (wire201 ?
                              reg249 : reg218)) ?
                      ((&(8'hbe)) > {reg251}) : ((reg214 ? reg229 : reg230) ?
                          $unsigned(wire196) : (wire205 | reg240))) & $signed(((reg229 || (8'ha8)) <<< reg219[(1'h0):(1'h0)]))) : $unsigned((~^$signed(reg240[(3'h6):(2'h3)]))));
            end
          else
            begin
              reg240 <= wire196[(1'h1):(1'h1)];
              reg241 <= ($unsigned(($signed((reg235 ?
                  reg216 : reg217)) ~^ wire199)) - $signed(($signed({reg225}) ?
                  (^(reg228 >> (8'hbb))) : reg219[(1'h0):(1'h0)])));
            end
          reg242 <= wire224;
          reg243 <= ($unsigned(reg231) ?
              $unsigned(reg216) : wire204[(3'h4):(2'h2)]);
        end
      reg252 <= ($unsigned((((reg225 ? (7'h44) : reg213) ?
                  (reg234 ? reg220 : reg247) : (8'hae)) ?
              $signed((^~wire198)) : $signed($unsigned(reg218)))) ?
          (^wire197) : (8'hac));
    end
  assign wire253 = $unsigned(($signed(wire208) <= $unsigned(($signed(reg240) ?
                       (reg240 ? wire224 : reg237) : {wire202}))));
  assign wire254 = {((reg218 ?
                           $signed(reg244) : (^~reg229)) ~^ $unsigned((!$unsigned((8'ha9))))),
                       (reg220 ?
                           ($unsigned({reg227}) ?
                               (8'ha2) : wire253[(3'h4):(2'h3)]) : (wire253[(1'h0):(1'h0)] >= (8'h9d)))};
  assign wire255 = wire202[(1'h0):(1'h0)];
  assign wire256 = ($signed($signed(reg222)) ?
                       (^~$signed(wire223)) : (-{($unsigned(wire203) & wire206)}));
  assign wire257 = (wire254[(1'h0):(1'h0)] ?
                       reg215[(1'h1):(1'h1)] : ($signed((^{wire207})) >>> $signed(((8'ha4) && wire212))));
  assign wire258 = ($signed((((8'ha5) >>> ((8'ha7) ^~ reg219)) >> ((reg217 >>> reg230) ?
                       (+reg236) : reg244))) > (reg221 <<< reg245[(1'h0):(1'h0)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module418
#( parameter param454 = (((((~|(7'h44)) ? ((8'hb0) != (7'h42)) : ((8'ha1) ? (8'ha3) : (8'ha6))) || ({(8'hb0), (8'hbd)} ~^ ((8'hb6) & (8'hb2)))) - ((((8'hb4) >>> (8'hbe)) ? ((8'h9f) <= (8'hae)) : (~^(8'ha4))) >= (|((8'haf) * (8'hac))))) ? (-{(((8'ha9) ? (7'h42) : (8'hb6)) << ((8'ha3) <= (8'ha4)))}) : ((~({(8'ha3)} || ((8'had) << (8'h9e)))) >>> ((|((8'ha1) * (8'ha3))) == (((7'h41) ? (8'hb9) : (8'ha4)) > ((8'h9f) ~^ (8'ha3))))))
, parameter param455 = ((((!{param454, param454}) ~^ (param454 ? (param454 <<< (8'ha9)) : (~|param454))) & (((8'hbd) < (param454 ? param454 : param454)) ~^ (-param454))) >> (!(8'hb3))) )
(y, clk, wire423, wire422, wire421, wire420, wire419);
  output wire [(32'h128):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire423;
  input wire [(4'hc):(1'h0)] wire422;
  input wire [(5'h12):(1'h0)] wire421;
  input wire [(4'ha):(1'h0)] wire420;
  input wire [(5'h12):(1'h0)] wire419;
  reg [(2'h2):(1'h0)] reg453 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg452 = (1'h0);
  reg [(4'ha):(1'h0)] reg451 = (1'h0);
  reg [(3'h6):(1'h0)] reg450 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg449 = (1'h0);
  reg [(4'hb):(1'h0)] reg448 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg447 = (1'h0);
  reg [(3'h5):(1'h0)] reg446 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg445 = (1'h0);
  reg signed [(4'he):(1'h0)] reg444 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg443 = (1'h0);
  reg [(4'hc):(1'h0)] reg442 = (1'h0);
  reg [(5'h14):(1'h0)] reg441 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg440 = (1'h0);
  reg [(3'h5):(1'h0)] reg439 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg438 = (1'h0);
  reg [(3'h5):(1'h0)] reg437 = (1'h0);
  reg [(2'h2):(1'h0)] reg436 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg435 = (1'h0);
  wire [(4'hc):(1'h0)] wire434;
  reg signed [(5'h13):(1'h0)] reg433 = (1'h0);
  reg signed [(4'he):(1'h0)] reg432 = (1'h0);
  reg [(2'h3):(1'h0)] reg431 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire430;
  wire signed [(4'hb):(1'h0)] wire429;
  wire [(4'ha):(1'h0)] wire428;
  wire signed [(3'h7):(1'h0)] wire427;
  wire [(4'h9):(1'h0)] wire426;
  wire [(4'hb):(1'h0)] wire425;
  wire [(5'h10):(1'h0)] wire424;
  assign y = {reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 reg447,
                 reg446,
                 reg445,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 wire434,
                 reg433,
                 reg432,
                 reg431,
                 wire430,
                 wire429,
                 wire428,
                 wire427,
                 wire426,
                 wire425,
                 wire424,
                 (1'h0)};
  assign wire424 = (($unsigned($signed((wire420 ?
                       (8'had) : wire421))) && $unsigned($unsigned({wire422,
                       wire419}))) >>> (wire423 || $signed(wire422[(4'hb):(3'h5)])));
  assign wire425 = wire420[(4'h8):(3'h4)];
  assign wire426 = wire419[(3'h6):(1'h0)];
  assign wire427 = $signed({($unsigned(wire419) ?
                           wire426[(4'h8):(2'h3)] : $signed((8'had)))});
  assign wire428 = (wire426 ?
                       (wire427 ?
                           ((|(wire423 ? wire427 : wire422)) ?
                               (8'hb8) : (8'ha1)) : ($signed(wire426[(3'h7):(1'h1)]) ?
                               ($unsigned((8'ha3)) ^ (+wire421)) : $signed((wire426 <<< wire420)))) : (wire426 ^~ ({$unsigned(wire420),
                               $unsigned(wire424)} ?
                           $unsigned($unsigned(wire423)) : (|$signed(wire419)))));
  assign wire429 = (~&((wire426[(2'h2):(2'h2)] ~^ $unsigned((wire419 ?
                           wire427 : wire424))) ?
                       wire424 : (wire425[(4'ha):(4'ha)] ?
                           (((8'h9d) ? wire422 : wire426) ?
                               wire427 : (wire423 ^~ wire423)) : wire427)));
  assign wire430 = {$signed((~|(^wire429))),
                       ({$signed((wire425 ? (8'ha8) : wire422))} ?
                           (({wire425, wire423} ?
                                   $signed((8'ha4)) : ((8'hb1) != wire426)) ?
                               (wire423[(3'h4):(2'h2)] ?
                                   (wire424 ^ wire429) : wire423) : $unsigned(wire419)) : {((wire420 != wire428) ^~ {wire425})})};
  always
    @(posedge clk) begin
      if ($signed(wire425))
        begin
          reg431 <= (~&wire429);
        end
      else
        begin
          reg431 <= $signed((&reg431[(1'h1):(1'h0)]));
        end
      reg432 <= (~(^(~|($signed(wire420) ? (8'hbb) : (!wire425)))));
      reg433 <= wire430;
    end
  assign wire434 = (($signed(({wire420} != (wire419 ?
                           wire428 : wire424))) >> ((8'ha8) ?
                           $unsigned($unsigned(reg432)) : $unsigned((reg433 ?
                               wire427 : reg432)))) ?
                       ($signed($unsigned($signed(wire421))) ?
                           $unsigned(wire420) : $unsigned(wire428[(4'ha):(3'h6)])) : wire420);
  always
    @(posedge clk) begin
      if (wire427)
        begin
          reg435 <= wire423[(3'h4):(3'h4)];
          if ($unsigned((&$signed($signed(reg432[(1'h1):(1'h1)])))))
            begin
              reg436 <= (wire419 ?
                  $unsigned($unsigned((+$signed(wire426)))) : wire420[(2'h2):(1'h1)]);
            end
          else
            begin
              reg436 <= $unsigned(($unsigned(wire419) ?
                  $signed((wire424 ?
                      $signed(wire434) : ((8'ha8) == wire434))) : $signed(((wire423 ?
                          wire420 : (8'hb5)) ?
                      (wire423 >>> (8'ha2)) : $signed(wire421)))));
              reg437 <= wire427[(3'h4):(3'h4)];
              reg438 <= wire421[(4'h9):(2'h3)];
            end
          reg439 <= $signed($unsigned(($unsigned((|reg435)) && $unsigned($signed((7'h41))))));
          if ($signed((($unsigned({reg435, reg439}) ?
                  (((8'hb6) > reg438) ?
                      wire426[(2'h3):(2'h2)] : (~^wire434)) : (~|wire428)) ?
              $unsigned(((reg439 > wire424) < {wire425})) : $signed((8'hab)))))
            begin
              reg440 <= (wire428 >> reg435);
              reg441 <= $signed((8'ha2));
              reg442 <= {$signed(($signed(wire434) * $unsigned((~^wire430)))),
                  (({wire428[(3'h7):(2'h3)]} <<< reg437[(1'h0):(1'h0)]) ^ ($unsigned(((8'ha6) ?
                      wire428 : reg437)) ^~ (~^{reg439, wire428})))};
              reg443 <= (reg442[(3'h4):(3'h4)] ?
                  $unsigned($unsigned({(~&wire425)})) : wire428[(3'h6):(3'h6)]);
            end
          else
            begin
              reg440 <= {((wire420 == ((wire434 ~^ wire425) & {wire425})) ?
                      ({wire422, $unsigned((8'hac))} == (~&reg443)) : (8'hb0))};
              reg441 <= wire421;
              reg442 <= (reg438 >>> reg437[(2'h2):(1'h0)]);
              reg443 <= wire423;
              reg444 <= $unsigned({($unsigned(reg443) + $signed($signed(reg432)))});
            end
          if (wire430[(2'h3):(2'h3)])
            begin
              reg445 <= $unsigned($unsigned(wire434));
            end
          else
            begin
              reg445 <= (|{(((reg436 ?
                      wire423 : wire426) ^ $unsigned((8'hb5))) & reg442),
                  ($signed(wire421) ?
                      (reg433[(1'h0):(1'h0)] | $unsigned(reg433)) : reg439[(2'h2):(1'h1)])});
              reg446 <= $signed($signed(reg443));
              reg447 <= (wire427 != (~|$signed(reg437)));
              reg448 <= (~&wire428);
              reg449 <= reg433[(4'h8):(1'h0)];
            end
        end
      else
        begin
          reg435 <= $unsigned(((8'hb5) & reg436[(2'h2):(2'h2)]));
        end
      reg450 <= $unsigned((~|($signed($signed(reg432)) ~^ $signed(wire430[(3'h6):(3'h5)]))));
      reg451 <= {$signed((reg440[(2'h2):(2'h2)] ?
              $signed($unsigned(reg438)) : {((7'h41) ? reg449 : reg439),
                  $signed(reg446)}))};
      reg452 <= $signed((({{(8'had), reg438},
              (wire430 >>> wire428)} + $unsigned(reg436[(1'h1):(1'h0)])) ?
          wire419 : (($signed(reg442) ?
              (|wire421) : {reg448}) ^~ wire427[(3'h5):(1'h1)])));
      reg453 <= {{(-((^~reg445) ? $unsigned(wire420) : wire419))}};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module330
#( parameter param395 = (((~&(|((8'hbf) ? (8'ha4) : (8'haa)))) ? (~((~|(8'hb0)) ? ((8'ha3) ? (8'hb7) : (8'ha6)) : ((7'h41) ? (8'hb2) : (8'ha8)))) : {{((8'hb5) ? (8'hba) : (8'hb8))}}) != (({((8'hb2) ^ (8'hac))} ^~ (~&((7'h43) * (8'hbb)))) ? (+(((8'hba) ? (8'hbd) : (8'hbf)) ^ ((8'h9f) ? (8'h9e) : (8'ha3)))) : (&(((8'hb1) ? (8'ha3) : (8'h9c)) > ((8'hbe) ? (7'h44) : (8'ha5))))))
, parameter param396 = ((7'h43) >= (^~(((+param395) ? {param395, param395} : (~&param395)) ? {(param395 > param395), (param395 ^ param395)} : (&(^~param395))))) )
(y, clk, wire335, wire334, wire333, wire332, wire331);
  output wire [(32'h29f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire335;
  input wire signed [(2'h3):(1'h0)] wire334;
  input wire [(3'h5):(1'h0)] wire333;
  input wire [(4'hf):(1'h0)] wire332;
  input wire signed [(4'he):(1'h0)] wire331;
  wire [(5'h12):(1'h0)] wire394;
  reg [(4'hd):(1'h0)] reg393 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg392 = (1'h0);
  reg [(2'h2):(1'h0)] reg391 = (1'h0);
  reg [(4'hc):(1'h0)] reg390 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg389 = (1'h0);
  reg [(4'ha):(1'h0)] reg388 = (1'h0);
  reg [(2'h2):(1'h0)] reg387 = (1'h0);
  reg [(5'h12):(1'h0)] reg386 = (1'h0);
  reg [(3'h7):(1'h0)] reg385 = (1'h0);
  reg [(3'h5):(1'h0)] reg384 = (1'h0);
  reg [(2'h3):(1'h0)] reg383 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg382 = (1'h0);
  reg [(4'hf):(1'h0)] reg381 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg380 = (1'h0);
  reg [(5'h13):(1'h0)] reg379 = (1'h0);
  reg [(4'ha):(1'h0)] reg378 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg377 = (1'h0);
  reg [(5'h10):(1'h0)] reg376 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg375 = (1'h0);
  reg [(5'h11):(1'h0)] reg374 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg373 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg372 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg370 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire369;
  wire signed [(3'h5):(1'h0)] wire368;
  wire [(5'h14):(1'h0)] wire367;
  wire [(2'h3):(1'h0)] wire366;
  wire signed [(3'h4):(1'h0)] wire365;
  wire signed [(5'h10):(1'h0)] wire364;
  wire signed [(5'h11):(1'h0)] wire363;
  reg signed [(3'h6):(1'h0)] reg362 = (1'h0);
  reg [(5'h13):(1'h0)] reg361 = (1'h0);
  reg [(3'h7):(1'h0)] reg360 = (1'h0);
  reg [(4'hf):(1'h0)] reg359 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg358 = (1'h0);
  reg [(2'h3):(1'h0)] reg357 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg356 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg355 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg354 = (1'h0);
  reg signed [(4'he):(1'h0)] reg353 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg352 = (1'h0);
  wire [(5'h14):(1'h0)] wire351;
  reg signed [(3'h7):(1'h0)] reg350 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg349 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg348 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg347 = (1'h0);
  reg [(4'hf):(1'h0)] reg346 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg345 = (1'h0);
  reg [(3'h6):(1'h0)] reg344 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg342 = (1'h0);
  reg [(5'h13):(1'h0)] reg341 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg340 = (1'h0);
  reg signed [(4'he):(1'h0)] reg339 = (1'h0);
  reg [(5'h15):(1'h0)] reg338 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg337 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire336;
  assign y = {wire394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 wire369,
                 wire368,
                 wire367,
                 wire366,
                 wire365,
                 wire364,
                 wire363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 wire351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 wire336,
                 (1'h0)};
  assign wire336 = $signed($unsigned($signed($signed((wire334 ?
                       wire335 : wire333)))));
  always
    @(posedge clk) begin
      reg337 <= ($unsigned($unsigned((&$unsigned(wire335)))) ?
          (^~wire336[(3'h7):(3'h4)]) : wire335);
      if ($signed({(+{$unsigned(wire331)})}))
        begin
          if (((!wire333) << (~$signed($unsigned({wire331, (8'h9f)})))))
            begin
              reg338 <= reg337;
              reg339 <= (wire334[(2'h2):(1'h1)] ?
                  reg338[(5'h15):(3'h4)] : $signed({{$unsigned((8'ha8))},
                      (reg337 ^~ wire332[(4'hc):(2'h2)])}));
              reg340 <= {(^~$signed((~^((8'hac) ? wire333 : reg338))))};
              reg341 <= (reg339[(4'ha):(2'h2)] - $unsigned({((wire336 ?
                      wire334 : (8'h9f)) <<< $unsigned(wire332)),
                  ($unsigned((8'hab)) && $signed(wire331))}));
            end
          else
            begin
              reg338 <= $signed((($unsigned($unsigned(reg338)) >>> wire334) ?
                  reg337 : {(wire336 ? (~|reg339) : reg340[(3'h5):(2'h3)])}));
            end
          reg342 <= $unsigned(wire333);
        end
      else
        begin
          reg338 <= $unsigned(reg338);
        end
      if ($signed(($unsigned(($unsigned(reg340) != reg337[(3'h6):(1'h1)])) ?
          (~&($unsigned(reg341) ?
              (wire336 < (8'ha2)) : $unsigned((8'h9d)))) : ((8'h9f) ^~ $unsigned((~wire331))))))
        begin
          reg343 <= wire331;
          reg344 <= ((~wire332) ?
              (&(wire333[(1'h0):(1'h0)] ^ $signed($unsigned(wire335)))) : ((&((reg337 ?
                      wire332 : wire335) | (+reg338))) ?
                  $signed($signed($unsigned((8'hbb)))) : {(+((8'h9c) & wire334))}));
          reg345 <= $unsigned(reg337[(3'h4):(2'h3)]);
        end
      else
        begin
          if ($unsigned({(reg344[(1'h1):(1'h1)] | (8'hbe)), wire331}))
            begin
              reg343 <= (8'hac);
              reg344 <= {wire331[(4'hc):(3'h7)], reg339[(3'h5):(3'h5)]};
              reg345 <= ({(~^(reg341[(4'hf):(2'h3)] ^ $unsigned(reg344))),
                  {wire333}} >>> (8'hab));
              reg346 <= (^~(~|$signed((wire335[(4'hb):(3'h6)] == (reg340 >>> (8'hb6))))));
            end
          else
            begin
              reg343 <= (wire332[(3'h4):(1'h0)] ?
                  ((reg341 ?
                      reg339[(1'h0):(1'h0)] : (~(wire334 ?
                          wire336 : wire332))) ^~ reg337) : (reg337[(3'h6):(2'h2)] <<< {(-$signed(reg342))}));
              reg344 <= $unsigned(reg337);
              reg345 <= (&$signed(({(reg337 ? reg342 : (8'hba)),
                  $unsigned(wire335)} == ($unsigned((8'ha6)) != $unsigned(reg343)))));
              reg346 <= reg342[(4'h9):(3'h6)];
              reg347 <= (~^{$signed((&(wire331 && reg337))),
                  $unsigned(($signed(wire335) ^ (wire336 ?
                      wire334 : reg344)))});
            end
          reg348 <= ((8'hb5) ?
              {((~|{wire335}) <<< (wire335[(5'h13):(5'h11)] << $unsigned(reg346))),
                  $unsigned((reg344[(3'h4):(2'h3)] <= reg345))} : (reg347[(4'hf):(1'h1)] >= reg340[(3'h5):(2'h3)]));
        end
      reg349 <= (8'hb2);
      reg350 <= (reg341[(3'h7):(2'h3)] <<< reg343);
    end
  assign wire351 = (((8'hbb) ?
                       (($signed(reg345) ? $unsigned(reg349) : reg348) ?
                           $unsigned($signed(wire333)) : {(wire334 - reg349)}) : (reg340[(4'h9):(4'h8)] ?
                           (8'ha5) : ($unsigned(reg344) ?
                               (~&reg340) : $signed((8'hbe))))) - $unsigned((wire336 ^ ((&reg343) >>> (reg343 ?
                       wire332 : reg349)))));
  always
    @(posedge clk) begin
      if (reg349[(2'h2):(2'h2)])
        begin
          if ((8'had))
            begin
              reg352 <= (reg349 ?
                  (+(7'h44)) : {((8'hb2) <<< $unsigned({wire334}))});
              reg353 <= wire351[(5'h13):(5'h12)];
              reg354 <= (^(($signed((~&(8'ha4))) ?
                  ($signed((8'hb5)) ?
                      (reg352 & reg343) : $signed(reg340)) : $signed($signed(reg349))) <<< (^(wire351 ?
                  ((8'had) ? wire334 : reg347) : $unsigned(reg338)))));
            end
          else
            begin
              reg352 <= $signed({{$unsigned((reg340 < wire331)),
                      ($signed(reg352) ^ (wire336 || reg347))}});
              reg353 <= $unsigned((^$unsigned($signed((^~reg354)))));
              reg354 <= ((reg337[(1'h0):(1'h0)] > {{$unsigned(wire336),
                          (&reg344)},
                      (wire335[(3'h6):(2'h2)] ?
                          {reg353, (8'ha0)} : (wire334 > (8'hbe)))}) ?
                  $signed($unsigned(((&reg338) | $signed(reg348)))) : (($signed($unsigned(reg345)) * (reg353[(1'h1):(1'h0)] & reg340[(2'h3):(1'h0)])) <<< (reg344 & $unsigned($signed(wire351)))));
              reg355 <= $signed(reg354[(5'h12):(4'hf)]);
              reg356 <= reg346;
            end
          reg357 <= ($signed((($unsigned(wire332) ?
                  reg341[(4'ha):(1'h0)] : $unsigned(reg354)) ?
              reg352[(3'h6):(3'h6)] : $signed((reg355 ?
                  wire331 : reg346)))) * ($unsigned(((~reg356) ?
              $unsigned(reg341) : $signed(wire336))) ~^ reg350));
          if (reg339)
            begin
              reg358 <= (((~^wire331[(2'h3):(2'h3)]) ?
                  (8'hba) : (({reg346, (8'hb3)} ?
                      (wire335 ?
                          reg356 : wire332) : $unsigned(wire336)) + wire331)) < $unsigned(($signed((reg347 ?
                  wire351 : wire334)) != reg339)));
              reg359 <= (~|($unsigned(reg348[(2'h2):(1'h0)]) ?
                  $unsigned((8'ha6)) : $signed(($unsigned(reg340) >> (reg358 ?
                      wire332 : wire336)))));
            end
          else
            begin
              reg358 <= reg343;
              reg359 <= (wire333 > reg342);
              reg360 <= reg344;
            end
        end
      else
        begin
          if (($unsigned(reg348[(1'h1):(1'h0)]) << $unsigned((~&(^~$unsigned(reg337))))))
            begin
              reg352 <= reg338;
            end
          else
            begin
              reg352 <= (7'h44);
              reg353 <= reg354;
              reg354 <= (!reg352[(4'ha):(2'h3)]);
              reg355 <= $signed(((~^reg355[(2'h3):(2'h3)]) ?
                  (&$signed(reg350[(1'h0):(1'h0)])) : {($signed(wire334) <<< (reg357 ?
                          reg355 : reg358)),
                      reg358}));
            end
          reg356 <= {$unsigned((^~wire336[(1'h1):(1'h1)])),
              reg348[(1'h0):(1'h0)]};
          reg357 <= reg357;
          reg358 <= $signed((wire332[(3'h5):(2'h2)] ?
              reg337[(3'h5):(1'h0)] : $signed($unsigned(reg354[(5'h14):(2'h2)]))));
          reg359 <= $signed({(~&($signed(reg354) ?
                  {reg339, (8'hba)} : $signed(reg355))),
              (+reg337[(5'h10):(5'h10)])});
        end
      reg361 <= $unsigned(reg339);
      reg362 <= $unsigned($signed(((~^{(7'h43)}) < reg343)));
    end
  assign wire363 = (~&(8'ha7));
  assign wire364 = {wire335, $signed((~^reg354))};
  assign wire365 = reg348;
  assign wire366 = $unsigned((^$unsigned(reg338)));
  assign wire367 = wire334;
  assign wire368 = ($unsigned(wire351[(3'h6):(3'h6)]) ?
                       reg362[(2'h3):(2'h3)] : {((^~(reg358 ?
                                   wire335 : reg339)) ?
                               ((~&wire333) ?
                                   reg360[(3'h6):(1'h0)] : $unsigned(reg338)) : wire365[(2'h2):(2'h2)])});
  assign wire369 = $unsigned($unsigned(($signed({reg346}) > (reg342[(4'hd):(3'h7)] ?
                       reg348 : $unsigned((8'hbb))))));
  always
    @(posedge clk) begin
      if (reg362[(1'h0):(1'h0)])
        begin
          reg370 <= $signed($signed(wire368[(2'h3):(2'h3)]));
        end
      else
        begin
          reg370 <= (reg359[(4'hc):(1'h0)] ?
              ($unsigned((reg360 << (^~reg360))) ?
                  ((+reg338[(3'h5):(3'h4)]) < ($unsigned(reg350) ?
                      (reg340 <= wire351) : $unsigned(reg343))) : reg361[(2'h3):(2'h2)]) : ((((reg337 ?
                          reg353 : reg360) >= (reg344 ? reg339 : reg342)) ?
                      $signed({wire366}) : $unsigned((^reg359))) ?
                  (!(!(~^reg370))) : (($signed(wire335) <= $signed(reg359)) + (~&(-wire351)))));
          reg371 <= wire369[(2'h3):(2'h2)];
          reg372 <= $signed((|$unsigned(((8'hab) >>> (wire351 ?
              reg343 : reg341)))));
        end
      reg373 <= (reg358[(4'ha):(2'h2)] ?
          $unsigned($signed(($unsigned(wire332) ?
              (reg347 ? wire351 : wire367) : $signed(wire332)))) : wire332);
      reg374 <= (+wire366[(2'h2):(1'h1)]);
      if ($signed((|reg354[(4'hf):(3'h5)])))
        begin
          if (reg342[(4'h8):(1'h0)])
            begin
              reg375 <= ($unsigned($signed((&reg342))) > wire333);
              reg376 <= ({(8'ha4)} ?
                  $signed($signed(((-wire351) ?
                      $signed(wire351) : (reg372 * reg348)))) : ({$signed((reg341 | (8'hb0))),
                          $signed($unsigned(reg355))} ?
                      $unsigned(reg360) : $unsigned(reg359[(3'h6):(3'h6)])));
              reg377 <= (!$signed((~|(|(~&reg349)))));
            end
          else
            begin
              reg375 <= ({{(-$signed(wire363))}} >= $signed(wire367[(5'h13):(2'h2)]));
            end
          if (wire363)
            begin
              reg378 <= {(|reg348[(1'h1):(1'h1)]), reg353[(3'h4):(2'h3)]};
              reg379 <= $signed(reg344[(2'h2):(1'h1)]);
              reg380 <= ($unsigned({($signed(reg374) ?
                      reg362 : $signed(reg356))}) | ((reg350[(3'h5):(2'h2)] && $signed((wire336 ?
                  reg354 : wire368))) == reg347[(4'he):(4'h9)]));
              reg381 <= (($unsigned(((^(7'h41)) ? (~^wire351) : {reg376})) ?
                      $unsigned(wire351) : {(((8'haa) ? reg352 : wire369) ?
                              (reg361 >= reg340) : (reg338 ?
                                  (8'haf) : reg350))}) ?
                  ($unsigned($signed(reg360)) ?
                      $signed({(reg353 > wire369)}) : $unsigned($signed((~reg360)))) : reg379[(4'h9):(4'h8)]);
              reg382 <= wire367;
            end
          else
            begin
              reg378 <= $unsigned((reg373[(1'h1):(1'h1)] ?
                  (~&{reg362}) : {$signed({reg370, reg373})}));
              reg379 <= (^wire363[(5'h10):(1'h0)]);
              reg380 <= (((^(wire334[(1'h0):(1'h0)] ?
                          $signed(reg382) : reg372[(4'h9):(4'h9)])) ?
                      wire363 : (+wire363)) ?
                  {$signed(wire363[(4'h9):(1'h1)])} : reg353[(1'h1):(1'h1)]);
              reg381 <= wire369;
              reg382 <= $unsigned($unsigned($signed((~$signed(wire366)))));
            end
          if ((+wire363))
            begin
              reg383 <= wire351;
              reg384 <= reg339[(4'he):(1'h1)];
            end
          else
            begin
              reg383 <= (+(&($signed(reg354) <= $unsigned((~^reg372)))));
              reg384 <= (^$signed((~(7'h40))));
              reg385 <= (($signed(((wire334 | reg370) ?
                  reg346 : {reg377})) <= $signed(reg360[(1'h1):(1'h1)])) <= reg339);
              reg386 <= {(((reg338[(5'h11):(5'h11)] ?
                          (reg347 <= reg347) : {wire334}) ?
                      $signed({reg370}) : $unsigned((+reg381))) < ((wire351[(5'h12):(2'h2)] <= $unsigned(reg370)) ?
                      $signed($signed(reg345)) : {wire364}))};
              reg387 <= $unsigned((wire333 ^~ (wire366[(2'h3):(1'h1)] ^ $signed(reg384[(2'h2):(1'h1)]))));
            end
          reg388 <= (-(((^$signed(reg362)) ?
              (reg360[(3'h7):(1'h1)] ?
                  (~|(8'hb5)) : $signed(reg344)) : reg360) ^ wire331[(4'h8):(2'h2)]));
        end
      else
        begin
          reg375 <= ((reg387[(2'h2):(1'h1)] ?
              reg345[(2'h3):(1'h0)] : (~$unsigned(reg343[(3'h7):(2'h2)]))) ^ reg372[(4'h8):(3'h6)]);
        end
      if (($signed(((|$signed(wire363)) | reg386)) ?
          $signed((+reg382[(3'h6):(3'h6)])) : reg355[(3'h4):(2'h3)]))
        begin
          reg389 <= wire367;
        end
      else
        begin
          if ((^~(7'h41)))
            begin
              reg389 <= (^~(^$unsigned(wire366[(2'h2):(1'h0)])));
              reg390 <= $signed($signed(reg389));
              reg391 <= (reg354 ?
                  $unsigned(($unsigned({reg385, (8'ha8)}) ?
                      ($signed((8'hb6)) ?
                          (^~(8'hbc)) : $unsigned(reg386)) : $unsigned($signed((8'hb2))))) : (!reg339));
              reg392 <= (8'had);
              reg393 <= {$unsigned($unsigned((~^$signed((8'h9d)))))};
            end
          else
            begin
              reg389 <= reg376;
              reg390 <= $unsigned(($unsigned(reg375[(4'hb):(1'h0)]) ?
                  reg373 : (wire332 ?
                      $unsigned(reg382[(1'h0):(1'h0)]) : (~|$signed(reg371)))));
              reg391 <= ($signed(wire369) ?
                  ($unsigned((reg362 != (!reg345))) ?
                      $signed(reg342[(4'he):(1'h1)]) : (((reg340 ?
                          reg355 : (8'hab)) << (reg392 * (8'hb5))) || (reg360[(2'h2):(1'h0)] >>> (wire334 ?
                          reg357 : reg376)))) : {reg379,
                      (reg350 || $unsigned($signed(reg341)))});
            end
        end
    end
  assign wire394 = reg389[(3'h6):(3'h5)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module304
#( parameter param326 = ({(((~(7'h44)) ? (~(8'had)) : ((7'h42) ? (7'h40) : (8'ha1))) == (|(^(8'ha0))))} ~^ (({{(8'hbd)}, ((8'hb0) ? (7'h42) : (7'h42))} ? {(&(8'hbc)), ((8'h9c) ? (8'ha8) : (8'hb9))} : ({(8'hb6)} & {(8'hbd), (8'haf)})) ? (~&(~&(8'ha2))) : ((&{(7'h41)}) != ((8'hbd) << (!(8'hb2))))))
, parameter param327 = (((~&(((8'hab) ? param326 : (8'ha1)) ^ (~param326))) && {((8'hbe) ? (param326 ? param326 : param326) : param326)}) == (^param326)) )
(y, clk, wire308, wire307, wire306, wire305);
  output wire [(32'hcc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire308;
  input wire [(4'h8):(1'h0)] wire307;
  input wire signed [(5'h15):(1'h0)] wire306;
  input wire [(2'h3):(1'h0)] wire305;
  wire signed [(4'hf):(1'h0)] wire325;
  reg signed [(3'h5):(1'h0)] reg324 = (1'h0);
  wire [(3'h5):(1'h0)] wire323;
  wire signed [(5'h10):(1'h0)] wire322;
  reg signed [(4'he):(1'h0)] reg321 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg320 = (1'h0);
  wire [(2'h2):(1'h0)] wire319;
  wire signed [(5'h15):(1'h0)] wire318;
  wire [(3'h5):(1'h0)] wire317;
  wire [(5'h12):(1'h0)] wire316;
  wire [(5'h14):(1'h0)] wire315;
  wire [(2'h3):(1'h0)] wire314;
  wire signed [(4'h9):(1'h0)] wire313;
  wire signed [(5'h15):(1'h0)] wire312;
  wire signed [(4'ha):(1'h0)] wire311;
  wire signed [(5'h12):(1'h0)] wire310;
  wire signed [(5'h12):(1'h0)] wire309;
  assign y = {wire325,
                 reg324,
                 wire323,
                 wire322,
                 reg321,
                 reg320,
                 wire319,
                 wire318,
                 wire317,
                 wire316,
                 wire315,
                 wire314,
                 wire313,
                 wire312,
                 wire311,
                 wire310,
                 wire309,
                 (1'h0)};
  assign wire309 = (wire308[(3'h6):(3'h5)] ?
                       {(&($signed(wire308) ? (&(7'h43)) : {wire306, wire306})),
                           (((wire307 && wire307) <= wire308[(2'h3):(1'h1)]) ?
                               wire306 : (wire306[(4'hf):(2'h3)] + (+wire306)))} : $unsigned((($unsigned((8'hb3)) - wire306[(2'h2):(2'h2)]) * wire307)));
  assign wire310 = (&{$unsigned(wire306[(3'h5):(2'h3)]),
                       (~(~$signed(wire308)))});
  assign wire311 = (8'h9c);
  assign wire312 = {(^(~^$unsigned($unsigned(wire310))))};
  assign wire313 = ((8'hae) | {(&wire312)});
  assign wire314 = (~$unsigned($unsigned(wire307[(3'h7):(3'h7)])));
  assign wire315 = (((~|wire314) ~^ ($unsigned(((8'had) ?
                           wire306 : wire307)) << wire307[(1'h0):(1'h0)])) ?
                       $unsigned(wire309[(5'h10):(4'hb)]) : wire306);
  assign wire316 = $unsigned((wire309[(1'h0):(1'h0)] ?
                       $signed((^~{(8'ha9)})) : ($signed({wire308}) ?
                           (~|{wire305}) : $signed((7'h41)))));
  assign wire317 = (&($unsigned(wire305) & (-(((8'hbf) ?
                       wire309 : wire305) << wire308))));
  assign wire318 = ($signed($unsigned(($signed(wire311) && $unsigned(wire312)))) ?
                       (wire311[(1'h0):(1'h0)] ?
                           {$unsigned($unsigned((8'hb7))),
                               wire309[(2'h2):(2'h2)]} : ($signed($signed(wire310)) ?
                               $signed((wire306 ?
                                   wire315 : wire315)) : ($signed(wire313) & (wire313 ?
                                   (8'h9d) : wire310)))) : $unsigned($unsigned($unsigned($signed(wire305)))));
  assign wire319 = (~^($unsigned(($signed(wire305) <= wire317)) > $unsigned(wire309[(4'hd):(4'hd)])));
  always
    @(posedge clk) begin
      reg320 <= wire311[(4'ha):(3'h4)];
      reg321 <= (((wire308 - (^(wire311 > wire314))) * $unsigned(wire317[(1'h0):(1'h0)])) > ($signed({wire308,
              wire318}) ?
          (((+wire307) & wire314[(2'h3):(2'h3)]) ?
              (wire317 < (^wire318)) : $signed((wire313 + wire310))) : ((8'haf) ?
              wire314 : ((wire317 ?
                  wire314 : wire308) && (wire308 >>> wire316)))));
    end
  assign wire322 = $unsigned(({wire307[(3'h4):(2'h3)], wire308} ?
                       reg320 : ((~&reg321) <<< (reg321 + {wire312,
                           wire312}))));
  assign wire323 = ($signed(wire305[(1'h1):(1'h1)]) ?
                       $signed((wire308[(1'h1):(1'h0)] == wire310)) : wire309[(4'hd):(2'h3)]);
  always
    @(posedge clk) begin
      reg324 <= wire318;
    end
  assign wire325 = $signed(wire309[(3'h5):(3'h4)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module555
#( parameter param1832 = ((((((8'hbf) >= (8'hbd)) ? ((8'haa) && (8'hbd)) : ((8'hba) ? (8'hb0) : (8'ha3))) ? (~(-(8'haf))) : (^~{(8'ha2), (8'hb8)})) ? {(((8'ha5) ? (8'hbc) : (8'h9f)) ? (8'hab) : ((7'h44) ? (8'ha5) : (8'hab))), (8'h9c)} : {{((8'hb8) <<< (8'hb8))}, ((~&(8'ha6)) ? (^(8'hb2)) : ((8'h9f) ? (7'h44) : (8'hba)))}) & {(((!(8'hbf)) ? (-(7'h44)) : {(8'hb8)}) ^~ ({(8'hb6)} ? {(8'hb3)} : (8'ha8)))})
, parameter param1833 = param1832 )
(y, clk, wire556, wire557, wire558, wire559, wire560);
  output wire [(32'h2f1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire556;
  input wire signed [(5'h12):(1'h0)] wire557;
  input wire [(5'h15):(1'h0)] wire558;
  input wire signed [(5'h15):(1'h0)] wire559;
  input wire [(5'h14):(1'h0)] wire560;
  wire [(4'h9):(1'h0)] wire1831;
  wire [(5'h13):(1'h0)] wire1830;
  wire [(3'h5):(1'h0)] wire1829;
  wire signed [(2'h2):(1'h0)] wire1828;
  wire signed [(4'h8):(1'h0)] wire1827;
  wire signed [(4'hf):(1'h0)] wire1826;
  wire [(5'h14):(1'h0)] wire1825;
  wire [(5'h10):(1'h0)] wire1824;
  wire [(4'h8):(1'h0)] wire1822;
  wire signed [(4'ha):(1'h0)] wire1821;
  wire signed [(4'ha):(1'h0)] wire1820;
  wire [(5'h12):(1'h0)] wire1818;
  wire [(5'h10):(1'h0)] wire561;
  wire signed [(5'h13):(1'h0)] wire903;
  wire [(4'h8):(1'h0)] wire905;
  reg [(4'ha):(1'h0)] reg906 = (1'h0);
  reg [(3'h6):(1'h0)] reg907 = (1'h0);
  reg [(4'hc):(1'h0)] reg908 = (1'h0);
  reg [(5'h14):(1'h0)] reg909 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg910 = (1'h0);
  reg [(4'ha):(1'h0)] reg911 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg912 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg913 = (1'h0);
  reg [(2'h3):(1'h0)] reg914 = (1'h0);
  reg [(5'h11):(1'h0)] reg915 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg916 = (1'h0);
  reg signed [(4'he):(1'h0)] reg917 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg918 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg919 = (1'h0);
  reg [(4'he):(1'h0)] reg920 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg921 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg922 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg923 = (1'h0);
  reg [(4'h9):(1'h0)] reg924 = (1'h0);
  reg [(4'hc):(1'h0)] reg925 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg926 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg927 = (1'h0);
  reg [(2'h2):(1'h0)] reg928 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg929 = (1'h0);
  reg [(3'h4):(1'h0)] reg930 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg931 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg932 = (1'h0);
  reg [(5'h11):(1'h0)] reg933 = (1'h0);
  reg [(4'hd):(1'h0)] reg934 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg935 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg936 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg937 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg938 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg939 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg940 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg941 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg942 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg943 = (1'h0);
  reg [(5'h15):(1'h0)] reg944 = (1'h0);
  reg [(4'h9):(1'h0)] reg945 = (1'h0);
  wire [(5'h11):(1'h0)] wire946;
  wire [(5'h11):(1'h0)] wire947;
  wire signed [(4'h9):(1'h0)] wire948;
  wire signed [(2'h3):(1'h0)] wire949;
  wire [(3'h6):(1'h0)] wire1004;
  wire [(2'h2):(1'h0)] wire1816;
  assign y = {wire1831,
                 wire1830,
                 wire1829,
                 wire1828,
                 wire1827,
                 wire1826,
                 wire1825,
                 wire1824,
                 wire1822,
                 wire1821,
                 wire1820,
                 wire1818,
                 wire561,
                 wire903,
                 wire905,
                 reg906,
                 reg907,
                 reg908,
                 reg909,
                 reg910,
                 reg911,
                 reg912,
                 reg913,
                 reg914,
                 reg915,
                 reg916,
                 reg917,
                 reg918,
                 reg919,
                 reg920,
                 reg921,
                 reg922,
                 reg923,
                 reg924,
                 reg925,
                 reg926,
                 reg927,
                 reg928,
                 reg929,
                 reg930,
                 reg931,
                 reg932,
                 reg933,
                 reg934,
                 reg935,
                 reg936,
                 reg937,
                 reg938,
                 reg939,
                 reg940,
                 reg941,
                 reg942,
                 reg943,
                 reg944,
                 reg945,
                 wire946,
                 wire947,
                 wire948,
                 wire949,
                 wire1004,
                 wire1816,
                 (1'h0)};
  assign wire561 = wire558[(4'hc):(4'ha)];
  module562 modinst904 (.clk(clk), .wire565(wire558), .wire566(wire557), .wire564(wire560), .wire563(wire559), .y(wire903));
  assign wire905 = ((($unsigned((8'haf)) > wire558) + wire557[(4'hd):(3'h4)]) ?
                       ((((8'ha9) ?
                           wire556[(4'hd):(4'h8)] : $signed(wire558)) != $signed({(8'ha7),
                           wire556})) * $signed(wire558)) : $signed(((^$unsigned(wire556)) + wire557)));
  always
    @(posedge clk) begin
      if ((wire905[(3'h6):(2'h3)] > $unsigned(wire561[(2'h3):(2'h2)])))
        begin
          reg906 <= (~^(&wire558));
        end
      else
        begin
          reg906 <= wire560;
          if (wire905)
            begin
              reg907 <= wire905[(3'h6):(2'h2)];
              reg908 <= wire558;
              reg909 <= $signed((!(reg906[(3'h7):(3'h4)] ?
                  $unsigned((~|wire559)) : wire560[(3'h7):(2'h3)])));
              reg910 <= ($unsigned((($signed((8'ha6)) ~^ wire556) + $unsigned((~(8'hb0))))) ?
                  wire558 : reg909);
            end
          else
            begin
              reg907 <= {$signed($signed((8'ha8)))};
              reg908 <= (8'hb7);
              reg909 <= (wire903 * {($unsigned(wire561[(2'h3):(1'h1)]) || {$signed((8'hbd)),
                      $signed(wire559)})});
            end
          reg911 <= (wire557 ?
              $signed(wire559) : ((($unsigned(reg906) ?
                  (reg908 ?
                      (8'ha0) : wire556) : reg910) > $signed({wire558})) ~^ (($signed(wire560) ?
                  {reg907, reg910} : ((8'hbf) ?
                      wire559 : wire903)) | {$unsigned(wire557),
                  $unsigned(wire561)})));
          reg912 <= ($signed(({(reg908 ? reg907 : (8'ha5)),
                  $signed(reg911)} <<< reg909[(4'hc):(1'h1)])) ?
              (+reg906) : wire558);
          if (reg908)
            begin
              reg913 <= $unsigned(wire557);
              reg914 <= $signed(((reg909[(5'h11):(5'h11)] < wire559[(5'h10):(5'h10)]) - ({(reg911 ?
                      wire560 : reg908)} * $signed((~&reg911)))));
              reg915 <= reg913;
            end
          else
            begin
              reg913 <= $unsigned((($signed(wire558[(5'h10):(1'h1)]) ~^ reg912[(2'h3):(2'h3)]) ?
                  $signed(($unsigned(reg913) >>> $unsigned(wire558))) : ($signed($unsigned(wire558)) != (((8'hab) >= wire556) <= $signed(wire556)))));
            end
        end
      if ($unsigned((|reg907[(2'h2):(1'h0)])))
        begin
          reg916 <= reg911[(3'h4):(1'h0)];
          reg917 <= (wire905 ?
              (^~$unsigned(reg907)) : $unsigned($signed($unsigned(reg913))));
          reg918 <= wire559[(4'h9):(4'h8)];
        end
      else
        begin
          reg916 <= {((reg916[(4'hf):(3'h4)] ?
                  reg911 : $signed((reg915 ? wire558 : reg911))) || {reg913})};
          if (((!$signed(reg917[(3'h4):(1'h0)])) ?
              reg916 : {({reg916} >= {{reg914}})}))
            begin
              reg917 <= {({wire557,
                          ((reg913 | reg918) ?
                              $unsigned(wire561) : $signed(reg908))} ?
                      (reg913 ?
                          (!((8'ha4) ?
                              (8'ha0) : wire556)) : (8'hb4)) : {($signed(reg918) ?
                              (|reg915) : (-wire561)),
                          $unsigned($signed(reg914))})};
              reg918 <= reg918;
              reg919 <= $unsigned((($unsigned((^wire561)) ?
                      $unsigned({(8'hab),
                          reg917}) : $signed(((8'hbd) > reg918))) ?
                  wire559 : (($signed((8'hba)) ?
                          $unsigned(reg911) : (wire903 ? reg907 : reg915)) ?
                      (~^(+reg912)) : $signed($signed(reg914)))));
              reg920 <= (wire557 ?
                  (reg910 ?
                      $unsigned(($signed(reg914) < $unsigned(reg917))) : ((~^(&(7'h40))) ?
                          (8'hbd) : wire905)) : $unsigned((((reg912 || reg919) == $signed(wire557)) ?
                      ((reg915 >>> reg909) ?
                          reg908 : (wire903 ^~ reg917)) : {$signed(reg916)})));
            end
          else
            begin
              reg917 <= ((&(((reg917 ?
                      reg917 : wire903) ~^ ((8'ha5) >> reg912)) ^ $signed(reg908))) ?
                  (wire559 ~^ $unsigned((~^(reg908 >>> reg913)))) : reg916);
              reg918 <= $signed(reg914);
              reg919 <= (^(^~(reg913[(3'h7):(3'h5)] << {$signed(reg910)})));
              reg920 <= $unsigned($unsigned($unsigned(wire558[(4'hc):(1'h0)])));
            end
          if ($signed((~($signed($signed(reg917)) && $unsigned(wire556)))))
            begin
              reg921 <= $unsigned(($unsigned($signed($signed(reg910))) >> (reg913 >>> (~&(wire561 || reg907)))));
              reg922 <= {(~(-reg910[(2'h3):(2'h2)])),
                  (^$unsigned(reg907[(3'h5):(3'h4)]))};
              reg923 <= wire557[(5'h11):(4'hf)];
            end
          else
            begin
              reg921 <= reg912;
              reg922 <= wire903[(1'h0):(1'h0)];
              reg923 <= reg908[(4'hc):(3'h4)];
              reg924 <= reg910;
            end
          reg925 <= {(($signed(reg912) < (reg912[(4'hd):(4'h8)] ?
                  (reg924 ?
                      wire557 : (7'h40)) : (~^reg916))) || reg915[(1'h1):(1'h1)]),
              $unsigned((&$unsigned(((8'ha9) ? reg920 : reg917))))};
        end
      if ((8'hac))
        begin
          reg926 <= $signed((&reg912[(1'h1):(1'h1)]));
        end
      else
        begin
          reg926 <= (reg912[(3'h6):(2'h3)] >= $unsigned(reg923[(2'h2):(1'h0)]));
          reg927 <= reg921[(4'he):(1'h0)];
          reg928 <= ($unsigned((reg927[(1'h0):(1'h0)] ?
              (&(&wire560)) : wire903[(4'ha):(1'h0)])) << {(~&reg906)});
        end
      reg929 <= $unsigned($unsigned({reg925[(4'hc):(4'hb)]}));
    end
  always
    @(posedge clk) begin
      reg930 <= {{{reg906, $signed((&wire561))}},
          $signed((+((+(8'ha5)) ? $signed(wire559) : reg911)))};
      if (($signed(((~^(reg907 ?
              reg926 : reg923)) && $unsigned($signed(wire561)))) ?
          reg921[(3'h6):(1'h0)] : (^reg925)))
        begin
          reg931 <= $unsigned((reg930 ?
              $signed((~^(wire559 == reg913))) : {reg927[(1'h0):(1'h0)]}));
          if (wire558[(3'h7):(3'h4)])
            begin
              reg932 <= $signed((8'haa));
            end
          else
            begin
              reg932 <= reg908;
              reg933 <= reg920;
              reg934 <= ($unsigned(reg921[(4'h9):(1'h1)]) ?
                  reg910 : (^~reg914[(1'h1):(1'h1)]));
              reg935 <= (7'h44);
              reg936 <= $signed($signed((reg926 != (~|{wire903}))));
            end
          reg937 <= (~^reg906);
          if ($unsigned($signed((+$unsigned((reg909 ? reg922 : reg928))))))
            begin
              reg938 <= $signed($unsigned(reg908[(4'h9):(1'h1)]));
            end
          else
            begin
              reg938 <= {(reg915 ?
                      $signed($signed($unsigned(wire905))) : wire557),
                  $unsigned(reg917[(1'h0):(1'h0)])};
            end
          if ($unsigned((8'ha3)))
            begin
              reg939 <= ((((&(~reg906)) | (!$signed(reg931))) | ((+$signed((8'ha1))) ~^ reg930[(2'h3):(2'h3)])) <= ({{reg926[(3'h4):(1'h1)]},
                      $unsigned($signed(reg913))} ?
                  reg926 : reg924[(4'h9):(1'h0)]));
              reg940 <= ($signed((~((~(8'hb2)) << $signed(reg926)))) * wire905[(1'h1):(1'h0)]);
            end
          else
            begin
              reg939 <= reg913;
              reg940 <= $unsigned(((reg925[(3'h5):(1'h0)] ?
                  $signed($unsigned(wire557)) : reg924) ^~ (!(|$signed(reg911)))));
              reg941 <= (^{$signed({(reg927 & reg911)})});
              reg942 <= {$signed((|{$unsigned((8'hb3)), (reg917 >= (8'ha8))}))};
            end
        end
      else
        begin
          reg931 <= $unsigned($signed(reg911));
          reg932 <= (!$unsigned((!((reg930 ? wire559 : reg914) ?
              $unsigned(reg907) : (wire557 ? reg927 : reg919)))));
          reg933 <= (!$signed($unsigned((~reg925[(4'h8):(1'h0)]))));
          reg934 <= reg906[(3'h4):(2'h3)];
          if ($unsigned(reg928))
            begin
              reg935 <= $unsigned($signed($unsigned($signed(reg910[(4'he):(1'h1)]))));
              reg936 <= (wire560 ^ (reg930 ?
                  reg910[(4'ha):(1'h1)] : (($signed(wire557) ?
                      (7'h44) : reg906) >> wire557[(4'h9):(2'h2)])));
            end
          else
            begin
              reg935 <= $unsigned((~(~|{{reg915}})));
              reg936 <= $signed({$unsigned($signed(reg914)), reg933});
              reg937 <= $unsigned(((reg941[(4'h9):(3'h7)] ?
                  reg927[(4'h8):(3'h7)] : $unsigned(reg925)) >>> {{((8'haa) <= reg913),
                      $unsigned(reg920)},
                  $signed({reg933})}));
              reg938 <= $unsigned((!reg940));
            end
        end
      reg943 <= $signed($signed(reg932[(4'hd):(2'h3)]));
      reg944 <= $unsigned(reg923[(1'h1):(1'h1)]);
      reg945 <= reg930;
    end
  assign wire946 = (^$signed($signed(reg906[(2'h2):(1'h1)])));
  assign wire947 = reg917[(3'h7):(2'h2)];
  assign wire948 = $signed(((+(reg933 || {reg911,
                       (8'ha5)})) == $unsigned($signed({reg908}))));
  assign wire949 = (reg907[(2'h2):(1'h1)] || reg913);
  module950 modinst1005 (.wire951(reg938), .wire954(reg919), .wire952(reg915), .y(wire1004), .clk(clk), .wire953(reg922));
  module1006 modinst1817 (.clk(clk), .wire1011(reg933), .y(wire1816), .wire1010(reg944), .wire1008(reg917), .wire1007(wire905), .wire1009(reg929));
  module675 modinst1819 (.wire679(reg938), .wire677(reg945), .clk(clk), .wire678(wire903), .wire676(reg915), .y(wire1818));
  assign wire1820 = (($unsigned((8'ha7)) ?
                            (reg921 & $unsigned($signed(reg928))) : $signed(((~^(8'hac)) && reg916[(3'h6):(1'h0)]))) ?
                        reg912 : $signed((((wire903 > wire561) ?
                            reg907 : {wire560}) < reg925)));
  assign wire1821 = reg934[(1'h1):(1'h0)];
  module675 modinst1823 (.wire679(wire561), .wire678(reg916), .wire676(reg938), .clk(clk), .wire677(wire948), .y(wire1822));
  assign wire1824 = (~&(($unsigned((reg932 ? reg926 : reg915)) ?
                        {wire1004} : ($unsigned(reg938) <= (reg937 ?
                            reg915 : reg911))) == (((reg923 ?
                            reg907 : wire949) ?
                        reg908[(1'h1):(1'h0)] : (~^wire946)) + wire948[(3'h4):(3'h4)])));
  assign wire1825 = (-$unsigned(reg912));
  assign wire1826 = (+((|(~(~^reg938))) == reg937[(4'h9):(4'h8)]));
  assign wire1827 = reg931[(1'h0):(1'h0)];
  assign wire1828 = {$unsigned(reg941[(5'h11):(3'h5)])};
  assign wire1829 = $unsigned(((8'hb9) ^ $signed(((reg929 ? wire947 : reg919) ?
                        $signed(wire1818) : (wire1825 > reg918)))));
  assign wire1830 = wire561[(4'hc):(1'h1)];
  assign wire1831 = wire1824[(4'he):(4'h9)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1006
#( parameter param1815 = ((^~{((^(8'hac)) ^~ ((8'hb2) <<< (8'hb3))), ((!(7'h44)) ? (8'hbd) : (^(8'hbd)))}) ? ((((^~(8'hb8)) ? (-(8'hb6)) : ((8'ha2) <<< (8'ha5))) ? {((8'haa) ? (8'had) : (8'ha2)), {(8'hb4)}} : (8'h9e)) ? ((~|((8'hbf) ? (8'hbc) : (8'hb6))) == (((7'h43) ? (8'hb6) : (8'hb6)) ? ((8'hbd) ? (8'ha2) : (8'hbb)) : ((8'hb4) ^ (8'hab)))) : (+(~^(~|(8'ha3))))) : (~&{({(8'ha1)} ? (~&(8'ha7)) : ((7'h44) >> (8'hba))), (^((8'hbc) ? (8'hae) : (7'h40)))})) )
(y, clk, wire1011, wire1010, wire1009, wire1008, wire1007);
  output wire [(32'h1d8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire1011;
  input wire [(5'h14):(1'h0)] wire1010;
  input wire [(5'h14):(1'h0)] wire1009;
  input wire [(4'he):(1'h0)] wire1008;
  input wire [(2'h3):(1'h0)] wire1007;
  wire [(4'ha):(1'h0)] wire1309;
  wire [(5'h10):(1'h0)] wire1155;
  wire signed [(4'ha):(1'h0)] wire1153;
  wire signed [(4'he):(1'h0)] wire1139;
  wire [(5'h15):(1'h0)] wire1138;
  wire [(5'h13):(1'h0)] wire1136;
  wire [(5'h13):(1'h0)] wire1067;
  wire [(5'h14):(1'h0)] wire1066;
  wire signed [(5'h13):(1'h0)] wire1064;
  wire [(5'h12):(1'h0)] wire1012;
  wire [(5'h13):(1'h0)] wire1311;
  wire signed [(4'hd):(1'h0)] wire1312;
  reg [(4'hf):(1'h0)] reg1313 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1314 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1315 = (1'h0);
  reg [(5'h13):(1'h0)] reg1316 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1317 = (1'h0);
  reg [(2'h3):(1'h0)] reg1318 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1319 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1320 = (1'h0);
  reg [(2'h3):(1'h0)] reg1321 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1322 = (1'h0);
  reg [(5'h14):(1'h0)] reg1323 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1324 = (1'h0);
  reg [(5'h12):(1'h0)] reg1325 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1326 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire1696;
  wire [(5'h13):(1'h0)] wire1713;
  wire signed [(4'hb):(1'h0)] wire1715;
  wire signed [(4'hf):(1'h0)] wire1716;
  wire [(3'h6):(1'h0)] wire1717;
  wire signed [(4'h9):(1'h0)] wire1718;
  wire signed [(4'h9):(1'h0)] wire1719;
  wire [(5'h12):(1'h0)] wire1813;
  assign y = {wire1309,
                 wire1155,
                 wire1153,
                 wire1139,
                 wire1138,
                 wire1136,
                 wire1067,
                 wire1066,
                 wire1064,
                 wire1012,
                 wire1311,
                 wire1312,
                 reg1313,
                 reg1314,
                 reg1315,
                 reg1316,
                 reg1317,
                 reg1318,
                 reg1319,
                 reg1320,
                 reg1321,
                 reg1322,
                 reg1323,
                 reg1324,
                 reg1325,
                 reg1326,
                 wire1696,
                 wire1713,
                 wire1715,
                 wire1716,
                 wire1717,
                 wire1718,
                 wire1719,
                 wire1813,
                 (1'h0)};
  assign wire1012 = (!wire1011[(3'h4):(3'h4)]);
  module1013 modinst1065 (wire1064, clk, wire1010, wire1008, wire1012, wire1011);
  assign wire1066 = {$signed(wire1007[(1'h1):(1'h1)]),
                        {$unsigned(((wire1010 ? wire1012 : wire1011) ?
                                wire1008 : $unsigned(wire1012)))}};
  assign wire1067 = wire1012[(5'h10):(4'ha)];
  module1068 modinst1137 (.wire1069(wire1007), .wire1072(wire1010), .clk(clk), .wire1071(wire1066), .y(wire1136), .wire1070(wire1067));
  assign wire1138 = {wire1067[(4'hf):(3'h5)], (8'ha0)};
  assign wire1139 = ($unsigned((~&(8'hbf))) + wire1067);
  module1140 modinst1154 (wire1153, clk, wire1008, wire1012, wire1011, wire1138);
  assign wire1155 = ((+($signed($signed(wire1138)) ?
                        {(wire1007 ? wire1008 : wire1066),
                            wire1010} : wire1009)) << $unsigned((&wire1067[(4'h8):(4'h8)])));
  module1156 modinst1310 (.y(wire1309), .wire1157(wire1010), .clk(clk), .wire1160(wire1008), .wire1159(wire1136), .wire1161(wire1012), .wire1158(wire1153));
  assign wire1311 = (+$unsigned({wire1155}));
  assign wire1312 = ($signed(wire1007[(2'h3):(2'h2)]) & ((($unsigned(wire1064) ?
                            $unsigned(wire1309) : $signed((8'ha5))) ?
                        $unsigned($signed(wire1067)) : $signed({wire1067,
                            wire1008})) * ($unsigned($unsigned(wire1153)) <<< (((7'h43) ?
                        wire1153 : (8'ha3)) >= $unsigned(wire1155)))));
  always
    @(posedge clk) begin
      reg1313 <= wire1311[(4'ha):(4'h9)];
      reg1314 <= ({{$unsigned(wire1007),
              (8'ha0)}} < (wire1155 && (({wire1012} ~^ {wire1010}) ?
          $unsigned($unsigned(wire1008)) : ((wire1138 ?
              (8'hac) : (8'hb6)) << (~&wire1007)))));
      if ($signed((({(wire1064 && wire1011), (|wire1309)} ?
          $signed($unsigned(wire1067)) : (wire1153 > ((8'hb2) ?
              wire1064 : reg1313))) ^ {$unsigned($signed(wire1064)),
          wire1155[(1'h1):(1'h1)]})))
        begin
          reg1315 <= {(8'ha9)};
          if (wire1011)
            begin
              reg1316 <= (({$signed((8'hba)),
                      $unsigned({(8'hb9), wire1312})} + wire1010) ?
                  $unsigned(($unsigned(((8'haa) - wire1012)) == ((~&wire1010) ~^ (reg1313 | wire1153)))) : $unsigned((+((wire1011 >= wire1012) ?
                      wire1311[(3'h4):(2'h2)] : (wire1312 ?
                          wire1312 : wire1312)))));
              reg1317 <= $signed(wire1007[(1'h0):(1'h0)]);
            end
          else
            begin
              reg1316 <= (|reg1315);
              reg1317 <= reg1315[(2'h3):(2'h3)];
              reg1318 <= (~|$signed(($unsigned((wire1153 < (8'ha4))) ?
                  $signed((8'hba)) : $signed($signed(wire1312)))));
              reg1319 <= wire1155;
            end
          reg1320 <= ($unsigned(wire1008) ?
              (^(wire1009 < ((wire1067 ^ (8'had)) ?
                  (wire1155 ?
                      reg1315 : reg1314) : (wire1136 - (8'hb3))))) : ((reg1319 | (wire1138[(4'hf):(2'h2)] - reg1316[(3'h5):(2'h3)])) > wire1009));
          if ((wire1139[(3'h5):(3'h4)] & ((8'hbd) && ($unsigned({wire1136}) ?
              (|(wire1312 & reg1320)) : ((reg1316 ^ wire1138) != $signed(wire1064))))))
            begin
              reg1321 <= $unsigned({{(~(!(7'h44))),
                      {((8'hb5) ? reg1319 : (8'ha6)), (+wire1009)}},
                  (wire1312[(2'h2):(1'h1)] >> reg1318[(2'h3):(2'h2)])});
              reg1322 <= {($signed((!(~^wire1007))) ?
                      ($unsigned((~&wire1139)) ?
                          $signed({wire1139}) : (^~wire1309[(1'h1):(1'h1)])) : wire1155)};
              reg1323 <= $signed(reg1322[(1'h1):(1'h1)]);
              reg1324 <= $unsigned($unsigned(($signed((reg1323 ?
                  reg1323 : wire1011)) != wire1136)));
            end
          else
            begin
              reg1321 <= reg1318;
              reg1322 <= $unsigned($signed((~reg1324[(1'h1):(1'h0)])));
              reg1323 <= (wire1009[(3'h5):(1'h0)] >>> reg1317);
              reg1324 <= (wire1066 * {(!$unsigned(wire1007)),
                  reg1318[(1'h0):(1'h0)]});
            end
          if ($signed($unsigned(reg1320[(1'h1):(1'h1)])))
            begin
              reg1325 <= ($signed(({{reg1320, reg1320}} ?
                      wire1139[(3'h5):(1'h1)] : reg1323)) ?
                  ((((-reg1318) ?
                              $signed(reg1318) : ((8'hbf) ?
                                  wire1067 : (8'haf))) ?
                          wire1139 : (reg1323 & wire1311[(4'he):(3'h4)])) ?
                      $unsigned(reg1323) : wire1009[(3'h6):(3'h4)]) : ((reg1315 >>> $unsigned(wire1009[(3'h6):(2'h3)])) + reg1322[(2'h3):(2'h2)]));
              reg1326 <= $signed($signed(reg1316));
            end
          else
            begin
              reg1325 <= ((($signed($unsigned(wire1007)) != wire1312) | $signed((~&reg1320))) <<< reg1326[(4'h8):(3'h6)]);
              reg1326 <= (+(7'h43));
            end
        end
      else
        begin
          reg1315 <= $unsigned($signed((~^$unsigned((reg1326 | wire1009)))));
          reg1316 <= {wire1008};
          if ($unsigned(reg1313[(3'h4):(1'h0)]))
            begin
              reg1317 <= (+wire1311[(4'hc):(4'hc)]);
              reg1318 <= (8'ha2);
            end
          else
            begin
              reg1317 <= (wire1009 ?
                  $signed($signed(reg1320)) : ($signed({(~^wire1008),
                      wire1064}) | wire1153[(2'h3):(2'h2)]));
              reg1318 <= wire1067[(1'h1):(1'h0)];
              reg1319 <= reg1319[(1'h0):(1'h0)];
            end
        end
    end
  module1327 modinst1697 (.wire1331(wire1155), .wire1328(wire1009), .clk(clk), .wire1330(reg1322), .wire1329(wire1011), .y(wire1696));
  module1698 modinst1714 (.wire1701(wire1155), .clk(clk), .wire1700(wire1312), .wire1702(wire1064), .y(wire1713), .wire1699(reg1326));
  assign wire1715 = $unsigned((^~{$unsigned((reg1319 & wire1067))}));
  assign wire1716 = $unsigned(((&wire1153[(3'h5):(1'h0)]) > wire1309));
  assign wire1717 = (~&$unsigned({wire1713[(2'h2):(1'h1)]}));
  assign wire1718 = reg1322[(4'h8):(1'h1)];
  assign wire1719 = wire1153[(3'h4):(2'h2)];
  module1720 modinst1814 (.clk(clk), .y(wire1813), .wire1722(wire1713), .wire1723(reg1316), .wire1721(wire1138), .wire1724(reg1323), .wire1725(reg1314));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module950
#( parameter param1002 = ((({((8'h9d) ? (8'hb9) : (8'hbb)), (|(8'ha1))} >> ((~&(8'ha5)) ? {(8'hae)} : ((8'hb3) < (8'hbc)))) ? (~^{{(8'hb0)}}) : (({(8'hbb), (8'ha9)} ? (+(7'h42)) : ((8'ha5) <<< (8'hac))) ? ((-(8'hb7)) + (~(8'hbe))) : ((~^(8'ha7)) ? {(8'hb3)} : ((8'h9c) ? (8'hab) : (7'h43))))) || ((^~(((8'ha7) >= (8'hb4)) | ((8'hac) || (7'h44)))) != (8'ha5)))
, parameter param1003 = (~&(~|(^~((param1002 <= param1002) ? (param1002 ? param1002 : param1002) : (!param1002))))) )
(y, clk, wire954, wire953, wire952, wire951);
  output wire [(32'h24f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire954;
  input wire [(5'h10):(1'h0)] wire953;
  input wire [(3'h4):(1'h0)] wire952;
  input wire signed [(5'h10):(1'h0)] wire951;
  wire [(5'h12):(1'h0)] wire1001;
  wire [(5'h11):(1'h0)] wire1000;
  wire [(4'he):(1'h0)] wire999;
  wire signed [(3'h6):(1'h0)] wire998;
  reg signed [(4'h8):(1'h0)] reg997 = (1'h0);
  reg [(5'h11):(1'h0)] reg996 = (1'h0);
  wire [(4'h9):(1'h0)] wire995;
  wire [(5'h13):(1'h0)] wire994;
  wire [(4'h9):(1'h0)] wire993;
  wire [(3'h5):(1'h0)] wire992;
  reg [(5'h13):(1'h0)] reg991 = (1'h0);
  reg [(4'hc):(1'h0)] reg990 = (1'h0);
  reg [(4'hb):(1'h0)] reg989 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg988 = (1'h0);
  reg [(4'hf):(1'h0)] reg987 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg986 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg985 = (1'h0);
  reg [(5'h14):(1'h0)] reg984 = (1'h0);
  reg [(3'h6):(1'h0)] reg983 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg982 = (1'h0);
  reg [(5'h12):(1'h0)] reg981 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg980 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg979 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg978 = (1'h0);
  reg [(3'h5):(1'h0)] reg977 = (1'h0);
  reg signed [(4'he):(1'h0)] reg976 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg975 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire974;
  wire signed [(3'h7):(1'h0)] wire973;
  wire signed [(3'h5):(1'h0)] wire972;
  reg [(5'h11):(1'h0)] reg971 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg970 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg969 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg968 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg967 = (1'h0);
  reg [(5'h12):(1'h0)] reg966 = (1'h0);
  reg [(4'ha):(1'h0)] reg965 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg964 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg963 = (1'h0);
  reg [(3'h6):(1'h0)] reg962 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg961 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire960;
  wire [(5'h14):(1'h0)] wire959;
  wire [(4'he):(1'h0)] wire958;
  wire [(4'h8):(1'h0)] wire957;
  wire signed [(4'h8):(1'h0)] wire956;
  wire [(4'he):(1'h0)] wire955;
  assign y = {wire1001,
                 wire1000,
                 wire999,
                 wire998,
                 reg997,
                 reg996,
                 wire995,
                 wire994,
                 wire993,
                 wire992,
                 reg991,
                 reg990,
                 reg989,
                 reg988,
                 reg987,
                 reg986,
                 reg985,
                 reg984,
                 reg983,
                 reg982,
                 reg981,
                 reg980,
                 reg979,
                 reg978,
                 reg977,
                 reg976,
                 reg975,
                 wire974,
                 wire973,
                 wire972,
                 reg971,
                 reg970,
                 reg969,
                 reg968,
                 reg967,
                 reg966,
                 reg965,
                 reg964,
                 reg963,
                 reg962,
                 reg961,
                 wire960,
                 wire959,
                 wire958,
                 wire957,
                 wire956,
                 wire955,
                 (1'h0)};
  assign wire955 = wire951[(3'h4):(2'h3)];
  assign wire956 = $signed(wire954);
  assign wire957 = wire951[(2'h2):(2'h2)];
  assign wire958 = (&wire956[(2'h3):(2'h3)]);
  assign wire959 = ($signed($unsigned(wire954[(3'h5):(3'h4)])) ?
                       wire952[(2'h3):(1'h0)] : ((8'ha9) != (!(wire951 ?
                           (wire958 ?
                               wire952 : wire955) : $unsigned(wire957)))));
  assign wire960 = wire958[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      if ((8'hae))
        begin
          reg961 <= ((wire956[(3'h6):(3'h5)] ^~ (~^{{wire957}, wire956})) ?
              ({($signed(wire957) >>> (~^wire952))} && (((^~wire956) ?
                  wire954 : wire953[(3'h5):(2'h2)]) << ($signed(wire951) > (+wire953)))) : ((((!(8'hbe)) ?
                      (wire959 ? wire951 : wire959) : wire957) ?
                  $signed($unsigned(wire951)) : ($unsigned(wire951) ?
                      (8'haf) : (+wire953))) + wire958));
          if ((&wire955))
            begin
              reg962 <= $signed((($signed((|wire956)) ?
                      (+wire952) : $signed((~wire959))) ?
                  ((wire953 ?
                      (wire951 != wire957) : (+(8'haa))) >= wire954[(2'h3):(1'h0)]) : $signed((~|((8'hab) ?
                      (8'hb2) : wire953)))));
              reg963 <= ((wire957 > (~&(wire956 ^~ $signed(wire951)))) < wire952[(3'h4):(1'h1)]);
              reg964 <= wire954;
              reg965 <= (wire953 ?
                  ($unsigned((wire953[(1'h1):(1'h1)] ?
                          $unsigned(wire955) : reg962)) ?
                      $unsigned(((|reg963) ?
                          reg962 : $signed((8'had)))) : reg962) : $signed($unsigned(((wire954 ?
                      wire954 : wire958) << (wire953 ~^ reg961)))));
            end
          else
            begin
              reg962 <= $unsigned((wire954[(4'h8):(2'h2)] | (&wire955[(4'ha):(3'h4)])));
            end
        end
      else
        begin
          reg961 <= wire956;
        end
      reg966 <= ((8'ha8) ?
          ($signed(($signed(reg964) ? wire958 : (wire952 ^ reg964))) ?
              (wire951 < $unsigned((wire957 >= wire954))) : wire960) : reg961);
      if ((|(wire953[(3'h4):(1'h0)] + ((^$signed((8'ha6))) ?
          (reg962[(3'h4):(2'h2)] >= (wire956 ?
              (8'ha4) : wire955)) : $signed(((7'h44) == wire955))))))
        begin
          reg967 <= ({{(|{wire952, wire956}), (+wire957[(3'h7):(3'h6)])},
                  (7'h40)} ?
              $unsigned({(~$signed(wire957))}) : (!(($unsigned(reg964) < $unsigned(reg964)) ?
                  $signed((~^wire954)) : {$unsigned((7'h44))})));
          if ($signed(((&(-$signed(wire953))) ?
              (($unsigned(wire959) ^~ $unsigned(reg961)) | $unsigned(((8'hb9) ^ wire951))) : wire960)))
            begin
              reg968 <= $unsigned(reg966);
              reg969 <= $unsigned(((~|reg962) >> {$unsigned((wire951 << reg965))}));
            end
          else
            begin
              reg968 <= reg964[(2'h3):(1'h0)];
              reg969 <= $unsigned($signed($unsigned($signed($signed(wire953)))));
              reg970 <= (($unsigned(((~^reg964) ? {(8'h9c)} : (~&wire956))) ?
                      (wire958[(4'hc):(4'ha)] ?
                          ($unsigned(wire953) >= (reg969 * reg969)) : (+(wire953 ?
                              (8'hbf) : wire960))) : (~($signed(wire952) > $signed(wire957)))) ?
                  ({$unsigned({wire955})} > $signed(((^(8'hba)) ^ wire953[(4'hb):(4'h8)]))) : {wire952});
              reg971 <= ((+((reg961[(4'h8):(2'h3)] + $unsigned(reg967)) ?
                  wire959[(4'hc):(4'hc)] : wire952[(1'h0):(1'h0)])) >= (~reg967));
            end
        end
      else
        begin
          reg967 <= $unsigned($unsigned($signed(wire955)));
          reg968 <= reg965;
          if (wire959)
            begin
              reg969 <= (8'ha1);
              reg970 <= reg963;
              reg971 <= $signed($unsigned(((reg968 ?
                      (&wire954) : (wire953 ? wire952 : wire959)) ?
                  reg971[(4'hb):(1'h1)] : (wire959 != wire955[(3'h5):(3'h5)]))));
            end
          else
            begin
              reg969 <= $unsigned({(~&reg970),
                  $signed($signed($signed((8'ha9))))});
            end
        end
    end
  assign wire972 = {(8'ha9), (~^reg961[(5'h10):(4'hb)])};
  assign wire973 = (!$unsigned($signed($signed(wire959))));
  assign wire974 = ((($signed($unsigned(reg965)) ?
                       (^~wire951) : (wire958 == $signed(wire954))) * $signed((&$signed(reg971)))) < (8'hb4));
  always
    @(posedge clk) begin
      if ({$unsigned(((wire974[(3'h6):(3'h4)] ?
              wire959[(4'h9):(2'h3)] : $signed(reg961)) + ((reg961 ?
              wire956 : reg969) >>> ((8'hb8) ? wire959 : reg971)))),
          (-$unsigned(($unsigned(wire956) ?
              wire954[(4'h9):(3'h7)] : {reg965})))})
        begin
          reg975 <= reg971[(2'h3):(2'h3)];
          reg976 <= {reg964};
        end
      else
        begin
          reg975 <= (wire955 ^ (($signed((+reg971)) ?
                  reg975 : reg965[(2'h2):(1'h0)]) ?
              wire956 : $unsigned(({wire957} ?
                  $unsigned(wire954) : (-wire957)))));
          reg976 <= (reg975[(3'h5):(2'h2)] ?
              $signed(({(reg963 ?
                      reg962 : wire953)} <<< (8'haa))) : (^{$unsigned((wire955 ?
                      reg971 : reg971)),
                  reg975}));
          reg977 <= reg962;
          reg978 <= (((-(+(~|reg970))) > {((wire955 << reg968) | $unsigned((8'hae)))}) ?
              ((~|$signed(reg963)) != $signed((8'h9e))) : $signed({reg971[(5'h10):(4'hb)],
                  (8'hba)}));
        end
      reg979 <= $signed(wire974[(4'h9):(1'h1)]);
      reg980 <= reg961;
      reg981 <= (($signed({wire956[(3'h4):(2'h2)],
          $unsigned(wire956)}) & (reg968[(3'h7):(2'h3)] ?
          ({wire956, wire952} ?
              $signed(wire959) : $signed((7'h44))) : (8'hb3))) ^ reg966[(4'hb):(2'h3)]);
      if ($unsigned((((^~reg970) ?
              ($signed(reg967) ?
                  (^~reg965) : wire974) : wire960[(4'he):(4'he)]) ?
          (&$signed((~|reg981))) : $signed($signed((reg980 ?
              wire957 : wire957))))))
        begin
          if ($signed(reg965[(3'h5):(2'h3)]))
            begin
              reg982 <= (8'ha5);
              reg983 <= $unsigned($unsigned(reg963[(2'h2):(2'h2)]));
            end
          else
            begin
              reg982 <= wire973[(2'h3):(1'h0)];
              reg983 <= reg967;
              reg984 <= reg979;
              reg985 <= reg981[(4'hb):(4'h8)];
            end
          reg986 <= (((({reg961} << reg976) ?
                      reg975[(4'h9):(3'h7)] : reg976[(3'h7):(2'h2)]) ?
                  (wire952[(2'h2):(2'h2)] * $unsigned(reg976[(3'h4):(1'h1)])) : ($signed({(8'hb2),
                      (7'h43)}) < (8'hbc))) ?
              (~|(~reg981)) : reg983);
          if (({$unsigned(($unsigned(reg980) ~^ $unsigned(wire954)))} - wire973))
            begin
              reg987 <= $signed(wire953);
              reg988 <= {reg970[(4'hc):(4'h9)],
                  (wire973[(2'h3):(2'h2)] <<< ($unsigned((~&wire955)) ?
                      wire951 : (reg983[(3'h6):(2'h3)] >= reg968)))};
              reg989 <= (8'hbc);
              reg990 <= reg966;
              reg991 <= reg966;
            end
          else
            begin
              reg987 <= reg969;
              reg988 <= (((~|((!reg977) ?
                      (reg965 ^~ (8'hb5)) : $unsigned(reg981))) <<< reg967) ?
                  $unsigned((-(^~(reg983 ?
                      reg980 : wire953)))) : $signed($signed((reg966[(4'hb):(4'hb)] ?
                      (reg985 + reg984) : (reg983 ? wire974 : reg967)))));
            end
        end
      else
        begin
          if ((reg988 ?
              $signed(reg965) : $signed((($unsigned(reg964) ?
                      (reg988 || (8'ha3)) : (wire959 ? (8'ha8) : reg979)) ?
                  (~(reg982 ? reg987 : reg971)) : {$unsigned(reg979)}))))
            begin
              reg982 <= ((8'hba) ?
                  (reg981[(4'hf):(4'h8)] <= $unsigned((8'hbe))) : reg977[(3'h5):(1'h0)]);
              reg983 <= $signed(wire953);
              reg984 <= reg979[(1'h0):(1'h0)];
              reg985 <= (reg983[(3'h6):(2'h3)] ~^ (|$unsigned(wire957)));
            end
          else
            begin
              reg982 <= ((^reg975) ?
                  ({(|{wire954, wire974}),
                      {(reg986 ?
                              reg982 : reg966)}} + reg961[(4'hc):(3'h4)]) : (+reg977[(2'h2):(1'h0)]));
              reg983 <= (!((-(~(8'ha3))) & ((~^$signed(reg977)) ?
                  $signed(reg981) : (^$signed(wire956)))));
              reg984 <= (reg983 ?
                  reg975[(3'h6):(3'h5)] : $signed((reg963[(3'h5):(2'h3)] >= reg989)));
              reg985 <= reg978[(1'h1):(1'h1)];
              reg986 <= $signed(reg985);
            end
          reg987 <= ({({$unsigned(wire974)} ? $signed(reg983) : (&reg966)),
                  (|((~wire956) ? {wire959, (8'hb4)} : (reg983 > (8'h9d))))} ?
              reg968[(3'h5):(3'h4)] : $unsigned(wire954[(3'h6):(3'h5)]));
          reg988 <= {$signed({{$unsigned(reg977)}, reg963[(2'h2):(1'h0)]})};
          reg989 <= reg971;
        end
    end
  assign wire992 = reg983[(3'h4):(2'h2)];
  assign wire993 = reg988;
  assign wire994 = (reg962 ? (|$unsigned(wire960)) : reg978[(1'h0):(1'h0)]);
  assign wire995 = reg968;
  always
    @(posedge clk) begin
      reg996 <= ((({(wire955 ~^ reg969)} ^~ (reg969 >> $unsigned(reg987))) || ((~^(~^reg978)) ?
              (reg983 >>> {reg991, (8'hae)}) : {$signed(reg963),
                  reg971[(4'ha):(3'h4)]})) ?
          $signed(($signed((reg970 || wire959)) ^~ {reg962[(1'h0):(1'h0)]})) : wire960[(4'hb):(1'h0)]);
      reg997 <= $unsigned(reg989);
    end
  assign wire998 = ((reg963 ?
                       {(wire992 ?
                               $signed(reg961) : wire957[(3'h5):(1'h0)])} : $signed($unsigned($signed(wire955)))) | $unsigned((($signed(reg987) ?
                       wire952[(3'h4):(3'h4)] : (~|wire957)) + $signed(wire959))));
  assign wire999 = ($unsigned(reg989[(1'h1):(1'h0)]) ?
                       reg962[(2'h2):(1'h0)] : reg989[(3'h4):(2'h2)]);
  assign wire1000 = ($signed(reg967[(4'hb):(4'h9)]) | reg961);
  assign wire1001 = reg963;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module562
#( parameter param902 = ((|{{((7'h40) ^~ (8'hb4)), ((7'h42) || (8'hb4))}, (|((8'hb0) ? (8'h9f) : (8'ha8)))}) <= {(~|{((8'hb0) ? (8'hbd) : (8'hae)), ((8'ha2) * (8'hb3))})}) )
(y, clk, wire563, wire564, wire565, wire566);
  output wire [(32'h259):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire563;
  input wire [(5'h14):(1'h0)] wire564;
  input wire [(5'h15):(1'h0)] wire565;
  input wire [(5'h12):(1'h0)] wire566;
  reg signed [(3'h4):(1'h0)] reg901 = (1'h0);
  reg [(4'ha):(1'h0)] reg900 = (1'h0);
  reg [(3'h6):(1'h0)] reg899 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg898 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg897 = (1'h0);
  reg [(3'h5):(1'h0)] reg896 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg895 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg894 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg893 = (1'h0);
  reg [(5'h15):(1'h0)] reg892 = (1'h0);
  reg [(4'hc):(1'h0)] reg891 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg890 = (1'h0);
  reg [(3'h6):(1'h0)] reg889 = (1'h0);
  reg [(4'h8):(1'h0)] reg888 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg887 = (1'h0);
  reg [(3'h6):(1'h0)] reg886 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg885 = (1'h0);
  wire [(3'h7):(1'h0)] wire884;
  wire signed [(4'ha):(1'h0)] wire883;
  reg [(5'h13):(1'h0)] reg882 = (1'h0);
  reg [(5'h11):(1'h0)] reg881 = (1'h0);
  reg [(5'h11):(1'h0)] reg880 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg879 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg878 = (1'h0);
  reg [(3'h6):(1'h0)] reg877 = (1'h0);
  reg [(4'hb):(1'h0)] reg876 = (1'h0);
  wire [(4'ha):(1'h0)] wire875;
  wire signed [(3'h7):(1'h0)] wire874;
  reg signed [(4'hc):(1'h0)] reg873 = (1'h0);
  reg [(5'h12):(1'h0)] reg872 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg871 = (1'h0);
  reg [(4'hc):(1'h0)] reg870 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg869 = (1'h0);
  reg [(2'h3):(1'h0)] reg868 = (1'h0);
  reg [(4'hb):(1'h0)] reg867 = (1'h0);
  reg [(4'hf):(1'h0)] reg866 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg865 = (1'h0);
  reg [(5'h13):(1'h0)] reg864 = (1'h0);
  reg [(4'hd):(1'h0)] reg863 = (1'h0);
  reg [(5'h15):(1'h0)] reg862 = (1'h0);
  reg [(5'h12):(1'h0)] reg861 = (1'h0);
  reg signed [(4'he):(1'h0)] reg860 = (1'h0);
  wire [(2'h2):(1'h0)] wire859;
  wire signed [(4'h8):(1'h0)] wire858;
  wire signed [(4'hf):(1'h0)] wire670;
  wire [(5'h14):(1'h0)] wire672;
  wire [(5'h12):(1'h0)] wire673;
  wire signed [(5'h14):(1'h0)] wire674;
  wire signed [(4'hb):(1'h0)] wire758;
  wire signed [(5'h12):(1'h0)] wire760;
  wire [(4'ha):(1'h0)] wire761;
  wire signed [(5'h12):(1'h0)] wire762;
  wire signed [(3'h7):(1'h0)] wire763;
  wire signed [(5'h11):(1'h0)] wire856;
  assign y = {reg901,
                 reg900,
                 reg899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 reg893,
                 reg892,
                 reg891,
                 reg890,
                 reg889,
                 reg888,
                 reg887,
                 reg886,
                 reg885,
                 wire884,
                 wire883,
                 reg882,
                 reg881,
                 reg880,
                 reg879,
                 reg878,
                 reg877,
                 reg876,
                 wire875,
                 wire874,
                 reg873,
                 reg872,
                 reg871,
                 reg870,
                 reg869,
                 reg868,
                 reg867,
                 reg866,
                 reg865,
                 reg864,
                 reg863,
                 reg862,
                 reg861,
                 reg860,
                 wire859,
                 wire858,
                 wire670,
                 wire672,
                 wire673,
                 wire674,
                 wire758,
                 wire760,
                 wire761,
                 wire762,
                 wire763,
                 wire856,
                 (1'h0)};
  module567 modinst671 (.wire572((8'hb6)), .wire568(wire565), .wire570(wire563), .wire571(wire566), .wire569(wire564), .clk(clk), .y(wire670));
  assign wire672 = wire563[(2'h3):(1'h1)];
  assign wire673 = (+($unsigned($signed({wire565, wire672})) ?
                       wire563[(3'h5):(2'h2)] : $signed($signed((wire563 ?
                           wire672 : wire563)))));
  assign wire674 = {($signed((~|$unsigned(wire565))) >>> wire565[(4'hb):(4'hb)]),
                       $unsigned(wire565)};
  module675 modinst759 (.wire676(wire564), .wire679(wire673), .clk(clk), .wire677(wire670), .wire678(wire674), .y(wire758));
  assign wire760 = $unsigned(wire758[(3'h4):(2'h3)]);
  assign wire761 = $unsigned(wire564[(5'h14):(4'h8)]);
  assign wire762 = (^~$unsigned(wire564));
  assign wire763 = (8'ha4);
  module764 modinst857 (wire856, clk, wire758, wire762, wire672, wire566, wire760);
  assign wire858 = (|wire674[(3'h4):(1'h0)]);
  assign wire859 = (-wire672[(5'h13):(2'h3)]);
  always
    @(posedge clk) begin
      reg860 <= ({(wire858[(3'h5):(1'h1)] ?
                  $unsigned($signed(wire760)) : $signed((wire563 | wire566))),
              wire760[(4'hd):(3'h4)]} ?
          wire762[(3'h4):(1'h0)] : ((~($signed((7'h44)) ?
              $unsigned(wire673) : (wire673 ? wire565 : wire566))) != wire758));
      reg861 <= $signed((wire673 >= wire760[(4'he):(3'h4)]));
      if ($signed({($unsigned(wire673[(4'h9):(4'h9)]) ?
              ((+wire762) * $unsigned(reg861)) : wire565)}))
        begin
          reg862 <= (($unsigned(($unsigned(reg861) ?
                  wire670[(3'h6):(3'h6)] : (^~wire565))) ?
              ($signed(wire762) != (&wire672[(1'h0):(1'h0)])) : $signed($unsigned($unsigned(wire672)))) - $signed((((~wire670) ?
              {(8'ha6)} : $signed(wire762)) == wire564[(5'h13):(3'h5)])));
          reg863 <= (8'hb5);
          reg864 <= wire856[(3'h7):(1'h0)];
          if ((reg863 & reg863))
            begin
              reg865 <= $unsigned((^~reg861[(3'h5):(1'h0)]));
              reg866 <= $unsigned(((($unsigned(wire758) ?
                          (reg861 ? (8'ha4) : wire858) : (wire674 ?
                              wire758 : wire858)) ?
                      $signed($signed(wire673)) : wire566[(4'he):(3'h4)]) ?
                  ($signed((wire762 ^ reg862)) && (~&{wire563})) : wire761[(2'h3):(2'h3)]));
            end
          else
            begin
              reg865 <= $signed($unsigned(($signed(wire672[(2'h3):(2'h3)]) ?
                  $signed((wire858 ?
                      wire859 : wire858)) : (~|(wire760 << wire763)))));
              reg866 <= wire670;
              reg867 <= {reg864[(4'he):(2'h2)]};
              reg868 <= (($signed($unsigned((wire566 * wire670))) << {{$unsigned(reg862)}}) ?
                  wire856 : reg865);
              reg869 <= wire763;
            end
          reg870 <= wire761;
        end
      else
        begin
          reg862 <= (!((~|wire856[(4'hc):(4'h9)]) >>> wire565));
          reg863 <= (~|$unsigned(wire758));
          if (($signed(reg869[(1'h1):(1'h1)]) && (|reg864)))
            begin
              reg864 <= (&(((!(wire564 ? reg864 : reg863)) ?
                      ($signed(reg866) <= (wire856 && reg867)) : wire563[(4'h9):(4'h9)]) ?
                  (reg860[(4'hd):(3'h7)] ?
                      reg867[(4'h9):(3'h5)] : {wire856}) : (^wire856[(3'h5):(3'h5)])));
              reg865 <= (|$unsigned(reg863));
              reg866 <= $unsigned((-wire758));
              reg867 <= (((-$signed({reg870})) <<< $signed((wire565 != wire858[(2'h3):(2'h2)]))) ?
                  wire566[(4'h8):(4'h8)] : wire566[(3'h4):(3'h4)]);
            end
          else
            begin
              reg864 <= $signed(((~|(~|(^~wire760))) << reg863[(4'hb):(4'h9)]));
              reg865 <= wire672[(5'h13):(4'he)];
              reg866 <= (wire673[(2'h2):(2'h2)] ?
                  ((!(^~$signed(wire673))) | (|((reg870 != (8'hbb)) || (wire762 ?
                      wire859 : wire674)))) : $unsigned({({wire763,
                          wire856} >= (reg867 >= wire670)),
                      $unsigned(wire565[(4'ha):(3'h6)])}));
              reg867 <= reg860[(4'h8):(4'h8)];
            end
          reg868 <= ((|($unsigned({reg867,
              wire762}) || wire673[(4'ha):(4'ha)])) <<< $unsigned($unsigned(reg863)));
        end
      reg871 <= $signed(($unsigned($unsigned((reg862 ? (8'ha3) : wire761))) ?
          reg865 : $signed(wire566[(4'hb):(4'h8)])));
      if ((~|$unsigned(wire762[(4'h8):(1'h0)])))
        begin
          reg872 <= $signed(((&wire674[(2'h3):(2'h3)]) <<< wire565[(4'hd):(4'hc)]));
        end
      else
        begin
          reg872 <= $unsigned((($signed($unsigned(wire856)) >= $signed((~reg871))) ?
              reg861 : ({$unsigned((8'ha8)), (~^wire566)} ?
                  reg871[(3'h7):(3'h5)] : wire858)));
          reg873 <= wire858;
        end
    end
  assign wire874 = reg864;
  assign wire875 = $signed($signed((+(+(reg869 ? wire762 : wire859)))));
  always
    @(posedge clk) begin
      if ((wire856[(4'hd):(3'h6)] ?
          (~&reg867[(3'h7):(2'h2)]) : ((wire859[(2'h2):(2'h2)] ?
              {$signed(reg872),
                  (reg870 && wire673)} : (|wire565[(4'hc):(2'h2)])) + wire670)))
        begin
          reg876 <= ($signed((8'hb1)) << reg861);
          reg877 <= ($signed({$signed((wire672 != wire874)),
                  wire674[(4'hc):(1'h0)]}) ?
              (wire874[(3'h7):(3'h5)] | reg867) : (wire875[(4'ha):(1'h1)] >> reg864));
          if (wire674)
            begin
              reg878 <= $unsigned($unsigned(($signed($signed(wire760)) ?
                  wire856[(3'h5):(2'h3)] : (!(!wire874)))));
              reg879 <= ($signed((reg866[(3'h5):(2'h2)] < (((8'haa) >>> reg865) ?
                  (&reg869) : ((8'h9f) ^~ reg869)))) > (&reg864));
              reg880 <= $unsigned({reg871,
                  ($unsigned(wire670[(1'h1):(1'h0)]) || ($signed(wire875) < (reg869 != (7'h42))))});
              reg881 <= reg861;
              reg882 <= $unsigned((~wire761[(3'h5):(2'h2)]));
            end
          else
            begin
              reg878 <= {$unsigned((!$signed((&reg878)))),
                  ($unsigned($unsigned($signed(wire758))) ?
                      $unsigned(({wire858, reg869} ?
                          reg869 : reg871)) : ((!$unsigned(reg866)) & ((wire763 ~^ reg873) <<< ((8'ha5) ?
                          wire670 : reg872))))};
              reg879 <= {($signed($signed(wire874)) ^ reg865),
                  $unsigned({wire760})};
              reg880 <= {reg862, (&(7'h44))};
              reg881 <= (8'hbb);
            end
        end
      else
        begin
          reg876 <= (^{reg881});
          if ($signed($unsigned($signed(wire856))))
            begin
              reg877 <= $unsigned($unsigned(wire761[(2'h2):(2'h2)]));
              reg878 <= $signed($unsigned($signed($unsigned((reg871 ?
                  reg869 : reg871)))));
              reg879 <= $signed({wire672, {$unsigned({wire565})}});
              reg880 <= ((wire670[(4'h8):(3'h6)] ?
                      $signed((8'hbc)) : (($signed(wire670) ?
                              (|reg870) : $unsigned(wire762)) ?
                          (((8'hb0) >= reg878) && (reg877 <= reg880)) : (-(wire762 ?
                              reg877 : wire856)))) ?
                  {wire674,
                      $unsigned($unsigned((reg862 << reg862)))} : wire858[(4'h8):(1'h1)]);
              reg881 <= $signed(reg877);
            end
          else
            begin
              reg877 <= ($signed((((^~reg861) - $unsigned(reg863)) ?
                  $unsigned($signed(wire674)) : reg882)) && $signed($signed((-(&wire674)))));
            end
          reg882 <= (~^({(((8'hb9) ?
                  wire563 : reg873) < reg867[(4'h9):(3'h7)])} << {(!(^~(8'hba))),
              reg865[(3'h5):(3'h5)]}));
        end
    end
  assign wire883 = $unsigned($signed((~&((~&wire565) ?
                       $unsigned(wire856) : $unsigned(reg862)))));
  assign wire884 = (-($signed($unsigned((reg867 ?
                       wire565 : (8'hb6)))) + $signed(reg866[(3'h5):(1'h0)])));
  always
    @(posedge clk) begin
      if ((((~reg868) ?
          reg868 : (((&wire673) && wire670[(3'h6):(3'h4)]) ?
              (~^wire672[(3'h4):(1'h0)]) : ($unsigned(reg864) ?
                  (reg864 >= (8'ha2)) : $signed(reg867)))) << ({(~|{reg861})} ?
          ($unsigned($unsigned(wire856)) ?
              ((~&wire761) ^ $unsigned((8'ha3))) : {{reg881},
                  (reg879 < wire858)}) : {((wire563 - (8'haf)) ?
                  reg868 : reg867[(3'h6):(2'h3)])})))
        begin
          if (((wire565 <= reg868[(1'h0):(1'h0)]) == $signed((reg876[(4'h8):(1'h1)] | $unsigned((reg863 ?
              wire874 : reg865))))))
            begin
              reg885 <= ((8'hbf) && (8'ha0));
              reg886 <= reg871;
            end
          else
            begin
              reg885 <= (~^((wire674 & $signed((reg877 ^ (8'hbf)))) ?
                  (&(wire564 ?
                      wire670[(3'h5):(1'h1)] : reg862[(4'he):(4'h9)])) : wire858));
              reg886 <= reg860[(3'h5):(1'h1)];
            end
        end
      else
        begin
          reg885 <= $signed($signed(($unsigned(((7'h42) <<< reg862)) ?
              ($signed(wire874) && ((8'ha5) << reg882)) : reg878[(3'h6):(3'h6)])));
          reg886 <= {reg868[(2'h2):(1'h1)],
              $signed(($unsigned((reg879 >= reg864)) < ($signed((8'ha9)) | $unsigned(wire564))))};
          reg887 <= (reg886 ?
              wire674[(4'hf):(3'h4)] : $unsigned((($signed(wire874) < (reg871 ?
                      wire672 : wire674)) ?
                  reg864 : (!(+reg869)))));
          if ($unsigned(((wire762[(1'h1):(1'h1)] << ($unsigned((8'h9c)) ?
              reg878 : (reg877 ? wire859 : wire859))) | $signed(reg886))))
            begin
              reg888 <= wire670;
              reg889 <= reg887[(2'h3):(1'h0)];
              reg890 <= (!$unsigned({(reg889[(3'h4):(1'h0)] && reg880[(4'h8):(3'h4)]),
                  wire763}));
              reg891 <= (!reg889);
            end
          else
            begin
              reg888 <= wire760;
              reg889 <= reg873;
              reg890 <= (reg872 ?
                  (wire565[(5'h11):(5'h10)] ?
                      (wire762[(3'h5):(3'h5)] ?
                          reg878 : wire856[(2'h3):(2'h3)]) : reg870[(4'hc):(4'h9)]) : {$signed($signed(reg878))});
            end
          reg892 <= (($unsigned((wire761[(3'h4):(3'h4)] ?
                  {reg860} : (reg888 + wire874))) ?
              $unsigned(reg881) : ($unsigned((wire762 >>> wire883)) - reg861)) & (reg870 >> {reg871,
              (8'hae)}));
        end
      reg893 <= ($unsigned($signed(((reg866 * reg866) ?
          (reg865 != (8'hb1)) : reg865))) >>> wire884[(2'h2):(1'h0)]);
      if ((wire856 >= $signed(($signed($unsigned(reg888)) <= $unsigned($unsigned(wire883))))))
        begin
          reg894 <= $unsigned((wire761 - reg879));
          reg895 <= ($signed((~|reg861[(4'h8):(3'h7)])) ~^ $unsigned({$unsigned((!reg864)),
              $unsigned((wire758 ? wire565 : reg877))}));
          if (((reg890 >>> wire566[(3'h5):(2'h3)]) <= {((reg869[(3'h5):(2'h2)] ?
                  wire674 : reg863) & wire673[(5'h12):(2'h2)])}))
            begin
              reg896 <= $signed(reg886);
              reg897 <= reg886;
              reg898 <= (~&(!$unsigned($signed((~wire875)))));
              reg899 <= {{$unsigned(reg896), (8'ha2)}};
            end
          else
            begin
              reg896 <= reg867;
              reg897 <= (reg870 ?
                  {$unsigned($unsigned($unsigned(reg894))),
                      $signed((!{(8'hab)}))} : $unsigned($signed(wire566[(4'hd):(2'h3)])));
            end
        end
      else
        begin
          reg894 <= ($unsigned((-reg889)) ?
              wire763 : (^$unsigned(($signed(reg889) <<< wire563))));
          reg895 <= ($unsigned($signed((+(reg870 ?
              (7'h40) : reg862)))) || reg861[(3'h6):(3'h5)]);
        end
      reg900 <= ((reg890 ?
          $signed((~&(wire674 || wire875))) : $signed((+$signed(reg882)))) != reg868[(2'h2):(1'h1)]);
      reg901 <= ((|$unsigned(reg900[(1'h0):(1'h0)])) != wire563);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module764  (y, clk, wire769, wire768, wire767, wire766, wire765);
  output wire [(32'h108):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire769;
  input wire [(4'h8):(1'h0)] wire768;
  input wire [(5'h14):(1'h0)] wire767;
  input wire [(5'h10):(1'h0)] wire766;
  input wire [(4'he):(1'h0)] wire765;
  wire signed [(4'hb):(1'h0)] wire854;
  reg signed [(3'h7):(1'h0)] reg791 = (1'h0);
  reg [(4'h9):(1'h0)] reg790 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg789 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg788 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg787 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg786 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg785 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg784 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg783 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg782 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg781 = (1'h0);
  reg [(5'h15):(1'h0)] reg780 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg779 = (1'h0);
  reg [(3'h7):(1'h0)] reg778 = (1'h0);
  reg [(3'h5):(1'h0)] reg777 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg776 = (1'h0);
  reg [(2'h2):(1'h0)] reg775 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg774 = (1'h0);
  reg [(5'h14):(1'h0)] reg773 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg772 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire771;
  wire signed [(5'h10):(1'h0)] wire770;
  assign y = {wire854,
                 reg791,
                 reg790,
                 reg789,
                 reg788,
                 reg787,
                 reg786,
                 reg785,
                 reg784,
                 reg783,
                 reg782,
                 reg781,
                 reg780,
                 reg779,
                 reg778,
                 reg777,
                 reg776,
                 reg775,
                 reg774,
                 reg773,
                 reg772,
                 wire771,
                 wire770,
                 (1'h0)};
  assign wire770 = {wire768, (8'hb8)};
  assign wire771 = wire765;
  always
    @(posedge clk) begin
      reg772 <= ({wire768[(4'h8):(3'h4)],
          wire767[(5'h10):(4'hb)]} ~^ $signed(($signed(wire767[(5'h14):(1'h1)]) << wire767[(3'h5):(1'h0)])));
      reg773 <= wire769;
      if ((wire768[(3'h5):(1'h1)] ?
          ($signed((wire765 <= (wire765 * reg772))) || reg773) : ($signed(wire766[(3'h6):(3'h5)]) ?
              (&{(~&(8'haa))}) : ($unsigned($signed(wire771)) ?
                  $signed(wire765[(2'h2):(1'h1)]) : (|wire769)))))
        begin
          reg774 <= {(-(8'haa))};
        end
      else
        begin
          if (reg773)
            begin
              reg774 <= wire769;
              reg775 <= (+(!$unsigned((~^$unsigned(reg774)))));
              reg776 <= (~^$signed(reg774[(4'ha):(3'h7)]));
              reg777 <= ((8'hb8) << (wire765[(3'h7):(1'h1)] ?
                  {({wire769, reg776} < wire765[(4'h8):(3'h4)]),
                      wire766} : (wire766 ^ wire766)));
            end
          else
            begin
              reg774 <= reg775[(1'h1):(1'h1)];
              reg775 <= (!wire767);
            end
          reg778 <= ((((!((8'hbc) ~^ wire766)) | $signed((8'hb8))) ~^ $signed(((~&wire770) ?
                  (wire769 >> wire768) : ((7'h40) ? wire766 : reg776)))) ?
              reg777 : wire770[(3'h4):(3'h4)]);
          reg779 <= (+$signed($unsigned($signed((8'hbe)))));
          reg780 <= {({(-$unsigned(reg777))} <= reg779[(5'h11):(4'h9)])};
        end
      if ({$signed((|{wire767[(4'h8):(3'h7)], ((8'ha9) ? (8'h9f) : wire767)})),
          ($signed({reg775, (!wire770)}) <<< $signed($signed(reg775)))})
        begin
          if (($signed((((8'h9f) ? $signed((8'ha4)) : reg779[(3'h5):(1'h1)]) ?
              (^~wire770) : (^wire765))) != ($unsigned((^~wire771[(2'h3):(2'h2)])) - ((((8'hae) || reg773) ?
                  {reg778, wire771} : $unsigned(wire770)) ?
              $signed(reg772) : (^(wire766 ? wire771 : wire771))))))
            begin
              reg781 <= (^reg780[(1'h0):(1'h0)]);
              reg782 <= (~reg772);
              reg783 <= wire770[(1'h1):(1'h0)];
              reg784 <= ((~&({$signed(reg782)} >> {(reg781 && reg776)})) <= ((~wire767) ?
                  $signed((reg781[(1'h1):(1'h1)] & wire768)) : ($signed((wire768 ?
                      reg775 : reg781)) << $unsigned($unsigned(reg778)))));
            end
          else
            begin
              reg781 <= (~&$unsigned({{(|wire767)}, (|{reg774, reg773})}));
            end
          reg785 <= (reg779[(2'h3):(1'h1)] >= (8'haa));
          reg786 <= {wire771};
          if ((^$signed((|$unsigned(reg773[(4'hc):(4'h8)])))))
            begin
              reg787 <= {reg774};
              reg788 <= ((reg787 ?
                  (wire770 == $signed($unsigned(reg783))) : $unsigned(((wire767 >>> (8'hb0)) & (reg782 ?
                      reg776 : reg774)))) * (&(~&$signed($signed(wire771)))));
            end
          else
            begin
              reg787 <= ((($unsigned((wire770 || reg776)) ?
                          (wire768[(3'h7):(3'h6)] ?
                              (reg788 <<< reg788) : (~|reg777)) : $unsigned(reg785)) ?
                      (reg788[(4'h9):(3'h7)] ?
                          {$unsigned(reg787),
                              (+reg785)} : (~reg777[(2'h3):(1'h0)])) : reg782) ?
                  (((~$signed(reg782)) ?
                      (wire765 ?
                          reg776[(1'h1):(1'h1)] : $unsigned(reg788)) : ((+wire770) + $unsigned(reg774))) <<< (^~wire771[(2'h3):(1'h0)])) : wire771);
              reg788 <= (((!{(wire765 ? reg788 : reg774), $signed(reg777)}) ?
                  $signed(reg775) : ($unsigned(reg788[(1'h1):(1'h0)]) ?
                      {(wire765 * reg777),
                          $unsigned(reg779)} : reg783[(2'h2):(1'h1)])) * $unsigned($signed($unsigned($signed(wire768)))));
              reg789 <= ($unsigned((((reg781 ? wire766 : wire766) ?
                      ((7'h41) ? wire765 : reg787) : reg783[(4'hf):(2'h3)]) ?
                  ($unsigned(reg778) | (&(8'hb1))) : (^reg782))) >>> wire770[(4'ha):(3'h7)]);
              reg790 <= ({(wire765 ?
                      {{wire770}} : (-$signed(reg787)))} ^~ (reg781 & (reg786 >>> ($unsigned((7'h41)) ?
                  reg784 : {wire769, reg785}))));
              reg791 <= ($signed(reg779) ^ (-reg782[(3'h5):(2'h3)]));
            end
        end
      else
        begin
          reg781 <= ($signed((({wire766} ?
                  $unsigned(reg781) : wire766[(4'hf):(1'h1)]) ^ $signed((reg783 ?
                  wire770 : (8'hb0))))) ?
              {(|($unsigned(reg779) >= $unsigned(reg786))),
                  (|$unsigned((8'ha8)))} : (~&{$signed(reg772[(1'h1):(1'h0)])}));
          if ((reg791 ? reg787 : reg780[(1'h0):(1'h0)]))
            begin
              reg782 <= ((~|(~$unsigned(((8'hbf) == wire769)))) ?
                  $unsigned((reg780 ?
                      reg785[(3'h7):(3'h7)] : reg783)) : ($unsigned(reg784) ^~ $signed($unsigned(wire770[(4'hb):(1'h0)]))));
            end
          else
            begin
              reg782 <= $signed((^wire769));
              reg783 <= (((~|reg778[(1'h1):(1'h1)]) < (~&(^(reg790 ?
                      reg791 : reg776)))) ?
                  {((~^(wire766 ? reg789 : reg774)) ?
                          {(8'had)} : (~^{wire766,
                              reg773}))} : $signed(((~|reg789) ^ $unsigned({reg786}))));
            end
          if ((((reg782 > reg785[(1'h1):(1'h1)]) | $signed(reg772)) + (^~(+reg772[(2'h2):(1'h0)]))))
            begin
              reg784 <= ({(~^((reg778 ? reg782 : reg775) ?
                      (~^reg790) : (8'ha7))),
                  (8'ha7)} * (reg791[(3'h4):(2'h2)] >>> ($unsigned((reg784 ?
                  reg775 : reg774)) * ($unsigned(reg782) >> {(8'hbc),
                  wire769}))));
              reg785 <= (((+(reg777 ? $unsigned(wire765) : $unsigned(reg776))) ?
                      ((+((8'ha5) ^~ wire767)) ?
                          (!$unsigned((8'ha4))) : reg787) : $signed({(reg779 ?
                              wire768 : wire769)})) ?
                  ({reg788, {wire766}} | wire769[(3'h4):(1'h1)]) : reg779);
            end
          else
            begin
              reg784 <= {($signed({(reg776 ? wire767 : (8'hb7)),
                      reg781}) < (^reg772[(1'h0):(1'h0)])),
                  reg775};
              reg785 <= ({$signed((~(reg782 ? reg786 : (8'hbd))))} ?
                  reg777 : ($signed(reg772[(1'h0):(1'h0)]) - wire767));
              reg786 <= reg791;
              reg787 <= ($signed((-($unsigned(reg785) >>> reg786))) ?
                  $signed(reg787) : ((&$unsigned($signed(wire767))) ?
                      reg787[(4'h8):(3'h4)] : (wire766 ^ $unsigned(wire770))));
            end
          reg788 <= reg779[(3'h6):(3'h5)];
          reg789 <= (reg785[(4'ha):(3'h6)] ?
              $unsigned(reg784) : $unsigned($unsigned(((reg788 || reg782) ?
                  (8'hbb) : (&reg788)))));
        end
    end
  module792 modinst855 (wire854, clk, reg773, reg776, reg779, reg784);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module675  (y, clk, wire679, wire678, wire677, wire676);
  output wire [(32'h195):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire679;
  input wire [(5'h13):(1'h0)] wire678;
  input wire signed [(2'h3):(1'h0)] wire677;
  input wire [(5'h11):(1'h0)] wire676;
  wire signed [(5'h15):(1'h0)] wire757;
  wire signed [(3'h4):(1'h0)] wire756;
  wire [(5'h12):(1'h0)] wire755;
  wire signed [(3'h6):(1'h0)] wire754;
  wire [(4'hd):(1'h0)] wire753;
  reg signed [(3'h7):(1'h0)] reg752 = (1'h0);
  reg [(4'h8):(1'h0)] reg751 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg750 = (1'h0);
  reg [(4'h8):(1'h0)] reg749 = (1'h0);
  reg [(4'hc):(1'h0)] reg748 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg747 = (1'h0);
  reg [(3'h4):(1'h0)] reg746 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg745 = (1'h0);
  reg [(5'h14):(1'h0)] reg744 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg743 = (1'h0);
  reg [(4'ha):(1'h0)] reg742 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg741 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg740 = (1'h0);
  reg [(5'h10):(1'h0)] reg739 = (1'h0);
  reg [(3'h6):(1'h0)] reg738 = (1'h0);
  reg [(4'ha):(1'h0)] reg737 = (1'h0);
  reg [(4'hf):(1'h0)] reg736 = (1'h0);
  reg [(2'h2):(1'h0)] reg735 = (1'h0);
  reg [(3'h6):(1'h0)] reg734 = (1'h0);
  reg signed [(4'he):(1'h0)] reg733 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg732 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg731 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg730 = (1'h0);
  reg [(5'h11):(1'h0)] reg729 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg728 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire727;
  wire [(4'hd):(1'h0)] wire726;
  wire [(3'h7):(1'h0)] wire725;
  wire signed [(4'he):(1'h0)] wire724;
  wire [(4'h8):(1'h0)] wire722;
  wire signed [(4'hf):(1'h0)] wire682;
  wire [(3'h6):(1'h0)] wire681;
  wire signed [(3'h7):(1'h0)] wire680;
  assign y = {wire757,
                 wire756,
                 wire755,
                 wire754,
                 wire753,
                 reg752,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 reg747,
                 reg746,
                 reg745,
                 reg744,
                 reg743,
                 reg742,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 reg730,
                 reg729,
                 reg728,
                 wire727,
                 wire726,
                 wire725,
                 wire724,
                 wire722,
                 wire682,
                 wire681,
                 wire680,
                 (1'h0)};
  assign wire680 = wire677;
  assign wire681 = (({(^~(-wire677))} << ($unsigned((wire678 ?
                           wire678 : wire680)) >>> ((wire676 ?
                           wire678 : wire679) << wire679[(3'h4):(1'h1)]))) ?
                       {($unsigned({wire677}) * wire678)} : wire678);
  assign wire682 = (~|$unsigned((wire681 != wire681)));
  module683 modinst723 (wire722, clk, wire682, wire676, wire678, wire679);
  assign wire724 = (({(!((8'hb4) ? wire678 : wire678)), (+wire677)} ?
                           wire678 : $signed(wire677[(1'h1):(1'h0)])) ?
                       (((wire678 ~^ (wire681 == wire722)) ?
                           wire677 : ((wire682 - wire680) - {wire722,
                               wire682})) * $unsigned($unsigned(((8'hbe) + wire681)))) : wire722);
  assign wire725 = ((!(wire724 ?
                           $signed({wire677, wire677}) : ((wire676 ?
                               wire676 : wire724) >> wire676[(2'h3):(2'h3)]))) ?
                       (^$signed($signed(wire724))) : $unsigned($signed({$unsigned(wire677),
                           wire677[(1'h1):(1'h0)]})));
  assign wire726 = $signed($unsigned((wire681[(2'h3):(2'h3)] ?
                       (wire724[(4'hd):(4'h8)] ?
                           wire678 : wire679[(3'h7):(3'h5)]) : ((wire678 ~^ (8'haf)) ?
                           wire680 : $signed((8'haf))))));
  assign wire727 = wire678;
  always
    @(posedge clk) begin
      reg728 <= ($unsigned($signed($signed({wire678,
          wire726}))) || $unsigned((!(wire681 + $signed(wire725)))));
      reg729 <= wire676[(4'h8):(3'h4)];
      reg730 <= ((~$signed(((reg728 ?
          wire678 : wire726) & $signed((8'hae))))) <<< (&(wire681 ?
          (wire722[(3'h7):(1'h0)] || $unsigned(reg728)) : ({wire682, reg728} ?
              (&reg728) : wire727))));
    end
  always
    @(posedge clk) begin
      if (((wire680[(2'h2):(1'h1)] << (((^~wire682) <= wire676) ?
              $unsigned(reg728[(3'h7):(3'h7)]) : reg728)) ?
          (!wire680[(1'h1):(1'h1)]) : ((~^$unsigned(wire679[(4'hf):(3'h4)])) >>> $signed(wire722))))
        begin
          reg731 <= wire724;
          reg732 <= $signed(wire679);
          reg733 <= ($unsigned($unsigned((-((8'hb9) ? (8'h9e) : wire677)))) ?
              (reg728[(3'h4):(3'h4)] * (!{{wire727,
                      (8'hb0)}})) : {(-$unsigned(((8'hae) >>> reg731)))});
          reg734 <= (8'ha6);
          reg735 <= {(+(($unsigned(wire725) ?
                  (wire680 < wire725) : (-reg730)) >> $signed(reg729[(2'h3):(2'h3)])))};
        end
      else
        begin
          reg731 <= (~^((8'ha6) ? (&reg730) : $signed((8'haf))));
          reg732 <= wire676;
          if ({$unsigned(reg735[(1'h0):(1'h0)]), wire676})
            begin
              reg733 <= wire680[(3'h5):(3'h4)];
              reg734 <= wire677[(2'h3):(1'h0)];
              reg735 <= (~((wire722 ?
                  reg728[(1'h0):(1'h0)] : $signed({reg731,
                      wire727})) ^ reg731));
            end
          else
            begin
              reg733 <= $unsigned(wire680[(3'h5):(3'h5)]);
            end
          reg736 <= $unsigned((7'h44));
          if ((~reg729))
            begin
              reg737 <= reg731;
              reg738 <= wire680[(2'h2):(2'h2)];
            end
          else
            begin
              reg737 <= (({(!wire724)} ?
                  (~^(wire681 == reg737[(4'ha):(4'h8)])) : ($unsigned(reg733) ~^ (+((8'ha6) && wire725)))) >>> (~|$signed((~^$unsigned(wire727)))));
              reg738 <= $signed((-$signed(((8'hb3) ?
                  (wire680 ? wire678 : (8'ha3)) : $signed(wire725)))));
              reg739 <= {(({reg729, ((7'h41) ? reg729 : wire722)} ?
                      reg738 : ((reg735 ? reg734 : wire722) ?
                          wire680 : $signed(wire676))) & $signed(($signed(reg729) == $signed(reg736)))),
                  ($signed($signed(reg729)) ~^ $signed((wire677 & $unsigned(reg738))))};
              reg740 <= (reg730 ?
                  $unsigned($unsigned($signed(wire722))) : {{{(reg738 ?
                                  reg732 : (8'ha6)),
                              $unsigned(wire680)}},
                      $signed(((reg735 >> wire678) != wire722[(4'h8):(3'h6)]))});
              reg741 <= (&(($unsigned((|wire680)) * (8'hb3)) ?
                  {(^(wire727 <<< (8'hb7))),
                      ($unsigned(reg734) ?
                          ((8'hb5) << wire725) : $unsigned((7'h44)))} : reg735));
            end
        end
      reg742 <= (reg738[(3'h5):(3'h5)] ?
          $unsigned(($signed(wire726) ?
              $signed((reg732 ?
                  reg730 : (8'ha1))) : (!(reg735 ~^ reg733)))) : ($signed(wire678[(3'h4):(2'h3)]) && $signed(($unsigned(reg729) ?
              $unsigned((8'hb6)) : $signed(wire676)))));
      if ($signed(wire682))
        begin
          reg743 <= $signed(wire676);
        end
      else
        begin
          reg743 <= $unsigned(reg743);
          reg744 <= wire725[(1'h1):(1'h1)];
          if (($unsigned((!($signed(reg729) < (wire681 + reg730)))) ?
              ((reg739 >>> ((wire677 ~^ reg734) ?
                      $signed(wire682) : (reg740 ~^ reg743))) ?
                  ($unsigned((~^(8'hb7))) | (^(reg732 <= reg735))) : (reg740 ?
                      reg744 : ($signed(wire727) ?
                          wire722[(2'h3):(2'h2)] : $unsigned(wire678)))) : (8'hb6)))
            begin
              reg745 <= $unsigned(wire727);
            end
          else
            begin
              reg745 <= ((&(((reg743 << reg728) ?
                      wire676 : (7'h42)) < (reg738[(2'h3):(2'h2)] ?
                      reg744 : ((8'hb6) ? reg737 : wire678)))) ?
                  $unsigned(reg734[(3'h6):(1'h0)]) : (8'h9f));
              reg746 <= {(!reg742[(3'h5):(3'h4)])};
              reg747 <= $signed(reg744[(5'h10):(4'h8)]);
              reg748 <= wire682;
            end
          if ($signed({(^~{wire682[(1'h1):(1'h1)], (!wire679)})}))
            begin
              reg749 <= $signed(wire726);
            end
          else
            begin
              reg749 <= {(8'ha2)};
              reg750 <= ($signed(($unsigned($unsigned((8'hb3))) ?
                      $unsigned((^(7'h42))) : $signed($unsigned(wire681)))) ?
                  (!wire726[(1'h1):(1'h0)]) : $unsigned({$signed(reg743[(1'h0):(1'h0)]),
                      $unsigned(reg748[(4'ha):(4'h9)])}));
              reg751 <= (wire678[(5'h13):(2'h3)] != (reg748[(3'h5):(3'h4)] <= ({{reg732}} ?
                  (+wire682) : (wire724 & (!reg740)))));
            end
          reg752 <= reg746[(2'h3):(1'h1)];
        end
    end
  assign wire753 = $unsigned(reg734[(1'h1):(1'h1)]);
  assign wire754 = reg728;
  assign wire755 = $signed($unsigned((wire678[(4'hd):(1'h1)] <= reg730)));
  assign wire756 = $unsigned($signed((8'hac)));
  assign wire757 = {(~^(~&reg743[(3'h4):(1'h0)])),
                       ((+$unsigned(reg730[(2'h2):(2'h2)])) < ((^~$unsigned(reg741)) - ({reg736,
                               (8'hb1)} ?
                           ((8'hab) - wire677) : $unsigned((8'haf)))))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module567  (y, clk, wire568, wire569, wire570, wire571, wire572);
  output wire [(32'h159):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire568;
  input wire [(5'h14):(1'h0)] wire569;
  input wire signed [(4'h9):(1'h0)] wire570;
  input wire [(5'h12):(1'h0)] wire571;
  input wire [(3'h7):(1'h0)] wire572;
  wire [(4'hb):(1'h0)] wire669;
  wire [(2'h2):(1'h0)] wire667;
  wire [(4'hf):(1'h0)] wire651;
  wire [(3'h5):(1'h0)] wire650;
  reg signed [(4'he):(1'h0)] reg649 = (1'h0);
  reg [(4'h8):(1'h0)] reg648 = (1'h0);
  reg [(2'h3):(1'h0)] reg647 = (1'h0);
  reg [(3'h7):(1'h0)] reg646 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg645 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg644 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg643 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg642 = (1'h0);
  reg [(5'h13):(1'h0)] reg641 = (1'h0);
  reg [(4'ha):(1'h0)] reg640 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg639 = (1'h0);
  wire signed [(4'he):(1'h0)] wire638;
  wire signed [(4'hf):(1'h0)] wire637;
  wire [(4'hd):(1'h0)] wire636;
  reg signed [(2'h3):(1'h0)] reg635 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg634 = (1'h0);
  reg [(4'h8):(1'h0)] reg633 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg632 = (1'h0);
  reg [(3'h7):(1'h0)] reg631 = (1'h0);
  wire [(5'h10):(1'h0)] wire630;
  wire signed [(4'ha):(1'h0)] wire629;
  wire signed [(4'hc):(1'h0)] wire628;
  wire [(5'h15):(1'h0)] wire573;
  wire [(3'h5):(1'h0)] wire574;
  wire [(4'hc):(1'h0)] wire575;
  wire [(5'h13):(1'h0)] wire576;
  wire [(4'h9):(1'h0)] wire626;
  assign y = {wire669,
                 wire667,
                 wire651,
                 wire650,
                 reg649,
                 reg648,
                 reg647,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 reg642,
                 reg641,
                 reg640,
                 reg639,
                 wire638,
                 wire637,
                 wire636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 wire630,
                 wire629,
                 wire628,
                 wire573,
                 wire574,
                 wire575,
                 wire576,
                 wire626,
                 (1'h0)};
  assign wire573 = wire571[(4'hb):(1'h1)];
  assign wire574 = (wire568 ?
                       $signed(wire570[(3'h4):(2'h3)]) : wire573[(1'h1):(1'h0)]);
  assign wire575 = (&wire569[(1'h1):(1'h0)]);
  assign wire576 = (7'h43);
  module577 modinst627 (.wire582(wire574), .y(wire626), .clk(clk), .wire580(wire571), .wire581(wire570), .wire579(wire573), .wire578(wire568));
  assign wire628 = wire573[(5'h10):(3'h7)];
  assign wire629 = (^{(~|$signed((7'h40)))});
  assign wire630 = ($unsigned(($signed($unsigned(wire626)) ?
                           $signed(((8'hb2) <= (8'ha5))) : (7'h44))) ?
                       wire571[(1'h1):(1'h0)] : wire573[(5'h15):(2'h3)]);
  always
    @(posedge clk) begin
      reg631 <= $signed((wire569[(5'h10):(2'h3)] < ({(wire569 ?
                  wire570 : wire628)} ?
          $unsigned(wire568) : (~&wire574))));
      reg632 <= (~|$unsigned({{$signed(wire568)}}));
      reg633 <= (wire626 + $unsigned(wire574));
      reg634 <= ((~&wire629) ?
          $unsigned(($signed((wire574 ? wire630 : wire571)) ?
              $signed((&reg633)) : wire570[(3'h7):(1'h1)])) : (!wire575));
      reg635 <= (((wire571[(5'h10):(3'h4)] != wire574[(2'h2):(1'h1)]) ^ ($signed($signed(wire629)) ?
          (wire630[(3'h4):(1'h1)] <= wire570[(4'h8):(3'h6)]) : ((|(8'ha8)) ?
              $unsigned(reg632) : wire628))) >>> wire569[(4'hf):(3'h5)]);
    end
  assign wire636 = (~&(~^$signed(((~^wire569) ?
                       (|wire574) : (reg632 ^~ wire628)))));
  assign wire637 = (wire576[(4'h8):(1'h0)] >> $unsigned($unsigned(reg632[(4'h9):(2'h2)])));
  assign wire638 = ($unsigned(reg633) || ((wire576 ?
                       (reg635[(1'h1):(1'h0)] + $unsigned(wire569)) : (-(-wire628))) | ($signed($signed(wire571)) ?
                       wire571[(2'h2):(1'h1)] : $unsigned($unsigned(wire636)))));
  always
    @(posedge clk) begin
      reg639 <= wire571;
      if (wire570[(4'h9):(3'h7)])
        begin
          if ((wire638 ?
              {(8'hbc),
                  $unsigned(wire575[(3'h5):(1'h0)])} : reg632[(5'h12):(4'hb)]))
            begin
              reg640 <= reg631;
              reg641 <= {reg639, (8'had)};
              reg642 <= (~^$signed(reg634));
              reg643 <= $unsigned((reg639[(2'h2):(1'h0)] ?
                  wire570[(1'h1):(1'h0)] : (reg633 || (|{wire638, wire628}))));
              reg644 <= (|{{wire630, (^wire568[(5'h12):(4'ha)])},
                  $signed(wire573[(4'he):(3'h5)])});
            end
          else
            begin
              reg640 <= wire629;
              reg641 <= wire629;
              reg642 <= reg642[(3'h6):(1'h0)];
              reg643 <= {(^~$signed(wire637))};
              reg644 <= reg631;
            end
          reg645 <= reg641;
          reg646 <= ((({$signed(wire568)} ? (~&$unsigned(wire571)) : wire571) ?
                  {(-reg633[(3'h5):(3'h4)])} : (+($signed(wire572) ?
                      (~^reg631) : (wire569 ? reg644 : wire576)))) ?
              ($signed(({reg640, reg641} ?
                      $unsigned(wire636) : (wire637 || reg634))) ?
                  $unsigned(($unsigned(reg645) & $signed(reg633))) : (+((reg645 ?
                      wire630 : wire630) ~^ wire573[(4'h8):(2'h2)]))) : reg640);
        end
      else
        begin
          if ((reg646 <<< ((!(~|(8'hab))) ?
              (wire575 ?
                  (&((8'hb5) >> wire571)) : wire630[(1'h1):(1'h1)]) : $unsigned({((8'had) ~^ reg640),
                  (reg634 ? wire626 : wire570)}))))
            begin
              reg640 <= $signed(wire629[(3'h7):(2'h2)]);
              reg641 <= wire568;
              reg642 <= wire636;
              reg643 <= (wire568[(4'h9):(3'h7)] ?
                  $unsigned(($unsigned((~^wire568)) ?
                      (reg641 || (|wire626)) : ((reg646 != reg642) + $signed(wire626)))) : (~^(reg632[(4'hf):(4'hb)] ?
                      (wire630[(1'h0):(1'h0)] ?
                          $unsigned(reg643) : (-(8'hae))) : $signed((^~(8'h9d))))));
              reg644 <= (($unsigned((wire630 == $signed(reg639))) ?
                  ((wire574 ?
                          (reg634 ? (8'ha2) : wire636) : ((8'hb8) ^ wire638)) ?
                      ((reg639 ? (8'ha9) : reg640) ?
                          {reg645, wire576} : {wire629,
                              wire568}) : $signed((wire576 ?
                          reg646 : reg632))) : reg635) < reg632[(5'h11):(5'h11)]);
            end
          else
            begin
              reg640 <= (!($unsigned(reg641) ^ (~|wire626[(2'h2):(1'h0)])));
              reg641 <= wire569;
              reg642 <= {reg633};
            end
          reg645 <= ($signed($unsigned({(wire628 ? wire638 : wire575)})) ?
              reg645 : wire626[(4'h9):(4'h8)]);
          reg646 <= $unsigned(($signed(({wire572, reg644} ?
                  wire626[(3'h4):(1'h0)] : wire626)) ?
              $unsigned(wire638[(4'hc):(4'h8)]) : wire638));
        end
      reg647 <= {{reg633[(3'h4):(3'h4)],
              (((-wire630) << (~^wire571)) << {reg635[(2'h2):(2'h2)],
                  (wire576 + wire637)})},
          (reg641[(4'h9):(3'h7)] ?
              (reg640 & (~&(wire636 ? (8'haf) : wire571))) : wire570)};
      reg648 <= wire636[(4'ha):(1'h0)];
      reg649 <= $signed(wire638);
    end
  assign wire650 = $unsigned(($unsigned({(reg647 ^~ reg640)}) ?
                       {(reg640[(4'h8):(2'h2)] ?
                               wire568 : $signed(reg643))} : ((reg632[(4'he):(3'h5)] ?
                               reg640 : wire572[(1'h1):(1'h0)]) ?
                           (~&(wire637 >>> wire571)) : $signed($signed(reg633)))));
  assign wire651 = (~^{(~^(((8'hb2) & reg643) ?
                           $unsigned(wire568) : (~&wire626)))});
  module652 modinst668 (wire667, clk, wire570, wire630, wire568, wire575);
  assign wire669 = {$signed($unsigned($unsigned(reg640[(2'h3):(2'h2)]))),
                       {((8'hbe) == {wire629}), (8'hbd)}};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module652
#( parameter param665 = (((({(7'h43), (8'ha4)} >> (&(8'hac))) != ((8'hbc) ? {(8'hbf), (8'hb4)} : (8'hb7))) == (!(~&(-(8'hb7))))) ? ((~&(&((8'h9c) ? (7'h40) : (8'hbf)))) ^~ (^~((~|(7'h42)) << {(8'ha4)}))) : ((8'h9f) >= (!{((8'ha5) & (8'ha8))})))
, parameter param666 = {(((~&{param665, param665}) ? {(param665 | param665), (~^param665)} : (((8'ha3) ? param665 : param665) ? param665 : (param665 ^~ param665))) ? param665 : {(7'h44)}), (param665 || {((!param665) ? (param665 ? param665 : param665) : (param665 > param665)), (^(param665 | param665))})} )
(y, clk, wire656, wire655, wire654, wire653);
  output wire [(32'h6d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire656;
  input wire [(5'h10):(1'h0)] wire655;
  input wire [(3'h6):(1'h0)] wire654;
  input wire signed [(3'h7):(1'h0)] wire653;
  wire [(4'hf):(1'h0)] wire664;
  wire signed [(2'h3):(1'h0)] wire663;
  wire [(5'h15):(1'h0)] wire662;
  wire signed [(5'h11):(1'h0)] wire661;
  wire [(2'h2):(1'h0)] wire660;
  wire [(5'h15):(1'h0)] wire659;
  wire signed [(4'ha):(1'h0)] wire658;
  wire [(5'h13):(1'h0)] wire657;
  assign y = {wire664,
                 wire663,
                 wire662,
                 wire661,
                 wire660,
                 wire659,
                 wire658,
                 wire657,
                 (1'h0)};
  assign wire657 = $unsigned(($signed($signed($signed((8'hb5)))) ?
                       ((wire656 ?
                               {wire655, wire654} : wire653[(2'h3):(1'h0)]) ?
                           $unsigned($signed(wire654)) : (-wire653)) : wire656));
  assign wire658 = {wire656[(4'h9):(3'h7)]};
  assign wire659 = $signed($signed(($unsigned($unsigned(wire655)) ^ (wire655 ?
                       wire658 : $signed(wire657)))));
  assign wire660 = (8'hac);
  assign wire661 = $signed(((wire658[(3'h5):(3'h5)] == {wire657}) ?
                       $unsigned(wire659) : (wire660[(1'h0):(1'h0)] < wire654)));
  assign wire662 = ({wire661} << {(~|(wire658[(3'h5):(3'h4)] + ((8'hb4) ?
                           wire658 : (8'ha9))))});
  assign wire663 = ((~($unsigned({(8'h9f)}) >>> wire657[(3'h6):(2'h2)])) & wire655[(4'he):(4'ha)]);
  assign wire664 = (8'hba);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module577
#( parameter param625 = ((8'hbe) ? (({(+(8'hb4)), ((8'ha3) <<< (8'had))} ? (~&((7'h43) >> (8'ha2))) : ((~|(8'ha3)) ? ((8'h9e) || (7'h44)) : (~^(7'h44)))) ? (!(^~(8'hbf))) : ((((8'hab) ? (8'hb4) : (8'h9c)) ? ((8'hb0) <= (8'ha0)) : ((8'hba) ? (8'hb3) : (8'hab))) <= (((8'ha6) <<< (8'hac)) >= {(8'ha2)}))) : ({{((8'hb7) >> (8'ha1)), ((8'hb2) ~^ (8'ha6))}, (~^{(8'hb4), (8'h9e)})} * (~(8'hbc)))) )
(y, clk, wire582, wire581, wire580, wire579, wire578);
  output wire [(32'h20b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire582;
  input wire signed [(4'h9):(1'h0)] wire581;
  input wire signed [(5'h12):(1'h0)] wire580;
  input wire [(5'h15):(1'h0)] wire579;
  input wire signed [(3'h5):(1'h0)] wire578;
  wire signed [(4'hd):(1'h0)] wire624;
  wire [(4'hf):(1'h0)] wire623;
  reg signed [(4'hd):(1'h0)] reg622 = (1'h0);
  reg [(4'h9):(1'h0)] reg621 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg620 = (1'h0);
  wire [(5'h12):(1'h0)] wire619;
  wire signed [(4'hd):(1'h0)] wire618;
  reg signed [(5'h13):(1'h0)] reg617 = (1'h0);
  reg [(5'h12):(1'h0)] reg616 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire615;
  wire signed [(5'h11):(1'h0)] wire614;
  wire signed [(4'he):(1'h0)] wire613;
  reg signed [(3'h6):(1'h0)] reg612 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg611 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg610 = (1'h0);
  reg [(3'h5):(1'h0)] reg609 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg608 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg607 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg606 = (1'h0);
  reg signed [(4'he):(1'h0)] reg605 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg604 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg603 = (1'h0);
  reg [(4'h9):(1'h0)] reg602 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg601 = (1'h0);
  reg [(5'h14):(1'h0)] reg600 = (1'h0);
  reg [(4'hd):(1'h0)] reg599 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg598 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg597 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg596 = (1'h0);
  reg [(4'h8):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg594 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg593 = (1'h0);
  reg [(3'h7):(1'h0)] reg592 = (1'h0);
  reg signed [(4'he):(1'h0)] reg591 = (1'h0);
  reg signed [(4'he):(1'h0)] reg590 = (1'h0);
  reg [(4'h8):(1'h0)] reg589 = (1'h0);
  reg signed [(4'he):(1'h0)] reg588 = (1'h0);
  reg [(2'h3):(1'h0)] reg587 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire586;
  wire signed [(5'h11):(1'h0)] wire585;
  wire signed [(4'ha):(1'h0)] wire584;
  wire [(4'he):(1'h0)] wire583;
  assign y = {wire624,
                 wire623,
                 reg622,
                 reg621,
                 reg620,
                 wire619,
                 wire618,
                 reg617,
                 reg616,
                 wire615,
                 wire614,
                 wire613,
                 reg612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 wire586,
                 wire585,
                 wire584,
                 wire583,
                 (1'h0)};
  assign wire583 = $unsigned(wire582[(3'h4):(2'h2)]);
  assign wire584 = $unsigned($unsigned((~^wire582[(3'h4):(3'h4)])));
  assign wire585 = (wire582 | $unsigned((~&wire578[(2'h2):(2'h2)])));
  assign wire586 = $unsigned((wire580[(3'h7):(1'h1)] != $unsigned(wire585[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      if ((({(wire578[(2'h2):(1'h1)] ?
              wire583[(4'hd):(3'h5)] : wire583[(4'hd):(3'h4)]),
          wire584[(3'h4):(1'h0)]} > ($signed((~&wire584)) ?
          $unsigned((+wire585)) : (((8'ha3) != wire581) || (~^wire579)))) <= ($signed($unsigned((^wire584))) ?
          $unsigned(({wire585} ?
              $signed(wire579) : wire580[(4'hb):(3'h7)])) : $signed(($unsigned(wire585) != (-wire579))))))
        begin
          if ({wire584[(4'h8):(1'h0)]})
            begin
              reg587 <= {wire585};
              reg588 <= wire586;
              reg589 <= $signed(wire585);
            end
          else
            begin
              reg587 <= reg588[(1'h0):(1'h0)];
            end
          reg590 <= $signed({$signed((((7'h41) - reg588) ?
                  (wire585 ? wire584 : wire582) : (wire580 == wire579)))});
          if (wire581[(1'h1):(1'h1)])
            begin
              reg591 <= $signed($unsigned(((wire584[(2'h3):(2'h3)] >= (reg587 > wire581)) | wire586)));
              reg592 <= ($unsigned((wire585[(4'h8):(2'h2)] ~^ reg591)) ^~ $signed(reg591));
              reg593 <= (wire586[(3'h5):(3'h4)] ?
                  $unsigned((reg592[(3'h6):(3'h5)] ?
                      (reg588[(2'h3):(1'h0)] ?
                          {(8'hb7),
                              wire580} : $signed(wire580)) : $unsigned((^reg592)))) : (~|(((~&(8'had)) ^ (wire585 ?
                      (8'hb3) : (8'hab))) <<< wire582[(3'h4):(2'h2)])));
            end
          else
            begin
              reg591 <= $unsigned(($unsigned(({reg591} ?
                  $signed(reg592) : $unsigned(wire584))) << ((^~$unsigned(wire583)) ^ ($unsigned(wire581) > reg593))));
              reg592 <= ((7'h40) <= {wire585,
                  (wire579[(3'h6):(2'h3)] <<< wire581)});
            end
          if (wire583[(3'h4):(2'h3)])
            begin
              reg594 <= reg588;
              reg595 <= (($signed((8'haf)) ?
                      (~^$signed((reg588 + wire579))) : (((wire586 ?
                          wire583 : wire584) ^ $signed((8'hbe))) - (~|$signed((8'h9d))))) ?
                  (~$unsigned($unsigned(wire583[(4'hc):(4'h8)]))) : reg594[(4'ha):(3'h6)]);
              reg596 <= reg587;
            end
          else
            begin
              reg594 <= {reg595[(1'h1):(1'h1)],
                  $unsigned($unsigned({(reg595 && reg593)}))};
              reg595 <= ($unsigned(((+(^reg587)) ~^ reg591)) ?
                  wire578 : reg587[(2'h3):(1'h0)]);
            end
          reg597 <= (~($unsigned(({reg592} ?
                  $unsigned(wire584) : $signed((8'hb5)))) ?
              wire583[(1'h0):(1'h0)] : ($signed(((8'hb8) ? wire582 : wire578)) ?
                  $unsigned($unsigned(wire579)) : {$unsigned(wire581)})));
        end
      else
        begin
          reg587 <= $unsigned((~^reg590));
          reg588 <= $unsigned((wire581[(2'h2):(1'h0)] ?
              (8'hba) : $unsigned($signed((wire580 ? reg592 : (8'hb7))))));
          reg589 <= $signed(((wire585 ?
                  wire578[(1'h0):(1'h0)] : $signed((+wire585))) ?
              (+(^(reg588 != wire580))) : (8'haa)));
          reg590 <= reg589;
        end
      if ({{wire585[(3'h6):(3'h4)]}})
        begin
          reg598 <= (|{(8'h9f), wire579[(4'ha):(2'h2)]});
          reg599 <= wire585;
        end
      else
        begin
          if (($unsigned(($signed(reg599[(1'h0):(1'h0)]) ?
                  wire585 : reg597[(4'h9):(4'h8)])) ?
              (^wire578) : $unsigned($unsigned(reg595))))
            begin
              reg598 <= (reg598[(1'h1):(1'h1)] != ((&$signed(wire585)) <<< wire582[(1'h1):(1'h1)]));
              reg599 <= $unsigned($signed((reg590[(4'hd):(3'h6)] >> (wire582[(2'h3):(1'h0)] ?
                  reg595 : {wire579}))));
            end
          else
            begin
              reg598 <= (reg587 ?
                  reg599 : $signed(($signed($unsigned(reg597)) + (~|(-wire581)))));
              reg599 <= $signed($signed((~&wire586)));
              reg600 <= $signed((|reg595));
              reg601 <= $signed({(^(~reg593[(2'h2):(1'h1)])), $signed(reg600)});
            end
          reg602 <= ((8'hb6) - (reg599 >>> {$unsigned(reg592[(2'h2):(1'h0)]),
              $signed((wire580 ? reg592 : wire581))}));
          if ((8'hb4))
            begin
              reg603 <= (^reg589[(3'h5):(1'h1)]);
              reg604 <= reg594;
            end
          else
            begin
              reg603 <= $signed(reg594[(2'h2):(1'h1)]);
              reg604 <= $unsigned({$unsigned(($signed(reg600) & (wire580 * reg598))),
                  (($unsigned(wire584) ?
                          {reg589} : (reg600 ? reg603 : (8'h9e))) ?
                      (8'ha9) : ((reg597 ? wire586 : wire580) ?
                          (+wire581) : $unsigned(reg587)))});
              reg605 <= ((8'h9e) <= (~{wire581}));
            end
          reg606 <= {(&reg587), reg599};
          reg607 <= (&$signed((^~$signed(wire583[(3'h5):(3'h5)]))));
        end
    end
  always
    @(posedge clk) begin
      reg608 <= ($unsigned(((~&(reg595 ?
          wire582 : reg605)) ~^ reg605)) - {(~$signed((wire579 | (8'hbf)))),
          reg590});
      reg609 <= (~|((reg598 ?
              reg599[(1'h0):(1'h0)] : {(&reg596), $signed(wire585)}) ?
          (($unsigned(reg602) & reg600) && wire581) : (reg587 ?
              ((~reg600) + (reg600 != reg595)) : reg598[(1'h0):(1'h0)])));
      reg610 <= $unsigned(reg599);
      reg611 <= $signed($unsigned(($unsigned(reg598) - ({wire582, reg589} ?
          $signed(reg594) : wire582[(2'h3):(1'h0)]))));
      reg612 <= wire586[(4'h9):(3'h6)];
    end
  assign wire613 = ($unsigned($signed($signed($unsigned(wire585)))) + (($unsigned($unsigned(wire583)) * $signed(reg597[(3'h6):(1'h1)])) ?
                       $unsigned(wire582) : $signed({(reg609 + reg609),
                           $signed((8'hb3))})));
  assign wire614 = (($unsigned((8'ha9)) ?
                           wire583[(3'h4):(3'h4)] : wire581[(4'h9):(1'h0)]) ?
                       wire583[(4'ha):(2'h3)] : ($signed((^~(!wire580))) >= (~^(reg611[(2'h2):(2'h2)] && $signed(wire613)))));
  assign wire615 = (!{wire614});
  always
    @(posedge clk) begin
      if (({$signed((wire578[(2'h2):(1'h1)] << reg596[(1'h0):(1'h0)])),
          reg599[(3'h7):(3'h4)]} < $unsigned($signed(($signed(wire615) ?
          (wire584 ? reg587 : reg588) : (-reg598))))))
        begin
          reg616 <= reg601;
          reg617 <= $unsigned(wire614[(3'h7):(3'h4)]);
        end
      else
        begin
          reg616 <= (8'hb5);
          reg617 <= (8'ha8);
        end
    end
  assign wire618 = reg601;
  assign wire619 = reg605[(3'h5):(1'h1)];
  always
    @(posedge clk) begin
      reg620 <= (8'hb9);
      reg621 <= (reg610[(3'h6):(1'h1)] ?
          ($signed($unsigned(((8'haf) & wire579))) > {(reg591[(2'h2):(1'h0)] >= (7'h42)),
              ($unsigned(reg595) ^ $unsigned(reg606))}) : (~&(wire583[(4'ha):(1'h1)] == ({reg602,
                  reg600} ?
              {wire614, wire585} : {reg594, reg610}))));
      reg622 <= wire615;
    end
  assign wire623 = ({{(8'ha0)},
                           (^((reg591 ?
                               reg595 : reg620) * ((8'ha8) - wire580)))} ?
                       $unsigned((wire581[(3'h6):(3'h5)] <= $signed((8'hb6)))) : $signed((8'had)));
  assign wire624 = $unsigned((~^reg593));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module683  (y, clk, wire687, wire686, wire685, wire684);
  output wire [(32'h1b0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire687;
  input wire [(2'h2):(1'h0)] wire686;
  input wire signed [(4'h9):(1'h0)] wire685;
  input wire [(5'h10):(1'h0)] wire684;
  wire signed [(3'h7):(1'h0)] wire721;
  wire [(4'hc):(1'h0)] wire720;
  wire [(4'he):(1'h0)] wire719;
  reg [(3'h7):(1'h0)] reg718 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg717 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg716 = (1'h0);
  reg [(3'h5):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg714 = (1'h0);
  reg [(3'h7):(1'h0)] reg713 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg712 = (1'h0);
  reg [(4'h9):(1'h0)] reg711 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire710;
  wire [(3'h5):(1'h0)] wire709;
  wire [(4'he):(1'h0)] wire708;
  reg [(4'h8):(1'h0)] reg707 = (1'h0);
  reg [(5'h10):(1'h0)] reg706 = (1'h0);
  reg [(5'h12):(1'h0)] reg705 = (1'h0);
  reg [(2'h2):(1'h0)] reg704 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg703 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg702 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg701 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg700 = (1'h0);
  reg [(5'h13):(1'h0)] reg699 = (1'h0);
  reg [(4'h9):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg697 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg696 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg695 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg694 = (1'h0);
  reg [(4'hd):(1'h0)] reg693 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg692 = (1'h0);
  reg [(4'h8):(1'h0)] reg691 = (1'h0);
  reg [(5'h15):(1'h0)] reg690 = (1'h0);
  reg [(4'ha):(1'h0)] reg689 = (1'h0);
  wire [(5'h10):(1'h0)] wire688;
  assign y = {wire721,
                 wire720,
                 wire719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 reg713,
                 reg712,
                 reg711,
                 wire710,
                 wire709,
                 wire708,
                 reg707,
                 reg706,
                 reg705,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 reg699,
                 reg698,
                 reg697,
                 reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 reg691,
                 reg690,
                 reg689,
                 wire688,
                 (1'h0)};
  assign wire688 = ({$signed((wire685 ?
                           ((8'ha2) | wire687) : $signed((8'hbd)))),
                       ($signed((wire687 <= wire684)) ?
                           wire687 : (+(-wire687)))} != (!(^~{$signed(wire685)})));
  always
    @(posedge clk) begin
      if ({$signed((wire684 & (8'hab))),
          ((|wire688[(4'hc):(3'h4)]) ? wire688 : {wire686})})
        begin
          reg689 <= $signed(wire688[(3'h6):(3'h4)]);
          reg690 <= {$signed(wire684[(4'hf):(4'ha)]), wire686};
          reg691 <= wire688;
          reg692 <= $signed((~{reg689[(4'h9):(1'h1)], wire687[(2'h2):(2'h2)]}));
        end
      else
        begin
          if (wire688[(4'he):(2'h3)])
            begin
              reg689 <= $signed($unsigned(reg692));
              reg690 <= ($signed(wire687[(3'h4):(2'h3)]) > $unsigned($unsigned(((~^(8'hae)) ?
                  {wire686} : (wire685 <<< wire684)))));
              reg691 <= (($unsigned(((reg689 >>> reg691) ?
                      {reg691,
                          wire687} : (wire687 < reg691))) >= wire685[(3'h4):(3'h4)]) ?
                  wire686[(1'h1):(1'h1)] : reg690[(5'h14):(3'h6)]);
            end
          else
            begin
              reg689 <= $signed($unsigned((|{(wire684 ? wire687 : wire684),
                  (&(7'h40))})));
              reg690 <= wire688;
              reg691 <= $signed(($signed((reg692 & $unsigned(reg690))) ?
                  (wire684 ?
                      (((8'hb8) ? reg690 : (8'hb1)) | (reg691 ?
                          wire686 : (8'ha7))) : ((|wire686) ?
                          $unsigned(reg692) : $unsigned(reg691))) : $signed((wire684[(3'h6):(3'h5)] & (!reg689)))));
              reg692 <= (^~reg691);
            end
          if (reg691[(3'h7):(2'h3)])
            begin
              reg693 <= reg689;
              reg694 <= ((|$signed(reg689[(1'h0):(1'h0)])) ?
                  $unsigned((reg691[(4'h8):(3'h4)] ?
                      ((|wire687) ~^ (!reg692)) : $unsigned((~|wire686)))) : $unsigned(reg691[(3'h4):(1'h1)]));
              reg695 <= {$signed(reg689),
                  (&((~^(reg694 ?
                      reg691 : wire686)) << $signed($signed(wire686))))};
            end
          else
            begin
              reg693 <= wire685[(3'h7):(2'h2)];
              reg694 <= (8'hb4);
              reg695 <= (|(!reg690[(3'h5):(1'h1)]));
              reg696 <= $unsigned((~|$signed((-$unsigned(wire685)))));
              reg697 <= wire686;
            end
          if (wire684)
            begin
              reg698 <= (~^wire687);
              reg699 <= $signed((wire685[(3'h5):(2'h3)] <= (((wire684 ?
                          reg690 : (8'hb4)) ?
                      reg698 : (reg696 ? reg691 : reg693)) ?
                  $unsigned((^reg691)) : wire686)));
            end
          else
            begin
              reg698 <= (reg690[(4'hf):(4'hb)] ?
                  $signed(($unsigned((~^reg694)) ? reg694 : reg690)) : reg696);
              reg699 <= $unsigned((($unsigned($unsigned((8'hbb))) & ((reg698 > reg690) || $unsigned(reg695))) ?
                  reg690 : (~|wire686)));
            end
        end
      reg700 <= reg692[(3'h6):(2'h2)];
      if (((~&reg692) ?
          ($signed(((wire686 >> (8'hb0)) <= reg694[(4'h8):(2'h2)])) ?
              ((~&(reg697 > (8'hb6))) ?
                  $signed(reg698) : wire685[(3'h7):(1'h1)]) : ($unsigned($signed((8'h9e))) ?
                  (&(^~reg698)) : (!reg700))) : (!reg700[(3'h4):(2'h2)])))
        begin
          if (reg689[(4'h9):(3'h4)])
            begin
              reg701 <= (~(((8'ha9) != ((8'ha1) ?
                  (wire688 ?
                      reg700 : reg695) : $unsigned(wire684))) * (((reg697 ?
                      reg692 : reg699) ?
                  wire684 : (+reg692)) & $signed($unsigned(reg689)))));
              reg702 <= {(~|(^$signed((reg692 != reg698))))};
            end
          else
            begin
              reg701 <= (8'hab);
              reg702 <= (reg694[(4'ha):(3'h4)] ?
                  reg694 : (~^$signed($signed($unsigned(reg698)))));
              reg703 <= {(reg702[(4'ha):(4'h9)] ?
                      ((~reg697) ?
                          (wire684[(2'h3):(1'h0)] ?
                              {reg700} : $signed(reg701)) : $signed($unsigned(wire688))) : (7'h44))};
              reg704 <= $unsigned(reg699[(5'h10):(1'h0)]);
              reg705 <= $unsigned($unsigned(reg703[(4'hb):(2'h2)]));
            end
        end
      else
        begin
          if ($signed($unsigned(reg698)))
            begin
              reg701 <= wire686;
            end
          else
            begin
              reg701 <= reg705;
            end
          reg702 <= $unsigned(($signed((8'ha9)) ?
              $unsigned($signed(reg703)) : reg697));
          if ((!reg695[(4'ha):(3'h5)]))
            begin
              reg703 <= $unsigned($signed((-reg691)));
              reg704 <= $signed({$unsigned(reg692[(4'hd):(3'h4)])});
              reg705 <= reg692;
              reg706 <= wire686[(2'h2):(2'h2)];
            end
          else
            begin
              reg703 <= $unsigned($unsigned($unsigned($signed($signed(reg701)))));
              reg704 <= reg703;
              reg705 <= (~|$signed($unsigned($signed($signed(reg695)))));
              reg706 <= ($signed(($signed(wire686[(2'h2):(1'h0)]) ?
                      $signed($signed(reg700)) : ((reg701 <<< reg690) >= ((8'hb1) ?
                          reg698 : reg698)))) ?
                  wire687[(3'h4):(3'h4)] : reg702);
              reg707 <= (((reg690[(5'h14):(5'h14)] ?
                      ($signed(reg699) ?
                          (^~reg696) : $signed(reg703)) : wire687) >> wire687[(3'h5):(3'h4)]) ?
                  ((($unsigned(reg691) ?
                              reg697 : (wire686 ? wire688 : (8'hb2))) ?
                          reg695[(3'h5):(1'h1)] : reg693) ?
                      $signed(wire687) : $unsigned($unsigned((reg689 ?
                          reg703 : reg694)))) : ({(wire686[(1'h1):(1'h1)] ~^ reg695[(3'h6):(1'h0)])} ?
                      (reg705 ?
                          (reg689[(3'h5):(3'h5)] ?
                              ((8'hb9) ?
                                  (8'hb4) : (8'hb6)) : reg691[(3'h6):(1'h1)]) : reg694) : wire684[(4'ha):(3'h7)]));
            end
        end
    end
  assign wire708 = {($signed(({(8'hb2), reg693} ?
                               (!reg693) : $unsigned(wire686))) ?
                           ((~^(reg693 ? wire686 : reg702)) ?
                               (7'h44) : (~^$unsigned(reg696))) : {$signed(wire686)}),
                       (wire685 || wire685[(3'h4):(1'h1)])};
  assign wire709 = (reg695[(4'hb):(4'hb)] || reg700[(5'h14):(1'h1)]);
  assign wire710 = (((({(7'h41)} - $signed(wire686)) <<< (&(reg704 ?
                       reg704 : reg702))) * (-$signed(reg696[(4'he):(4'h9)]))) & reg699);
  always
    @(posedge clk) begin
      if ((((reg691[(2'h3):(2'h2)] != $signed((reg701 ? wire685 : reg694))) ?
          $signed($unsigned((reg704 > (8'hb5)))) : (~|reg705[(4'h9):(2'h3)])) <= $signed((-({reg694} > reg691)))))
        begin
          reg711 <= reg692[(3'h7):(3'h4)];
        end
      else
        begin
          reg711 <= ((~$unsigned($signed(reg698))) ?
              $signed(($unsigned((8'haa)) <<< reg705[(4'h8):(3'h5)])) : (($signed(wire710[(3'h4):(1'h0)]) >= $signed(((8'h9e) ?
                      reg689 : wire709))) ?
                  $unsigned($signed((reg690 << (7'h41)))) : reg694));
        end
      if ((~&reg699))
        begin
          reg712 <= reg702[(2'h2):(1'h1)];
          if (reg690)
            begin
              reg713 <= $unsigned(reg700);
              reg714 <= ($unsigned({(8'hbd)}) ?
                  wire684[(2'h3):(2'h3)] : ((((~^reg705) ?
                          (!reg697) : (reg691 ?
                              (8'had) : reg698)) > (reg691[(2'h3):(2'h3)] || reg702[(5'h12):(4'h9)])) ?
                      $signed((reg690[(4'h9):(3'h7)] <= (reg704 ?
                          wire688 : reg711))) : ((reg707[(3'h4):(2'h3)] && ((8'hbe) * wire685)) <= $unsigned(reg693))));
              reg715 <= ({(8'hb0),
                  ((~$signed(wire686)) ?
                      ($signed((8'hac)) - (reg694 << (8'had))) : wire685)} << reg702[(5'h10):(4'h8)]);
              reg716 <= reg689[(3'h5):(3'h5)];
              reg717 <= $unsigned(reg702);
            end
          else
            begin
              reg713 <= $signed({($signed($unsigned(reg701)) ?
                      ((reg703 ?
                          reg712 : reg702) <= (wire686 | reg699)) : (reg697[(3'h6):(2'h3)] | {wire709}))});
              reg714 <= (((wire709 ?
                      reg716[(2'h2):(1'h1)] : $signed({wire685})) ?
                  (8'ha0) : wire686[(2'h2):(1'h0)]) >>> wire710[(1'h1):(1'h1)]);
              reg715 <= (+((|reg698[(3'h6):(3'h4)]) ?
                  (($signed(reg715) & $unsigned((8'ha4))) > ({wire709} ?
                      $unsigned(wire688) : reg707)) : {$signed($signed(reg711)),
                      ((reg712 ? (8'haa) : reg700) << $signed((8'hb1)))}));
            end
        end
      else
        begin
          if ((&reg699[(4'hc):(4'ha)]))
            begin
              reg712 <= ((~^reg706) >= ((^~{reg691}) << (reg697[(4'hf):(4'h9)] >>> $unsigned($signed(wire709)))));
            end
          else
            begin
              reg712 <= (reg706 ^ reg716);
              reg713 <= reg715[(1'h0):(1'h0)];
              reg714 <= ((~&$unsigned((8'h9e))) <= reg714);
              reg715 <= reg714[(4'ha):(4'ha)];
            end
        end
      reg718 <= (~^reg712);
    end
  assign wire719 = (wire685[(2'h3):(2'h2)] << {$signed($unsigned($signed(reg698))),
                       {reg696}});
  assign wire720 = reg707;
  assign wire721 = (8'ha0);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module792
#( parameter param852 = {((((~^(8'hae)) >= (^(8'haf))) <= {((8'hae) ? (8'ha5) : (8'ha5)), (!(7'h43))}) ? (!(|((8'ha3) || (8'hb8)))) : (~{(8'haf), (!(8'h9f))}))}
, parameter param853 = (&{(^param852), param852}) )
(y, clk, wire796, wire795, wire794, wire793);
  output wire [(32'h24f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire796;
  input wire signed [(5'h11):(1'h0)] wire795;
  input wire [(3'h7):(1'h0)] wire794;
  input wire signed [(5'h15):(1'h0)] wire793;
  reg [(2'h2):(1'h0)] reg851 = (1'h0);
  reg [(4'h9):(1'h0)] reg850 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg849 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg848 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg847 = (1'h0);
  wire [(4'h8):(1'h0)] wire846;
  wire signed [(4'h8):(1'h0)] wire845;
  wire signed [(5'h10):(1'h0)] wire844;
  wire signed [(4'h9):(1'h0)] wire843;
  wire [(4'he):(1'h0)] wire842;
  wire signed [(3'h6):(1'h0)] wire841;
  reg [(5'h15):(1'h0)] reg840 = (1'h0);
  reg [(5'h14):(1'h0)] reg839 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg838 = (1'h0);
  reg [(5'h10):(1'h0)] reg837 = (1'h0);
  reg [(4'ha):(1'h0)] reg836 = (1'h0);
  wire [(3'h4):(1'h0)] wire835;
  reg signed [(5'h12):(1'h0)] reg834 = (1'h0);
  reg [(3'h6):(1'h0)] reg833 = (1'h0);
  reg [(4'hb):(1'h0)] reg832 = (1'h0);
  reg [(4'hf):(1'h0)] reg831 = (1'h0);
  reg [(2'h2):(1'h0)] reg830 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg829 = (1'h0);
  reg [(2'h2):(1'h0)] reg828 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg827 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg826 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg825 = (1'h0);
  reg [(2'h3):(1'h0)] reg824 = (1'h0);
  reg [(4'hb):(1'h0)] reg823 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg822 = (1'h0);
  reg [(4'hf):(1'h0)] reg821 = (1'h0);
  reg [(2'h3):(1'h0)] reg820 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg819 = (1'h0);
  wire [(3'h4):(1'h0)] wire818;
  wire signed [(5'h14):(1'h0)] wire817;
  wire signed [(3'h7):(1'h0)] wire816;
  wire signed [(3'h6):(1'h0)] wire815;
  wire [(4'he):(1'h0)] wire814;
  wire signed [(5'h14):(1'h0)] wire813;
  wire signed [(3'h7):(1'h0)] wire812;
  reg signed [(4'hb):(1'h0)] reg811 = (1'h0);
  reg [(5'h11):(1'h0)] reg810 = (1'h0);
  reg [(4'he):(1'h0)] reg809 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg808 = (1'h0);
  reg [(5'h13):(1'h0)] reg807 = (1'h0);
  reg [(5'h15):(1'h0)] reg806 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg805 = (1'h0);
  reg [(5'h15):(1'h0)] reg804 = (1'h0);
  reg [(2'h2):(1'h0)] reg803 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg802 = (1'h0);
  reg [(5'h11):(1'h0)] reg801 = (1'h0);
  reg [(2'h2):(1'h0)] reg800 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire799;
  wire [(3'h4):(1'h0)] wire798;
  wire signed [(3'h4):(1'h0)] wire797;
  assign y = {reg851,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 wire846,
                 wire845,
                 wire844,
                 wire843,
                 wire842,
                 wire841,
                 reg840,
                 reg839,
                 reg838,
                 reg837,
                 reg836,
                 wire835,
                 reg834,
                 reg833,
                 reg832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 reg827,
                 reg826,
                 reg825,
                 reg824,
                 reg823,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 wire818,
                 wire817,
                 wire816,
                 wire815,
                 wire814,
                 wire813,
                 wire812,
                 reg811,
                 reg810,
                 reg809,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg802,
                 reg801,
                 reg800,
                 wire799,
                 wire798,
                 wire797,
                 (1'h0)};
  assign wire797 = wire795[(3'h7):(1'h0)];
  assign wire798 = wire796;
  assign wire799 = wire793;
  always
    @(posedge clk) begin
      if ($unsigned($signed((({wire793} ?
              wire795[(4'hf):(3'h4)] : wire799[(3'h5):(2'h2)]) ?
          (((8'ha9) != wire798) >>> ((8'hb9) >= wire795)) : ((wire797 ?
                  wire797 : wire797) ?
              (^~wire796) : wire794)))))
        begin
          reg800 <= wire795;
          reg801 <= ((wire798 ? wire798[(2'h2):(2'h2)] : wire797) ?
              (~^(~|$unsigned((wire794 ?
                  wire799 : wire796)))) : $signed($unsigned((8'haf))));
          if ($unsigned((wire796 ?
              (wire798 ^~ wire798) : $unsigned(wire797[(3'h4):(1'h1)]))))
            begin
              reg802 <= {reg800[(2'h2):(1'h0)]};
              reg803 <= $signed({wire796[(5'h10):(4'hf)]});
              reg804 <= $signed(((((8'h9e) ?
                      reg801[(4'he):(1'h0)] : wire798) + (|{wire797})) ?
                  wire797[(2'h3):(1'h0)] : wire795));
              reg805 <= wire794[(3'h7):(3'h7)];
            end
          else
            begin
              reg802 <= (((wire799[(2'h2):(2'h2)] != (&reg804[(5'h12):(3'h7)])) < ({$signed((8'ha1)),
                  {wire794,
                      reg801}} < reg800[(1'h0):(1'h0)])) || $signed((|reg802)));
              reg803 <= ($signed((~|$unsigned((wire797 | reg803)))) & $unsigned($signed((|$signed(reg803)))));
            end
          reg806 <= $unsigned($unsigned({($unsigned(reg804) ?
                  $signed(wire799) : (reg805 ? wire793 : wire797))}));
          reg807 <= wire793[(5'h10):(1'h1)];
        end
      else
        begin
          if ((reg805 || reg802))
            begin
              reg800 <= (+(reg800[(2'h2):(1'h1)] >= $unsigned(wire796[(5'h10):(3'h6)])));
              reg801 <= $signed($unsigned((wire799 != $unsigned((reg800 | wire793)))));
              reg802 <= (((wire794 ?
                          ({(8'ha6), wire796} ?
                              $unsigned(wire797) : $unsigned((8'hb9))) : wire799) ?
                      $unsigned((8'hba)) : reg807[(4'he):(4'he)]) ?
                  wire797[(2'h3):(2'h3)] : ($unsigned($signed((^~reg802))) ^ {wire794}));
              reg803 <= $unsigned((|(+wire794)));
            end
          else
            begin
              reg800 <= {$unsigned(wire799)};
              reg801 <= wire796;
              reg802 <= (reg803 ^~ reg803);
              reg803 <= ((|$signed(wire796[(3'h7):(2'h2)])) ^~ (($signed($unsigned(wire793)) ?
                      ($signed(wire794) ?
                          reg807 : ((8'hbe) != wire794)) : wire796) ?
                  wire797[(1'h0):(1'h0)] : (+(reg802[(3'h7):(2'h2)] >> $unsigned(reg801)))));
              reg804 <= (|$unsigned($signed((wire797[(1'h1):(1'h0)] != (reg804 ?
                  wire798 : reg802)))));
            end
          if (reg807)
            begin
              reg805 <= reg801;
              reg806 <= (7'h43);
            end
          else
            begin
              reg805 <= {($signed(((&(7'h42)) ?
                      (reg804 ?
                          reg802 : reg805) : ((8'ha5) > (8'ha2)))) < (wire793[(2'h2):(1'h0)] | $signed((wire795 & (8'ha1))))),
                  (^(({reg804} ? $signed(reg803) : $signed(reg801)) - reg805))};
            end
          reg807 <= (|(!reg801));
          reg808 <= (reg805 ?
              ($unsigned({$signed(wire798)}) + $signed(((wire799 ?
                      wire795 : wire795) ?
                  wire797 : (reg806 ?
                      reg801 : reg806)))) : $signed($signed(((~^(7'h42)) | (reg806 >>> reg800)))));
        end
      reg809 <= reg807[(3'h7):(3'h6)];
      reg810 <= $unsigned(wire797);
      reg811 <= ((($unsigned((~^(8'hab))) >= $unsigned((8'hab))) >>> (wire798[(2'h3):(1'h0)] ?
          reg806[(4'hd):(2'h2)] : (wire796[(1'h0):(1'h0)] ?
              reg801[(2'h2):(2'h2)] : $signed(wire795)))) * wire796);
    end
  assign wire812 = reg802;
  assign wire813 = wire797[(1'h0):(1'h0)];
  assign wire814 = {(^~wire795[(2'h3):(1'h0)])};
  assign wire815 = ($unsigned(wire813[(2'h2):(1'h1)]) || reg803[(1'h1):(1'h0)]);
  assign wire816 = $signed(((reg800 ? wire793 : $unsigned((+(8'ha0)))) ?
                       $signed($signed({wire799})) : ($signed(wire812[(1'h1):(1'h0)]) != (wire813[(4'ha):(3'h5)] * reg801[(3'h5):(2'h2)]))));
  assign wire817 = ((-wire796) ?
                       $unsigned((~&(~|wire793))) : (^~(wire796 ?
                           (+{wire814}) : (^reg804))));
  assign wire818 = $unsigned($signed($unsigned(reg807)));
  always
    @(posedge clk) begin
      reg819 <= (~|$signed($signed(reg807)));
      if (wire818)
        begin
          if ($signed((wire798 ?
              (((^~(7'h42)) ?
                  (wire817 || wire813) : (reg804 ?
                      reg803 : (8'ha5))) >= (~|$unsigned(reg805))) : {($signed(reg806) & (|reg805))})))
            begin
              reg820 <= wire795[(3'h7):(1'h1)];
              reg821 <= (+$signed((~$unsigned(reg802[(4'he):(2'h2)]))));
              reg822 <= $signed((-$unsigned(((wire814 ? wire793 : (8'ha4)) ?
                  $unsigned(reg821) : (wire799 ? wire817 : reg805)))));
            end
          else
            begin
              reg820 <= wire814;
              reg821 <= $signed(reg806);
              reg822 <= wire798[(2'h2):(1'h1)];
              reg823 <= ($signed((!{((8'haf) ?
                      wire815 : reg807)})) - $signed(reg802[(4'ha):(4'h9)]));
              reg824 <= ($unsigned(reg800[(1'h1):(1'h0)]) <<< $unsigned($unsigned((^reg802))));
            end
          if ((|(+$signed({(~^wire817), wire816}))))
            begin
              reg825 <= (((wire797 >> reg805[(3'h6):(1'h0)]) ?
                      $unsigned(($unsigned(wire799) == wire816[(3'h5):(1'h1)])) : {((wire813 ^~ wire797) <<< $signed(wire812))}) ?
                  wire796 : $signed({$signed((reg806 ? wire816 : wire818))}));
              reg826 <= (($unsigned($unsigned((reg811 ?
                      wire799 : wire814))) ^ $unsigned(reg824)) ?
                  (&(reg802[(3'h5):(2'h3)] ~^ $signed($unsigned(reg806)))) : (wire814[(4'h8):(2'h3)] ?
                      (|$signed($signed(reg824))) : $unsigned($unsigned((reg811 || wire794)))));
              reg827 <= reg804[(1'h0):(1'h0)];
            end
          else
            begin
              reg825 <= $signed($signed((((~|reg806) < reg807) < reg808)));
              reg826 <= $signed(wire812);
              reg827 <= (&(wire793 - reg801));
              reg828 <= {wire815[(3'h4):(2'h2)]};
            end
          if (((|($unsigned((reg826 ?
                  reg828 : reg822)) && $signed($signed(reg804)))) ?
              (|($signed((wire816 < (8'hbf))) ?
                  wire812[(1'h0):(1'h0)] : reg807)) : $signed(reg819)))
            begin
              reg829 <= (&reg822[(2'h3):(1'h0)]);
            end
          else
            begin
              reg829 <= (reg826 ? $signed((8'h9d)) : wire817);
              reg830 <= ((((8'hac) ^ $signed({wire814,
                  wire818})) > (reg826[(1'h1):(1'h1)] > $signed(((8'ha7) >= reg819)))) >>> $signed((~|($signed(wire797) || $signed((8'hbd))))));
            end
          reg831 <= (reg825 <= ($signed(reg820) ?
              $signed($signed((wire816 <= wire793))) : (!wire794)));
          reg832 <= (($unsigned($signed(reg808[(2'h2):(2'h2)])) ?
              $unsigned($unsigned((|reg822))) : ($unsigned($unsigned(wire818)) >>> ({reg801,
                      reg811} ?
                  {reg823} : reg801))) << (^~((+(8'hbe)) ?
              (~^(^reg803)) : ($unsigned((8'ha4)) ^ wire815))));
        end
      else
        begin
          reg820 <= ($signed((((8'hb0) + $signed(wire797)) > ((reg804 != reg801) && wire816))) ?
              $signed((~|{reg811,
                  {reg821}})) : ({$signed(wire799[(3'h5):(1'h1)])} <<< ($unsigned({wire815,
                      reg810}) ?
                  reg805 : ($unsigned(reg801) * reg819[(4'he):(4'hd)]))));
        end
      reg833 <= (~(^~(&$signed($unsigned(reg831)))));
      reg834 <= $unsigned(($unsigned(((reg831 ? wire817 : (8'hbb)) ?
              $signed(wire815) : (^reg820))) ?
          (-$signed((8'hb0))) : (&$signed((!wire816)))));
    end
  assign wire835 = wire795[(4'hb):(2'h2)];
  always
    @(posedge clk) begin
      reg836 <= $unsigned(reg801);
      reg837 <= (8'h9d);
      reg838 <= {($unsigned((!reg833[(2'h2):(1'h1)])) ?
              $unsigned($signed((-wire795))) : ((reg807 ?
                      wire793 : reg810[(4'hc):(1'h1)]) ?
                  (~&reg824[(2'h2):(1'h0)]) : ({reg801,
                      wire814} >= $unsigned((8'hb1)))))};
      reg839 <= reg824[(1'h0):(1'h0)];
      reg840 <= reg821;
    end
  assign wire841 = wire793;
  assign wire842 = (((reg808 ?
                           $unsigned(wire814) : ((reg830 ? reg827 : wire812) ?
                               reg830[(2'h2):(1'h1)] : wire798[(2'h3):(1'h0)])) >= $unsigned(((reg822 ?
                               reg819 : reg834) ?
                           ((8'hba) && wire796) : $unsigned((8'hbe))))) ?
                       $unsigned($unsigned($signed(wire794))) : (^~(+reg820[(2'h2):(1'h0)])));
  assign wire843 = reg824[(1'h1):(1'h0)];
  assign wire844 = reg806[(1'h0):(1'h0)];
  assign wire845 = wire842;
  assign wire846 = $unsigned($unsigned(wire798));
  always
    @(posedge clk) begin
      reg847 <= (~^(~|reg820));
      reg848 <= (^{$signed(({wire797, wire841} ? {reg840} : reg810))});
    end
  always
    @(posedge clk) begin
      reg849 <= (reg839[(4'h8):(3'h7)] == ((((+(8'had)) < wire843[(1'h1):(1'h1)]) ?
              reg834 : (reg848 || $unsigned(wire841))) ?
          $signed($signed(reg848)) : wire798[(2'h2):(1'h1)]));
      reg850 <= $unsigned($signed($signed($signed($signed((8'h9f))))));
      reg851 <= (($signed(reg825[(1'h1):(1'h0)]) ?
              (~|((wire794 ? reg806 : reg839) >>> reg807)) : reg839) ?
          reg829 : ((wire797 ?
                  $unsigned(reg820[(1'h1):(1'h1)]) : (((8'ha7) <= reg848) != wire817)) ?
              (reg805[(4'h8):(3'h7)] ?
                  ($unsigned(reg807) >> (~|reg806)) : reg820[(1'h0):(1'h0)]) : ($unsigned($signed(wire798)) ?
                  wire799[(3'h7):(3'h5)] : $unsigned((reg834 || wire842)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1720
#( parameter param1812 = (({{(8'hab), (~&(7'h43))}, (((8'hba) ? (8'hb9) : (8'hb1)) ? {(8'h9d), (8'hb0)} : ((8'haa) == (8'hb7)))} ? ((~^((8'hb0) ? (8'hb7) : (7'h41))) ^~ {((8'hbc) >>> (8'hbd))}) : (((~^(8'ha4)) ? (8'ha1) : (+(8'hbd))) ? (((7'h40) ? (8'hb8) : (8'hb5)) ? {(7'h43)} : {(7'h42), (8'hb1)}) : (((8'hba) ? (8'hbe) : (8'ha9)) ? (-(7'h40)) : {(8'ha7), (8'ha1)}))) ? {(8'hb1), (((^(8'ha5)) == ((8'hbd) ? (8'hb0) : (8'hb4))) - (((8'ha6) ? (8'hbb) : (8'hb4)) < {(8'hb7)}))} : {({(^~(8'ha2)), ((8'hb4) ? (8'hb1) : (8'hbf))} != ((-(8'hbc)) ^~ (~^(7'h43)))), {(((8'h9d) ? (8'ha5) : (8'hb4)) ? (~|(8'ha5)) : ((7'h41) - (8'ha1))), (((7'h41) > (8'h9f)) ? {(8'hbe), (7'h40)} : ((7'h44) | (8'ha9)))}}) )
(y, clk, wire1721, wire1722, wire1723, wire1724, wire1725);
  output wire [(32'h273):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire1721;
  input wire signed [(4'hc):(1'h0)] wire1722;
  input wire signed [(5'h13):(1'h0)] wire1723;
  input wire [(5'h14):(1'h0)] wire1724;
  input wire signed [(4'ha):(1'h0)] wire1725;
  reg signed [(3'h7):(1'h0)] reg1811 = (1'h0);
  reg [(4'h9):(1'h0)] reg1810 = (1'h0);
  reg [(3'h7):(1'h0)] reg1809 = (1'h0);
  reg [(4'hc):(1'h0)] reg1808 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1807 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1806 = (1'h0);
  reg [(3'h6):(1'h0)] reg1805 = (1'h0);
  reg [(4'h8):(1'h0)] reg1804 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1803 = (1'h0);
  reg [(4'ha):(1'h0)] reg1802 = (1'h0);
  reg [(5'h15):(1'h0)] reg1801 = (1'h0);
  reg [(3'h7):(1'h0)] reg1800 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1799 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1798 = (1'h0);
  reg [(4'hb):(1'h0)] reg1797 = (1'h0);
  reg [(4'hb):(1'h0)] reg1796 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1795 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1794 = (1'h0);
  reg [(3'h6):(1'h0)] reg1793 = (1'h0);
  reg [(4'h9):(1'h0)] reg1792 = (1'h0);
  reg [(2'h3):(1'h0)] reg1791 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1790 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1789 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1788 = (1'h0);
  reg [(5'h13):(1'h0)] reg1787 = (1'h0);
  reg [(4'hf):(1'h0)] reg1786 = (1'h0);
  reg [(2'h2):(1'h0)] reg1785 = (1'h0);
  wire [(4'hd):(1'h0)] wire1784;
  wire signed [(3'h4):(1'h0)] wire1783;
  wire signed [(5'h10):(1'h0)] wire1782;
  wire signed [(4'ha):(1'h0)] wire1781;
  wire [(4'hc):(1'h0)] wire1780;
  reg signed [(3'h5):(1'h0)] reg1779 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1778 = (1'h0);
  wire [(4'hc):(1'h0)] wire1777;
  wire [(3'h6):(1'h0)] wire1776;
  wire [(4'h8):(1'h0)] wire1775;
  wire signed [(3'h7):(1'h0)] wire1774;
  wire signed [(4'he):(1'h0)] wire1773;
  wire signed [(4'he):(1'h0)] wire1772;
  reg signed [(4'hf):(1'h0)] reg1726 = (1'h0);
  reg [(2'h3):(1'h0)] reg1727 = (1'h0);
  reg [(4'hd):(1'h0)] reg1728 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1729 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire1730;
  reg [(5'h14):(1'h0)] reg1731 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1732 = (1'h0);
  reg [(4'ha):(1'h0)] reg1733 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1734 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1735 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1736 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1737 = (1'h0);
  reg [(4'ha):(1'h0)] reg1738 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1739 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1740 = (1'h0);
  reg [(4'ha):(1'h0)] reg1741 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1742 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1770;
  assign y = {reg1811,
                 reg1810,
                 reg1809,
                 reg1808,
                 reg1807,
                 reg1806,
                 reg1805,
                 reg1804,
                 reg1803,
                 reg1802,
                 reg1801,
                 reg1800,
                 reg1799,
                 reg1798,
                 reg1797,
                 reg1796,
                 reg1795,
                 reg1794,
                 reg1793,
                 reg1792,
                 reg1791,
                 reg1790,
                 reg1789,
                 reg1788,
                 reg1787,
                 reg1786,
                 reg1785,
                 wire1784,
                 wire1783,
                 wire1782,
                 wire1781,
                 wire1780,
                 reg1779,
                 reg1778,
                 wire1777,
                 wire1776,
                 wire1775,
                 wire1774,
                 wire1773,
                 wire1772,
                 reg1726,
                 reg1727,
                 reg1728,
                 reg1729,
                 wire1730,
                 reg1731,
                 reg1732,
                 reg1733,
                 reg1734,
                 reg1735,
                 reg1736,
                 reg1737,
                 reg1738,
                 reg1739,
                 reg1740,
                 reg1741,
                 reg1742,
                 wire1770,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1726 <= $unsigned(wire1723[(5'h13):(4'he)]);
      reg1727 <= (^~(($signed((wire1725 ?
              wire1724 : reg1726)) > ((wire1722 | wire1725) ?
              $unsigned((8'hb5)) : (-wire1723))) ?
          $signed((+$signed(wire1724))) : $signed(wire1725)));
      reg1728 <= ((~|$signed((|reg1727[(1'h0):(1'h0)]))) ?
          (8'hbc) : (^~wire1721[(2'h2):(2'h2)]));
      reg1729 <= (^(reg1726 ?
          (~$unsigned({wire1725})) : (wire1725[(2'h2):(1'h1)] * (-((8'hb3) ?
              wire1721 : wire1722)))));
    end
  assign wire1730 = $unsigned((((|(8'ha3)) <<< {reg1727,
                            reg1727[(2'h3):(1'h1)]}) ?
                        $signed(reg1726[(4'he):(4'ha)]) : ({wire1722[(4'h9):(3'h4)],
                            (^wire1721)} >= $signed((wire1724 >= reg1729)))));
  always
    @(posedge clk) begin
      reg1731 <= (((^~(^~$signed(reg1728))) ?
              $unsigned((&wire1725)) : ((~^wire1721) ?
                  (^{(8'hb8)}) : ($unsigned(wire1725) ?
                      (wire1725 + wire1724) : reg1728))) ?
          {$signed($signed((~|wire1725))),
              wire1725[(2'h3):(1'h1)]} : $signed((wire1725 << $unsigned($signed(wire1730)))));
      reg1732 <= $signed($unsigned(($unsigned(reg1728[(3'h7):(1'h1)]) ?
          wire1723[(1'h1):(1'h0)] : $unsigned((wire1723 && reg1727)))));
      reg1733 <= reg1731;
      if ((wire1725 ^~ ($signed(wire1722[(3'h7):(3'h6)]) ?
          reg1726[(3'h4):(1'h1)] : ((-(wire1721 ?
              (7'h42) : wire1730)) < reg1733[(3'h4):(3'h4)]))))
        begin
          if ((reg1727 && (({{wire1724}, wire1730} ?
                  {{reg1731, (8'haf)}} : wire1721[(2'h3):(1'h0)]) ?
              {(reg1727 ? ((8'hae) ~^ (8'h9f)) : wire1724)} : {(-wire1722),
                  (&$unsigned(wire1724))})))
            begin
              reg1734 <= $signed(($signed({reg1732}) >= (+((reg1732 ?
                  wire1722 : reg1727) - (wire1725 ? reg1727 : wire1724)))));
              reg1735 <= $unsigned(($signed((&$unsigned(wire1721))) + (((reg1727 <<< wire1723) && (~&wire1724)) << ({wire1725,
                      reg1728} ?
                  (|wire1721) : (reg1728 >= wire1721)))));
              reg1736 <= reg1734[(4'hf):(1'h1)];
            end
          else
            begin
              reg1734 <= (~&({$unsigned(reg1735[(3'h4):(2'h3)]),
                  $unsigned((wire1724 + reg1726))} < {reg1728[(3'h4):(2'h3)]}));
              reg1735 <= $unsigned($signed(reg1727[(1'h1):(1'h1)]));
            end
          reg1737 <= (!(({{wire1721}, $unsigned(reg1732)} ?
                  reg1729 : reg1733[(4'h9):(3'h4)]) ?
              reg1731 : (($signed(wire1721) != wire1730[(4'he):(4'ha)]) | (~&reg1735))));
          if ((reg1728[(1'h0):(1'h0)] ?
              ($signed($signed((~&reg1736))) ?
                  (^~reg1734) : $unsigned(reg1728[(4'h9):(1'h1)])) : $signed($unsigned(((^reg1737) >>> reg1732[(1'h1):(1'h0)])))))
            begin
              reg1738 <= $unsigned((+$unsigned($signed($signed(reg1733)))));
              reg1739 <= (reg1735 ? wire1724 : {reg1732});
              reg1740 <= (wire1721[(1'h0):(1'h0)] << (-reg1738));
              reg1741 <= ((8'ha7) ?
                  ($signed(((wire1725 ? reg1732 : wire1722) ?
                      $signed(wire1721) : (7'h44))) - (wire1724 * ((reg1734 ?
                          reg1737 : reg1728) ?
                      $unsigned((8'hb4)) : (wire1730 ?
                          reg1737 : wire1724)))) : {(($unsigned(reg1733) ~^ wire1722) + ((^reg1726) ?
                          $signed(reg1732) : ((8'hb2) << reg1735)))});
            end
          else
            begin
              reg1738 <= $unsigned(($unsigned($signed((reg1738 ?
                  reg1727 : (8'ha3)))) << {($signed(reg1739) ^ $unsigned(wire1722))}));
              reg1739 <= $unsigned(($unsigned(($signed(wire1723) || (8'had))) ?
                  (~|(+reg1736[(2'h3):(1'h1)])) : {wire1722,
                      reg1732[(4'hc):(4'hc)]}));
              reg1740 <= (^((-(8'hb6)) - ((!{wire1725}) <<< wire1721)));
            end
        end
      else
        begin
          reg1734 <= wire1722;
          reg1735 <= reg1736[(4'hb):(3'h4)];
          reg1736 <= reg1732[(4'he):(3'h4)];
        end
      reg1742 <= (~|((~^reg1729[(4'h9):(4'h8)]) ?
          {$unsigned((reg1740 ? reg1732 : reg1731)),
              ((+wire1723) ?
                  reg1741[(4'ha):(3'h7)] : reg1727[(2'h3):(1'h1)])} : $signed((^(reg1736 < reg1728)))));
    end
  module1743 modinst1771 (.wire1748(reg1738), .clk(clk), .wire1745(wire1724), .wire1746(reg1734), .wire1747(reg1731), .wire1744(reg1728), .y(wire1770));
  assign wire1772 = ({wire1725[(4'h8):(2'h2)],
                            {(reg1737[(2'h3):(1'h1)] ?
                                    (8'hb9) : $unsigned(reg1736))}} ?
                        (((&$signed(reg1740)) != reg1736) ?
                            reg1739 : $unsigned($unsigned(reg1733))) : {reg1738[(2'h3):(1'h0)],
                            ($signed((wire1721 + reg1727)) >= reg1736)});
  assign wire1773 = (!$signed($unsigned((+((7'h42) ? wire1770 : reg1734)))));
  assign wire1774 = (&$unsigned(($unsigned($signed(reg1733)) != $unsigned((+reg1726)))));
  assign wire1775 = (((~$unsigned((wire1724 ? reg1726 : reg1738))) ?
                            ({((8'ha2) > reg1736),
                                wire1722} && reg1736[(4'ha):(4'h8)]) : $signed($signed(wire1725))) ?
                        wire1774[(3'h5):(1'h0)] : ({((reg1732 - reg1728) ?
                                    (!(8'hab)) : wire1723),
                                (|wire1770[(2'h3):(2'h3)])} ?
                            $unsigned({reg1739}) : $signed((reg1727 ?
                                (^~reg1734) : (reg1736 << reg1735)))));
  assign wire1776 = {$unsigned((((^~wire1724) ?
                            (+wire1730) : (+wire1723)) || $signed(wire1775[(3'h6):(1'h0)]))),
                        (-$signed($signed($unsigned(reg1727))))};
  assign wire1777 = $signed(($unsigned($signed(reg1731[(4'hd):(2'h3)])) ?
                        reg1726[(3'h7):(3'h5)] : (8'hae)));
  always
    @(posedge clk) begin
      reg1778 <= ($unsigned(reg1736[(2'h2):(2'h2)]) ?
          wire1730[(5'h13):(5'h11)] : reg1737[(3'h5):(3'h5)]);
      reg1779 <= reg1728;
    end
  assign wire1780 = (8'hb1);
  assign wire1781 = wire1730[(3'h4):(3'h4)];
  assign wire1782 = wire1774;
  assign wire1783 = $unsigned((~$unsigned(($signed(wire1725) ?
                        wire1722[(2'h2):(2'h2)] : $signed(wire1775)))));
  assign wire1784 = {(-(wire1775[(1'h1):(1'h1)] ?
                            $signed({reg1731,
                                reg1778}) : wire1773[(3'h6):(3'h4)]))};
  always
    @(posedge clk) begin
      reg1785 <= wire1776[(3'h5):(3'h4)];
      reg1786 <= reg1732[(2'h2):(1'h0)];
      reg1787 <= ($unsigned($signed(((~reg1739) ?
              wire1722[(2'h3):(2'h2)] : $signed(wire1777)))) ?
          reg1727 : (!$signed((reg1778[(3'h5):(1'h0)] ?
              (reg1785 == reg1785) : $signed(wire1770)))));
      reg1788 <= reg1728[(3'h6):(3'h5)];
    end
  always
    @(posedge clk) begin
      reg1789 <= (-(^~{(((8'ha5) ? reg1788 : reg1735) ?
              $signed(wire1724) : (~|reg1779))}));
      if ($unsigned((wire1780 << (~|wire1722[(4'h8):(3'h7)]))))
        begin
          if ((((-($signed(reg1741) + (wire1783 ? wire1776 : wire1784))) ?
              reg1736[(4'hb):(3'h7)] : ((8'hab) ?
                  $signed({reg1739, wire1775}) : {((7'h41) ? (8'had) : (8'hbb)),
                      (wire1782 ?
                          wire1724 : wire1784)})) ^ (&($signed(((8'h9d) >> wire1777)) < reg1787[(4'h9):(1'h1)]))))
            begin
              reg1790 <= $signed(wire1781[(2'h2):(1'h1)]);
              reg1791 <= wire1723[(2'h2):(1'h0)];
              reg1792 <= (($signed($signed((reg1789 ~^ reg1742))) ?
                      $unsigned($signed(reg1737[(2'h3):(1'h0)])) : (($signed(reg1787) ?
                              ((8'h9d) ? reg1779 : reg1742) : reg1731) ?
                          reg1727 : {wire1730, wire1724[(1'h1):(1'h0)]})) ?
                  $unsigned(reg1742[(1'h1):(1'h0)]) : wire1782[(5'h10):(3'h4)]);
              reg1793 <= $unsigned({$unsigned($signed({reg1788, wire1723})),
                  reg1729});
              reg1794 <= ($signed((~&reg1736)) ?
                  (reg1737[(3'h5):(1'h1)] ?
                      (&((reg1788 << (8'haf)) - (reg1729 ?
                          wire1781 : reg1792))) : reg1733[(2'h3):(1'h1)]) : (-wire1774[(3'h7):(2'h3)]));
            end
          else
            begin
              reg1790 <= (|reg1739);
              reg1791 <= $unsigned((~|{{(wire1784 ? reg1785 : wire1783),
                      reg1734[(3'h4):(2'h3)]}}));
              reg1792 <= (reg1737 >> $unsigned((($unsigned(wire1721) ?
                  ((7'h44) << reg1787) : reg1734) & $signed((reg1739 << wire1730)))));
              reg1793 <= ($unsigned(reg1729) ?
                  ((^($unsigned(wire1773) << $unsigned(wire1784))) >> $signed((&(~^reg1732)))) : reg1786[(3'h7):(3'h4)]);
            end
        end
      else
        begin
          reg1790 <= $unsigned({reg1733,
              ((~|(reg1790 ^ reg1736)) ?
                  {(&(7'h40)),
                      (reg1788 | wire1730)} : ({wire1723} | reg1785))});
          if ((!(reg1793[(2'h3):(1'h1)] > {$unsigned($signed(wire1721)),
              $signed(((8'hb8) ^ wire1725))})))
            begin
              reg1791 <= $signed($signed({{(~reg1792)},
                  $unsigned(reg1734[(2'h3):(2'h3)])}));
            end
          else
            begin
              reg1791 <= reg1790[(2'h2):(2'h2)];
              reg1792 <= wire1775[(3'h7):(3'h4)];
              reg1793 <= ($unsigned(($signed((reg1794 <= reg1787)) - $signed((~reg1791)))) >>> (reg1785[(1'h1):(1'h1)] ?
                  $unsigned($signed((reg1790 && wire1774))) : ($unsigned((^reg1789)) & (wire1723[(5'h11):(5'h10)] ?
                      reg1785[(1'h1):(1'h0)] : (8'ha4)))));
              reg1794 <= ((&wire1723) ?
                  $unsigned(((~&(~reg1729)) == reg1733)) : $signed((reg1788 ?
                      (-reg1785[(1'h0):(1'h0)]) : $signed($signed((8'hab))))));
              reg1795 <= reg1727[(2'h2):(2'h2)];
            end
          if (($unsigned((($signed(reg1790) ?
                      $signed(reg1729) : (wire1774 | (8'hb5))) ?
                  (&(~|reg1789)) : (~&(reg1791 ~^ reg1779)))) ?
              (~|reg1785) : {$unsigned((~|(reg1726 ? reg1733 : wire1784)))}))
            begin
              reg1796 <= {(~^(wire1770[(3'h4):(2'h2)] ?
                      $signed($unsigned(reg1726)) : wire1722[(1'h1):(1'h1)]))};
              reg1797 <= $unsigned(reg1793);
              reg1798 <= {reg1739[(3'h4):(1'h0)], reg1729[(4'h9):(3'h7)]};
              reg1799 <= ((((~reg1796[(4'h8):(3'h5)]) ?
                      (wire1773[(1'h1):(1'h0)] ?
                          {reg1738, reg1789} : (8'hba)) : {$unsigned(reg1795),
                          (reg1731 << reg1793)}) ?
                  (~(~&(+reg1738))) : {((-reg1797) & $unsigned(reg1727)),
                      reg1793}) & ((&$signed(wire1776[(1'h0):(1'h0)])) ?
                  (&((wire1775 ? (8'hba) : wire1725) ?
                      $unsigned(wire1781) : (wire1783 <<< wire1774))) : ({wire1725[(1'h1):(1'h1)]} ?
                      (((8'had) ?
                          reg1734 : wire1783) << $signed(wire1780)) : (^~reg1733))));
            end
          else
            begin
              reg1796 <= ({$signed($signed((reg1793 + reg1726)))} || reg1787);
            end
          reg1800 <= ((-$signed(($unsigned((8'hb6)) ^~ $signed((8'ha0))))) >>> wire1782[(4'h9):(2'h2)]);
        end
      if (reg1788[(2'h3):(2'h3)])
        begin
          if (reg1796)
            begin
              reg1801 <= $unsigned((-reg1729[(4'h9):(1'h1)]));
              reg1802 <= $unsigned(wire1774[(1'h1):(1'h1)]);
              reg1803 <= wire1781[(3'h6):(1'h0)];
              reg1804 <= reg1736[(3'h4):(2'h3)];
            end
          else
            begin
              reg1801 <= (($unsigned((+$unsigned((7'h42)))) ?
                      $signed(($signed(reg1795) ?
                          $unsigned(reg1739) : (&reg1738))) : (reg1803[(5'h10):(1'h0)] ?
                          {(~^reg1733)} : ((+(8'h9f)) ^~ reg1799))) ?
                  (wire1783[(2'h2):(2'h2)] <<< $unsigned((|$signed(reg1741)))) : (&wire1781));
            end
          reg1805 <= ((!$unsigned({wire1776})) == $signed(($unsigned((^reg1794)) ?
              reg1801 : $signed(reg1787[(5'h13):(4'h8)]))));
        end
      else
        begin
          reg1801 <= {(8'hb0), $unsigned(reg1786)};
          reg1802 <= $signed(reg1788);
          if (($signed($signed($unsigned({reg1788}))) ?
              (~&({(reg1731 ?
                      reg1741 : reg1793)} <<< $signed(reg1794[(1'h1):(1'h0)]))) : $unsigned(reg1796[(3'h7):(3'h5)])))
            begin
              reg1803 <= $unsigned((reg1801[(1'h0):(1'h0)] ?
                  $signed(wire1780[(1'h0):(1'h0)]) : ($unsigned($unsigned(wire1775)) ?
                      reg1804[(3'h5):(1'h1)] : (&reg1742[(2'h3):(2'h2)]))));
              reg1804 <= (~&(8'ha3));
              reg1805 <= reg1739;
              reg1806 <= (-wire1770);
              reg1807 <= (reg1732[(4'hf):(4'hf)] ~^ (^($unsigned($unsigned(reg1792)) ?
                  ($unsigned(reg1787) ?
                      (reg1729 ?
                          wire1783 : reg1728) : wire1722[(1'h0):(1'h0)]) : $signed((reg1733 ?
                      reg1740 : wire1725)))));
            end
          else
            begin
              reg1803 <= reg1789;
              reg1804 <= (&(~wire1784));
              reg1805 <= (($unsigned(reg1805[(1'h1):(1'h0)]) > ($signed($unsigned((8'hb9))) ?
                  ((&(8'haf)) * reg1793) : ($unsigned(wire1783) <<< reg1804))) << (~|reg1800[(3'h4):(3'h4)]));
              reg1806 <= wire1784;
              reg1807 <= ((&wire1781) ?
                  (!{((reg1803 <= (8'ha5)) ?
                          reg1793[(3'h5):(3'h5)] : $unsigned(wire1723)),
                      (~^(-reg1726))}) : reg1739[(2'h3):(1'h0)]);
            end
          reg1808 <= wire1780;
          reg1809 <= wire1775[(3'h7):(2'h2)];
        end
      reg1810 <= wire1725[(4'h9):(2'h2)];
      reg1811 <= {{$signed(reg1808[(4'h8):(3'h6)]), reg1737},
          ((((reg1805 <= (8'hbb)) ? reg1798[(4'h8):(1'h1)] : $signed(reg1798)) ?
              $signed(wire1777) : ((&reg1740) ?
                  $unsigned(reg1803) : (reg1738 + reg1797))) <= (+$unsigned($unsigned(reg1789))))};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1698
#( parameter param1711 = ((8'ha7) >> (((^((8'ha2) ? (8'ha2) : (8'ha1))) << (^(&(8'ha4)))) && ((((8'h9c) ? (8'haa) : (8'hbd)) ^ {(8'hb1), (8'ha7)}) ? (((8'hbf) || (8'hb8)) ? ((7'h44) ? (8'hbf) : (8'hbb)) : {(8'hb0), (8'hbe)}) : (((8'h9f) ? (8'ha8) : (7'h42)) ? {(7'h41), (8'ha2)} : (~|(8'h9f))))))
, parameter param1712 = (~|{(!(((8'h9f) ? param1711 : param1711) ? (|param1711) : param1711))}) )
(y, clk, wire1702, wire1701, wire1700, wire1699);
  output wire [(32'h63):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire1702;
  input wire signed [(4'hf):(1'h0)] wire1701;
  input wire [(4'hd):(1'h0)] wire1700;
  input wire [(4'hc):(1'h0)] wire1699;
  wire [(4'hd):(1'h0)] wire1710;
  wire [(4'ha):(1'h0)] wire1709;
  wire [(2'h3):(1'h0)] wire1708;
  wire [(3'h7):(1'h0)] wire1707;
  wire [(3'h4):(1'h0)] wire1706;
  wire signed [(5'h15):(1'h0)] wire1705;
  wire signed [(5'h13):(1'h0)] wire1704;
  wire [(5'h15):(1'h0)] wire1703;
  assign y = {wire1710,
                 wire1709,
                 wire1708,
                 wire1707,
                 wire1706,
                 wire1705,
                 wire1704,
                 wire1703,
                 (1'h0)};
  assign wire1703 = wire1699;
  assign wire1704 = {(!$signed(((~^wire1703) ?
                            wire1703 : wire1699[(4'hb):(2'h2)])))};
  assign wire1705 = (wire1699[(2'h3):(2'h3)] ?
                        (~$unsigned(((^wire1699) - $signed(wire1703)))) : wire1704[(4'h9):(4'h8)]);
  assign wire1706 = $unsigned($unsigned((~({(7'h40)} <= $signed(wire1705)))));
  assign wire1707 = {wire1699,
                        {$unsigned((((7'h40) <= wire1706) ?
                                $signed((8'hb9)) : (wire1702 << wire1700))),
                            wire1706}};
  assign wire1708 = $unsigned(((((wire1705 ? wire1706 : wire1701) ?
                            $signed(wire1703) : wire1706) ?
                        ({(8'hae)} - (wire1699 ?
                            wire1707 : wire1703)) : (wire1699[(1'h1):(1'h0)] ?
                            (~^wire1702) : $unsigned(wire1703))) - $unsigned(wire1700)));
  assign wire1709 = ($unsigned($signed($signed($unsigned((8'hb7))))) || $signed($signed({wire1701})));
  assign wire1710 = $unsigned($signed(((8'hbd) ?
                        wire1708[(2'h2):(2'h2)] : (!wire1704[(4'hc):(4'hc)]))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1327
#( parameter param1695 = ((((~&((7'h43) >> (8'hb4))) ? (8'ha1) : (~&((8'hba) ? (7'h40) : (8'h9e)))) != ((((8'hb2) ? (8'hb0) : (8'hbb)) ? (8'ha8) : {(8'hae)}) >>> ((~^(8'hbd)) ? {(8'hba), (8'hb2)} : ((8'hb0) ? (8'hb2) : (7'h42))))) - (((~^((8'haa) ? (8'hb0) : (8'hbb))) != (((8'ha8) >>> (8'ha0)) || {(8'hae)})) > (-(~|(^~(7'h44)))))) )
(y, clk, wire1331, wire1330, wire1329, wire1328);
  output wire [(32'h306):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire1331;
  input wire signed [(5'h15):(1'h0)] wire1330;
  input wire signed [(5'h11):(1'h0)] wire1329;
  input wire signed [(5'h14):(1'h0)] wire1328;
  reg signed [(4'hc):(1'h0)] reg1694 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1693 = (1'h0);
  reg [(2'h3):(1'h0)] reg1692 = (1'h0);
  reg [(4'hf):(1'h0)] reg1691 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1690 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1689 = (1'h0);
  wire [(3'h6):(1'h0)] wire1688;
  wire [(4'ha):(1'h0)] wire1687;
  wire signed [(3'h5):(1'h0)] wire1686;
  reg [(4'hb):(1'h0)] reg1685 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1684 = (1'h0);
  reg [(3'h7):(1'h0)] reg1683 = (1'h0);
  reg [(2'h3):(1'h0)] reg1682 = (1'h0);
  reg [(5'h13):(1'h0)] reg1681 = (1'h0);
  reg [(4'he):(1'h0)] reg1680 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1679 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1678 = (1'h0);
  reg [(4'h8):(1'h0)] reg1677 = (1'h0);
  reg [(5'h14):(1'h0)] reg1676 = (1'h0);
  reg [(4'he):(1'h0)] reg1675 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1674 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1673 = (1'h0);
  reg [(4'h8):(1'h0)] reg1672 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1671 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1670 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1669 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1668 = (1'h0);
  reg [(3'h4):(1'h0)] reg1667 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1666 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1665 = (1'h0);
  reg [(4'hb):(1'h0)] reg1664 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1663 = (1'h0);
  reg [(3'h4):(1'h0)] reg1662 = (1'h0);
  reg [(3'h6):(1'h0)] reg1661 = (1'h0);
  reg [(4'hb):(1'h0)] reg1660 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1659 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1658 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1657 = (1'h0);
  reg [(3'h5):(1'h0)] reg1656 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1655 = (1'h0);
  reg [(4'h8):(1'h0)] reg1654 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1653 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1652 = (1'h0);
  reg [(4'hf):(1'h0)] reg1651 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1650 = (1'h0);
  reg [(2'h3):(1'h0)] reg1649 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1648 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1647 = (1'h0);
  reg [(5'h13):(1'h0)] reg1646 = (1'h0);
  reg [(4'hb):(1'h0)] reg1645 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1644 = (1'h0);
  reg [(5'h14):(1'h0)] reg1643 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1642 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1641 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1640 = (1'h0);
  wire [(4'he):(1'h0)] wire1570;
  wire signed [(5'h15):(1'h0)] wire1506;
  wire signed [(5'h11):(1'h0)] wire1372;
  wire signed [(4'hd):(1'h0)] wire1332;
  wire [(4'hb):(1'h0)] wire1543;
  reg signed [(4'he):(1'h0)] reg1572 = (1'h0);
  reg [(3'h6):(1'h0)] reg1573 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1574 = (1'h0);
  wire [(4'hd):(1'h0)] wire1575;
  reg signed [(3'h6):(1'h0)] reg1576 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1577 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1578 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1579 = (1'h0);
  wire [(4'h8):(1'h0)] wire1638;
  assign y = {reg1694,
                 reg1693,
                 reg1692,
                 reg1691,
                 reg1690,
                 reg1689,
                 wire1688,
                 wire1687,
                 wire1686,
                 reg1685,
                 reg1684,
                 reg1683,
                 reg1682,
                 reg1681,
                 reg1680,
                 reg1679,
                 reg1678,
                 reg1677,
                 reg1676,
                 reg1675,
                 reg1674,
                 reg1673,
                 reg1672,
                 reg1671,
                 reg1670,
                 reg1669,
                 reg1668,
                 reg1667,
                 reg1666,
                 reg1665,
                 reg1664,
                 reg1663,
                 reg1662,
                 reg1661,
                 reg1660,
                 reg1659,
                 reg1658,
                 reg1657,
                 reg1656,
                 reg1655,
                 reg1654,
                 reg1653,
                 reg1652,
                 reg1651,
                 reg1650,
                 reg1649,
                 reg1648,
                 reg1647,
                 reg1646,
                 reg1645,
                 reg1644,
                 reg1643,
                 reg1642,
                 reg1641,
                 reg1640,
                 wire1570,
                 wire1506,
                 wire1372,
                 wire1332,
                 wire1543,
                 reg1572,
                 reg1573,
                 reg1574,
                 wire1575,
                 reg1576,
                 reg1577,
                 reg1578,
                 reg1579,
                 wire1638,
                 (1'h0)};
  assign wire1332 = wire1331;
  module1333 modinst1373 (wire1372, clk, wire1328, wire1332, wire1329, wire1330);
  module1374 modinst1507 (.y(wire1506), .wire1376(wire1329), .wire1377(wire1372), .wire1378(wire1331), .clk(clk), .wire1375(wire1330), .wire1379(wire1332));
  module1508 modinst1544 (wire1543, clk, wire1328, wire1372, wire1330, wire1506, wire1329);
  module1545 modinst1571 (wire1570, clk, wire1330, wire1331, wire1328, wire1506, wire1543);
  always
    @(posedge clk) begin
      reg1572 <= (wire1332 > wire1570);
      reg1573 <= $unsigned(((((wire1331 == (8'hb9)) <= $signed(wire1330)) >>> ({wire1332,
          wire1330} >> (wire1570 * wire1331))) + wire1331));
      reg1574 <= ($unsigned($signed(reg1573)) >> ($signed((~|(^~wire1543))) >> ($signed((7'h44)) ?
          (wire1543[(3'h6):(1'h1)] ?
              (~&wire1543) : $signed(wire1570)) : (|(wire1543 ?
              (8'hb7) : wire1330)))));
    end
  assign wire1575 = $unsigned($unsigned({({wire1506, wire1506} ?
                            (reg1573 ?
                                reg1574 : wire1506) : $unsigned(wire1570)),
                        {(^~wire1543)}}));
  always
    @(posedge clk) begin
      reg1576 <= $signed(wire1575[(1'h1):(1'h1)]);
      reg1577 <= ((!$signed((~|$signed(wire1372)))) ?
          $unsigned($unsigned(wire1332)) : (wire1332 <<< (wire1372 & wire1506)));
      reg1578 <= (^((reg1577 <= reg1573) | $unsigned($unsigned($unsigned(wire1372)))));
      reg1579 <= (-{reg1576[(3'h6):(2'h2)]});
    end
  module1580 modinst1639 (.clk(clk), .wire1583(reg1577), .wire1584(reg1579), .wire1581(reg1574), .wire1582(wire1330), .y(wire1638), .wire1585(wire1543));
  always
    @(posedge clk) begin
      if (wire1543)
        begin
          reg1640 <= (!$signed((wire1328[(4'hb):(2'h2)] <<< ((wire1331 ?
              wire1328 : wire1543) >>> $unsigned(wire1332)))));
          reg1641 <= {($signed(((8'ha0) ? {reg1572} : $signed(wire1329))) ?
                  (^~((&reg1579) ~^ reg1576)) : ($signed(wire1330) > wire1328))};
          if (wire1331[(3'h4):(1'h1)])
            begin
              reg1642 <= (reg1578[(4'hf):(4'hd)] ^ $unsigned(wire1543[(4'h9):(2'h3)]));
              reg1643 <= (^($signed({(reg1579 && reg1641)}) & (((wire1506 < wire1330) + (wire1506 ~^ (8'hae))) ?
                  ($signed(reg1642) ?
                      (^~wire1638) : $unsigned((8'ha2))) : $signed(((8'had) ?
                      wire1575 : (7'h40))))));
            end
          else
            begin
              reg1642 <= ($signed((~(-reg1642[(3'h4):(2'h2)]))) ?
                  (~^$signed(reg1576)) : $signed($unsigned(((-reg1579) ?
                      (reg1577 >> reg1573) : $signed(reg1577)))));
              reg1643 <= wire1506[(4'h9):(4'h9)];
            end
          if ((~|(((reg1578 & (reg1573 ? wire1332 : wire1575)) ?
                  wire1331 : reg1640) ?
              $signed(wire1506[(5'h15):(4'hb)]) : $unsigned(((7'h42) < $signed(reg1578))))))
            begin
              reg1644 <= (8'hac);
              reg1645 <= ({$signed($unsigned(wire1575[(3'h5):(1'h1)])),
                  ((wire1331[(4'hf):(3'h6)] ?
                      ((8'hb8) ? wire1372 : (8'hb0)) : (wire1332 ?
                          reg1574 : reg1573)) >> ({wire1543,
                      reg1642} >= {reg1640,
                      reg1641}))} == ((((^~(8'ha7)) * $signed(wire1331)) ?
                      ((-wire1543) ?
                          (!reg1641) : wire1330) : $signed((^reg1644))) ?
                  wire1570[(2'h2):(1'h1)] : $signed(((reg1574 >> (8'hb1)) ?
                      wire1331 : wire1575[(4'hb):(4'h8)]))));
              reg1646 <= (~^$unsigned(wire1331));
              reg1647 <= (8'hbc);
            end
          else
            begin
              reg1644 <= (~wire1638[(3'h4):(2'h2)]);
            end
        end
      else
        begin
          if (reg1647[(1'h1):(1'h1)])
            begin
              reg1640 <= (((((|(7'h41)) ?
                      $unsigned((7'h42)) : (wire1570 || reg1572)) ?
                  (((8'hbd) ? reg1646 : reg1574) ?
                      ((8'hbc) ?
                          reg1574 : reg1577) : (wire1372 ~^ reg1643)) : {{wire1543}}) ^ $unsigned($signed(reg1579))) < (~|{(~|(reg1646 ?
                      wire1329 : reg1577)),
                  {reg1579[(3'h4):(1'h0)]}}));
              reg1641 <= (reg1577 ?
                  ((^reg1572[(3'h4):(1'h0)]) <= reg1579) : (wire1328[(4'hb):(2'h2)] ~^ (|reg1573)));
            end
          else
            begin
              reg1640 <= $signed($unsigned(reg1644[(1'h0):(1'h0)]));
            end
          reg1642 <= {wire1575[(4'hd):(3'h5)],
              ((($unsigned(reg1645) ?
                  $unsigned(reg1640) : (reg1646 | reg1579)) ^~ ((8'hb5) << $signed((8'hb1)))) >> (reg1578 ?
                  $unsigned(reg1642[(2'h3):(1'h1)]) : reg1643))};
        end
      if ((~(reg1643[(4'h8):(1'h1)] ? wire1372 : (~reg1642[(2'h3):(1'h1)]))))
        begin
          reg1648 <= $signed((!({{reg1644, (7'h41)}, wire1372[(5'h10):(3'h7)]} ?
              (7'h43) : (reg1642 >>> (^~wire1331)))));
          reg1649 <= wire1332[(1'h1):(1'h0)];
          reg1650 <= ($unsigned($unsigned($signed(((7'h40) ?
                  reg1643 : wire1506)))) ?
              reg1573[(1'h0):(1'h0)] : {wire1330[(4'ha):(3'h4)],
                  (((reg1642 ? reg1645 : (8'hae)) & $signed(reg1642)) ?
                      reg1643[(4'hd):(2'h2)] : ($signed(wire1575) ?
                          (reg1578 >>> wire1332) : (8'ha5)))});
          reg1651 <= ((8'hab) + $unsigned($signed(reg1574[(5'h10):(1'h1)])));
          reg1652 <= wire1372;
        end
      else
        begin
          if (reg1652)
            begin
              reg1648 <= {$unsigned((~|$signed(wire1330)))};
              reg1649 <= reg1643;
              reg1650 <= $signed($unsigned($unsigned((-(^~wire1570)))));
              reg1651 <= (reg1648 > ($unsigned($signed($signed((7'h42)))) ?
                  (($signed(reg1651) < wire1331) ?
                      ({wire1330} ?
                          wire1638[(1'h0):(1'h0)] : $unsigned((8'had))) : $signed(reg1578)) : (+($signed(reg1651) & wire1543))));
              reg1652 <= reg1646;
            end
          else
            begin
              reg1648 <= $unsigned($signed((^~$signed((wire1332 ^~ reg1640)))));
              reg1649 <= ({reg1647[(3'h5):(1'h1)]} ?
                  $signed(reg1574) : (reg1572[(1'h1):(1'h0)] == wire1372));
              reg1650 <= (|wire1638);
            end
          reg1653 <= (^~reg1652[(3'h6):(3'h4)]);
          if ((wire1331[(3'h7):(3'h4)] ?
              (8'ha8) : (((8'hb9) ? $unsigned($signed(reg1651)) : reg1652) ?
                  (({reg1644} ?
                      (&reg1651) : (+(8'hbb))) >= {$unsigned(wire1570)}) : (8'ha3))))
            begin
              reg1654 <= (&reg1577[(5'h13):(4'h9)]);
              reg1655 <= (~$signed(($unsigned((reg1578 ? reg1578 : reg1644)) ?
                  $signed((+wire1372)) : (^$signed(wire1638)))));
              reg1656 <= ($unsigned(($unsigned($unsigned(reg1649)) ?
                      (-reg1578[(4'hc):(3'h7)]) : reg1573[(1'h1):(1'h1)])) ?
                  $unsigned(((8'ha9) ?
                      wire1543[(3'h6):(2'h2)] : $unsigned((wire1506 ?
                          (8'ha3) : wire1330)))) : reg1576);
            end
          else
            begin
              reg1654 <= reg1656;
            end
          if ((reg1650[(4'h8):(2'h2)] || (8'h9e)))
            begin
              reg1657 <= (($signed(reg1646) ?
                      reg1652[(1'h1):(1'h0)] : (((~wire1330) >= {wire1575,
                              reg1655}) ?
                          $signed((wire1506 ?
                              reg1648 : (8'had))) : {(~&reg1574)})) ?
                  wire1638 : reg1651[(1'h1):(1'h1)]);
              reg1658 <= reg1642[(3'h4):(2'h2)];
              reg1659 <= ((wire1332[(4'hd):(1'h1)] >>> (~$unsigned(wire1543))) ?
                  (8'hbb) : reg1640);
            end
          else
            begin
              reg1657 <= reg1656[(3'h4):(2'h2)];
              reg1658 <= (reg1645 ?
                  ($signed((!(reg1578 <<< (8'ha9)))) ?
                      $unsigned(wire1372[(5'h11):(4'he)]) : (^$unsigned(reg1659))) : {(((reg1647 != reg1645) ?
                              {reg1574, reg1641} : (!wire1332)) ?
                          $unsigned(reg1645) : ((wire1328 ?
                              (8'ha0) : reg1640) && $unsigned(reg1649))),
                      reg1650});
              reg1659 <= wire1575[(1'h0):(1'h0)];
              reg1660 <= wire1331;
              reg1661 <= $signed({wire1575[(4'hd):(2'h3)]});
            end
          reg1662 <= (reg1645[(3'h7):(2'h2)] ?
              $unsigned((8'hb6)) : reg1660[(3'h7):(1'h0)]);
        end
      if ($unsigned($signed(reg1661[(3'h4):(1'h0)])))
        begin
          if (($signed(reg1659[(4'hb):(2'h3)]) ~^ ($unsigned({(reg1651 > wire1329),
              (^reg1649)}) >> (~(-((8'hb1) ? reg1654 : reg1656))))))
            begin
              reg1663 <= (~(8'hbd));
              reg1664 <= (8'ha7);
            end
          else
            begin
              reg1663 <= reg1647[(3'h4):(1'h1)];
              reg1664 <= reg1576;
              reg1665 <= (^({$signed($unsigned(reg1655))} ?
                  reg1647[(2'h3):(1'h0)] : {((reg1647 ? reg1655 : reg1572) ?
                          (-reg1652) : $unsigned(reg1664))}));
              reg1666 <= $signed((8'ha1));
              reg1667 <= reg1657[(4'h8):(3'h5)];
            end
        end
      else
        begin
          reg1663 <= reg1577[(3'h7):(3'h6)];
        end
      reg1668 <= (wire1372[(4'h8):(3'h4)] <<< $signed((!(|(8'hae)))));
      if ((|reg1640[(4'h9):(3'h5)]))
        begin
          if ({reg1661, wire1543})
            begin
              reg1669 <= $signed(({$unsigned((reg1662 ? reg1649 : reg1658)),
                  ({wire1506, (8'haf)} ?
                      $unsigned((8'had)) : (wire1330 && reg1641))} || {$signed({reg1574,
                      reg1662})}));
            end
          else
            begin
              reg1669 <= reg1573[(3'h5):(3'h4)];
              reg1670 <= {(&wire1506[(4'hd):(3'h5)])};
              reg1671 <= wire1331;
              reg1672 <= $unsigned((reg1653[(1'h0):(1'h0)] ?
                  wire1331[(4'hd):(3'h6)] : $unsigned(({(8'hb4),
                      (8'hac)} < reg1662))));
            end
          if ($signed(((+{(reg1649 == reg1577)}) ?
              $signed((8'h9d)) : wire1332[(1'h0):(1'h0)])))
            begin
              reg1673 <= $signed((-reg1644));
              reg1674 <= $unsigned(reg1574[(5'h15):(5'h10)]);
              reg1675 <= reg1649;
            end
          else
            begin
              reg1673 <= {($signed($unsigned({reg1578})) ?
                      $unsigned({(reg1648 && reg1573)}) : reg1670[(1'h1):(1'h1)]),
                  reg1664};
              reg1674 <= (8'hba);
              reg1675 <= (8'haa);
            end
          if ((~reg1643[(5'h11):(4'hd)]))
            begin
              reg1676 <= (&{((reg1666 >>> (reg1640 ?
                      reg1652 : reg1646)) & $signed($signed(reg1657)))});
              reg1677 <= (reg1576 > (8'ha4));
              reg1678 <= ((~&(reg1572[(4'hb):(3'h6)] ?
                  (~((8'hb7) ?
                      wire1332 : reg1677)) : (8'hb7))) < (|(wire1506[(3'h4):(1'h1)] ?
                  reg1644[(2'h2):(2'h2)] : (8'had))));
            end
          else
            begin
              reg1676 <= ($signed($signed(reg1654)) <<< reg1667);
              reg1677 <= $signed(reg1674);
              reg1678 <= (-$signed($signed((^$unsigned(reg1647)))));
            end
          reg1679 <= (reg1649[(1'h0):(1'h0)] ?
              $unsigned(((-reg1659[(5'h10):(2'h3)]) ?
                  wire1638 : reg1678)) : $signed(($unsigned(((8'hbc) - reg1666)) ?
                  $signed(reg1644) : $signed(reg1640))));
        end
      else
        begin
          reg1669 <= $signed((reg1576 ?
              (~^$unsigned(reg1658)) : ($signed(reg1671[(2'h3):(1'h0)]) ?
                  reg1572[(3'h7):(1'h1)] : (wire1506 ?
                      reg1659[(5'h11):(3'h5)] : $signed(wire1328)))));
          reg1670 <= $unsigned($signed($signed({{reg1655}})));
        end
    end
  always
    @(posedge clk) begin
      if (reg1665[(4'hb):(3'h5)])
        begin
          reg1680 <= wire1329[(5'h11):(3'h5)];
          if (reg1663[(1'h1):(1'h1)])
            begin
              reg1681 <= (-(-wire1570[(3'h4):(3'h4)]));
              reg1682 <= wire1332;
              reg1683 <= $signed(reg1680[(2'h2):(1'h1)]);
              reg1684 <= {reg1650[(3'h6):(3'h4)], reg1643[(5'h12):(4'hb)]};
            end
          else
            begin
              reg1681 <= $unsigned(({(^~(reg1577 >>> (8'h9f)))} == $unsigned(($unsigned(wire1328) != (reg1656 > wire1330)))));
              reg1682 <= {{(^reg1678)}};
              reg1683 <= (reg1684 <= $signed((+$unsigned((reg1578 << reg1648)))));
              reg1684 <= (8'ha4);
              reg1685 <= (~&{{$unsigned(reg1659), $unsigned((+reg1645))}});
            end
        end
      else
        begin
          reg1680 <= (~|{$unsigned(((~|reg1678) ?
                  (reg1667 >= reg1648) : (reg1577 ? reg1677 : reg1646)))});
          reg1681 <= $signed((((reg1646[(4'he):(3'h7)] ^ ((8'ha9) ?
              reg1646 : reg1664)) == reg1659) + $signed((|$signed(reg1684)))));
        end
    end
  assign wire1686 = wire1331;
  assign wire1687 = ($unsigned(reg1656[(1'h1):(1'h0)]) ?
                        ((reg1640 ? (~&reg1651) : wire1332) ?
                            (&(~^wire1575[(1'h0):(1'h0)])) : wire1328[(5'h14):(4'ha)]) : (reg1579[(1'h0):(1'h0)] << $unsigned(($unsigned((8'ha5)) ?
                            $signed(reg1680) : $signed((8'hbd))))));
  assign wire1688 = (-wire1506[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg1689 <= wire1686[(2'h3):(1'h0)];
      if (($signed(reg1666) <= (!$unsigned(reg1689))))
        begin
          reg1690 <= $unsigned({reg1685[(2'h3):(1'h1)]});
          reg1691 <= reg1679[(3'h5):(1'h0)];
          reg1692 <= reg1668;
        end
      else
        begin
          if ((^~reg1576[(3'h5):(1'h1)]))
            begin
              reg1690 <= wire1332;
            end
          else
            begin
              reg1690 <= reg1676;
              reg1691 <= ((+reg1572[(3'h7):(3'h7)]) || $unsigned($signed(((reg1675 - reg1691) ?
                  wire1330[(4'hd):(2'h2)] : (reg1670 ? (8'had) : reg1689)))));
              reg1692 <= $unsigned($unsigned(($unsigned($unsigned((8'hb7))) <<< wire1372[(5'h10):(1'h1)])));
            end
        end
      reg1693 <= {(reg1689[(4'hc):(4'h8)] ?
              reg1654[(3'h4):(3'h4)] : {$unsigned((reg1663 << (8'hac)))}),
          reg1661[(3'h6):(1'h0)]};
      reg1694 <= (!(+reg1647));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1156
#( parameter param1307 = (((7'h42) ? ((((8'ha8) | (8'hbf)) - ((8'ha9) ? (8'h9d) : (8'ha7))) | (((8'hbf) ? (8'ha3) : (8'ha2)) - ((7'h44) || (8'hb2)))) : {(((8'ha7) <= (8'hb0)) && (~^(8'haf)))}) ^ (-((((8'hba) == (8'ha0)) <= ((7'h44) - (8'hb4))) ^ (((8'hb1) * (8'h9d)) ? ((8'hb6) ^ (8'ha6)) : {(7'h44)}))))
, parameter param1308 = {param1307} )
(y, clk, wire1161, wire1160, wire1159, wire1158, wire1157);
  output wire [(32'h25c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire1161;
  input wire signed [(4'he):(1'h0)] wire1160;
  input wire [(5'h13):(1'h0)] wire1159;
  input wire signed [(4'ha):(1'h0)] wire1158;
  input wire signed [(5'h14):(1'h0)] wire1157;
  wire [(4'he):(1'h0)] wire1306;
  wire signed [(3'h4):(1'h0)] wire1305;
  wire [(3'h7):(1'h0)] wire1304;
  wire [(2'h3):(1'h0)] wire1303;
  wire signed [(5'h13):(1'h0)] wire1302;
  wire [(4'hc):(1'h0)] wire1301;
  wire [(3'h7):(1'h0)] wire1300;
  wire signed [(5'h13):(1'h0)] wire1299;
  reg [(3'h4):(1'h0)] reg1298 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1297 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1296 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1295 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1294 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1293 = (1'h0);
  reg [(3'h7):(1'h0)] reg1292 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1291 = (1'h0);
  reg [(4'hc):(1'h0)] reg1290 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1289 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire1288;
  wire signed [(5'h10):(1'h0)] wire1287;
  wire signed [(4'ha):(1'h0)] wire1286;
  reg signed [(3'h5):(1'h0)] reg1285 = (1'h0);
  reg [(5'h12):(1'h0)] reg1284 = (1'h0);
  reg [(5'h14):(1'h0)] reg1283 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1282 = (1'h0);
  reg [(4'hb):(1'h0)] reg1281 = (1'h0);
  reg [(4'he):(1'h0)] reg1280 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1279 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1278 = (1'h0);
  reg [(3'h4):(1'h0)] reg1277 = (1'h0);
  reg [(4'h9):(1'h0)] reg1276 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1275 = (1'h0);
  reg [(4'ha):(1'h0)] reg1274 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1273 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1272 = (1'h0);
  reg [(2'h2):(1'h0)] reg1271 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1270 = (1'h0);
  reg [(4'hf):(1'h0)] reg1269 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1268 = (1'h0);
  reg [(5'h13):(1'h0)] reg1267 = (1'h0);
  reg [(4'hd):(1'h0)] reg1266 = (1'h0);
  reg [(4'h9):(1'h0)] reg1265 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1264 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1263 = (1'h0);
  reg [(4'ha):(1'h0)] reg1262 = (1'h0);
  reg [(4'hf):(1'h0)] reg1261 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire1260;
  wire signed [(4'hf):(1'h0)] wire1259;
  wire [(5'h10):(1'h0)] wire1257;
  reg [(4'hd):(1'h0)] reg1220 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1219 = (1'h0);
  wire [(3'h7):(1'h0)] wire1218;
  wire [(5'h13):(1'h0)] wire1217;
  wire signed [(3'h6):(1'h0)] wire1215;
  assign y = {wire1306,
                 wire1305,
                 wire1304,
                 wire1303,
                 wire1302,
                 wire1301,
                 wire1300,
                 wire1299,
                 reg1298,
                 reg1297,
                 reg1296,
                 reg1295,
                 reg1294,
                 reg1293,
                 reg1292,
                 reg1291,
                 reg1290,
                 reg1289,
                 wire1288,
                 wire1287,
                 wire1286,
                 reg1285,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1281,
                 reg1280,
                 reg1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 reg1275,
                 reg1274,
                 reg1273,
                 reg1272,
                 reg1271,
                 reg1270,
                 reg1269,
                 reg1268,
                 reg1267,
                 reg1266,
                 reg1265,
                 reg1264,
                 reg1263,
                 reg1262,
                 reg1261,
                 wire1260,
                 wire1259,
                 wire1257,
                 reg1220,
                 reg1219,
                 wire1218,
                 wire1217,
                 wire1215,
                 (1'h0)};
  module1162 modinst1216 (.wire1163(wire1161), .wire1165(wire1157), .wire1166(wire1158), .y(wire1215), .wire1164(wire1159), .clk(clk));
  assign wire1217 = (wire1160[(4'h8):(3'h4)] ?
                        (($signed({wire1215}) != wire1215) & (!wire1157)) : (~(wire1161 ?
                            (~^{wire1157}) : wire1161[(5'h12):(3'h5)])));
  assign wire1218 = $unsigned({wire1161[(4'hc):(2'h3)]});
  always
    @(posedge clk) begin
      reg1219 <= (^~(($unsigned(wire1161) << ((wire1159 != wire1215) == (8'hb0))) ?
          wire1159 : (^~((|wire1159) ? $unsigned(wire1158) : {(8'hab)}))));
      reg1220 <= wire1218;
    end
  module1221 modinst1258 (.wire1224(wire1217), .y(wire1257), .clk(clk), .wire1223(wire1159), .wire1225(wire1161), .wire1222(wire1157));
  assign wire1259 = wire1257[(3'h7):(1'h1)];
  assign wire1260 = {(wire1161[(3'h6):(1'h1)] ?
                            reg1220 : (({reg1220,
                                wire1161} || $signed((8'haa))) >> (&{wire1218}))),
                        (8'hb7)};
  always
    @(posedge clk) begin
      reg1261 <= {wire1260,
          $unsigned(({{(8'hae)}} ?
              ((wire1159 - wire1218) ?
                  (~&(7'h43)) : $unsigned((7'h44))) : $signed($unsigned(wire1158))))};
      reg1262 <= reg1261;
      if (wire1158[(4'ha):(1'h1)])
        begin
          reg1263 <= (~&(reg1220[(3'h4):(2'h2)] ?
              wire1159 : wire1260[(3'h5):(1'h1)]));
          if ($unsigned($unsigned((({wire1259,
              reg1263} << wire1217[(3'h7):(2'h2)]) + $signed((reg1219 <<< (8'hbe)))))))
            begin
              reg1264 <= (8'hb6);
              reg1265 <= (8'hb8);
              reg1266 <= $signed($signed(($signed($signed(reg1263)) ?
                  reg1265[(1'h1):(1'h1)] : $signed($unsigned((8'h9c))))));
              reg1267 <= $unsigned((((wire1218[(2'h2):(2'h2)] ?
                          (wire1161 ? wire1158 : wire1159) : (wire1260 ?
                              wire1260 : wire1257)) ?
                      wire1260[(4'hc):(4'hb)] : (((8'h9f) >= reg1262) - (~^wire1218))) ?
                  {(+(wire1215 ? (8'ha6) : (8'ha9)))} : (8'hb9)));
              reg1268 <= (7'h44);
            end
          else
            begin
              reg1264 <= {({($unsigned(wire1161) >= $unsigned(reg1267))} << $unsigned(wire1160[(4'ha):(3'h7)]))};
            end
          reg1269 <= {$unsigned(($unsigned({wire1260}) ?
                  $unsigned((wire1160 + reg1262)) : $unsigned((&wire1218))))};
          if (reg1220)
            begin
              reg1270 <= (reg1265[(3'h7):(1'h1)] ?
                  reg1265 : wire1215[(3'h6):(2'h3)]);
              reg1271 <= $signed($signed($unsigned((^~{wire1158}))));
              reg1272 <= ((reg1263[(3'h6):(3'h6)] & wire1218[(2'h3):(2'h2)]) > reg1262);
              reg1273 <= ($unsigned({($unsigned(wire1260) ?
                          (reg1265 ?
                              wire1218 : reg1266) : $unsigned((8'haa)))}) ?
                  reg1220 : {$signed(reg1271[(1'h1):(1'h0)])});
              reg1274 <= (^($unsigned($signed($unsigned(reg1220))) >= ((wire1161 ~^ $unsigned(wire1161)) << wire1157[(4'hd):(2'h2)])));
            end
          else
            begin
              reg1270 <= ((~{$signed(((8'hb8) > reg1269))}) || $signed(reg1268));
              reg1271 <= (8'h9d);
            end
        end
      else
        begin
          if (reg1267[(4'h9):(4'h9)])
            begin
              reg1263 <= reg1261;
            end
          else
            begin
              reg1263 <= reg1267[(3'h5):(1'h0)];
              reg1264 <= reg1268;
            end
          reg1265 <= {reg1261[(3'h6):(3'h6)]};
          if (($unsigned({$signed($signed(wire1218)),
                  $unsigned(reg1272[(3'h7):(2'h2)])}) ?
              ((8'ha7) - wire1260[(3'h4):(2'h2)]) : $signed((reg1265 * $unsigned((reg1267 ?
                  wire1260 : wire1159))))))
            begin
              reg1266 <= $signed(reg1267[(2'h3):(1'h0)]);
            end
          else
            begin
              reg1266 <= reg1266[(3'h5):(3'h5)];
            end
          if ($signed($unsigned((reg1220[(3'h4):(2'h2)] ?
              $unsigned($unsigned(wire1218)) : reg1264[(4'hb):(1'h1)]))))
            begin
              reg1267 <= (|(!$signed(wire1217)));
            end
          else
            begin
              reg1267 <= wire1157;
              reg1268 <= (&({reg1261[(3'h7):(2'h3)]} ?
                  reg1270[(4'hb):(3'h6)] : reg1261[(4'he):(3'h6)]));
              reg1269 <= wire1161;
              reg1270 <= $unsigned(wire1159[(2'h3):(1'h1)]);
              reg1271 <= reg1261;
            end
          if (wire1259)
            begin
              reg1272 <= ($unsigned($unsigned((~(wire1161 ?
                  (8'h9d) : reg1261)))) >= (|$signed({$signed(wire1257)})));
              reg1273 <= $unsigned(((8'h9d) + wire1158));
              reg1274 <= (~&wire1218[(3'h6):(3'h6)]);
              reg1275 <= ($signed((((reg1272 ? reg1272 : wire1217) ?
                      reg1219 : (8'ha5)) ^~ $signed($unsigned(reg1266)))) ?
                  reg1220 : reg1220);
            end
          else
            begin
              reg1272 <= {wire1157[(2'h2):(1'h0)],
                  (wire1157[(5'h12):(4'h9)] && (!reg1269[(4'hd):(4'h9)]))};
              reg1273 <= (((8'hb7) ?
                  (!($unsigned((8'ha4)) ?
                      {reg1268} : $unsigned(reg1269))) : $signed((^~wire1218[(2'h2):(1'h0)]))) + reg1264[(4'h8):(2'h2)]);
              reg1274 <= (reg1267[(3'h5):(1'h0)] ?
                  reg1271 : reg1267[(3'h6):(2'h2)]);
              reg1275 <= reg1268[(4'h9):(3'h6)];
            end
        end
      if (wire1217)
        begin
          if ((reg1262 ? (~&({reg1219} < wire1215[(1'h0):(1'h0)])) : (8'ha6)))
            begin
              reg1276 <= ($unsigned($unsigned($signed((wire1257 ?
                      reg1219 : reg1271)))) ?
                  wire1159 : {reg1219[(1'h0):(1'h0)]});
              reg1277 <= {((~(8'ha1)) ^~ $unsigned(wire1160)),
                  ($signed(reg1220) ?
                      $unsigned((((8'ha8) ?
                          reg1264 : wire1218) ^ (wire1157 ~^ wire1218))) : {wire1158[(4'h9):(1'h1)],
                          (reg1270 || {(8'hbb), reg1261})})};
              reg1278 <= (reg1261[(4'he):(3'h6)] << $unsigned(wire1217));
              reg1279 <= wire1158[(2'h2):(2'h2)];
              reg1280 <= ($unsigned({$unsigned($unsigned(reg1220))}) ?
                  $unsigned(reg1266) : (((&(reg1219 <= reg1271)) - $unsigned((8'hb8))) <<< (~^(8'had))));
            end
          else
            begin
              reg1276 <= (reg1279 ? $signed(reg1276) : wire1260);
            end
          reg1281 <= wire1260[(1'h0):(1'h0)];
          if ($unsigned((-wire1158)))
            begin
              reg1282 <= (8'hb3);
            end
          else
            begin
              reg1282 <= {((~|reg1271) ?
                      ((+((8'hb7) ? wire1260 : wire1259)) ?
                          ((|wire1217) ?
                              $unsigned((8'hb8)) : (reg1264 <= reg1282)) : ((reg1271 & reg1269) ?
                              $signed(reg1264) : $unsigned(reg1265))) : $signed($unsigned(reg1271))),
                  ((!(reg1278[(2'h2):(2'h2)] ?
                      (reg1281 < reg1268) : (reg1219 ?
                          reg1220 : reg1273))) || (~|(8'haf)))};
              reg1283 <= ((({(reg1275 ? reg1268 : reg1277), (+reg1279)} ?
                          (~|(reg1282 & reg1274)) : $signed(reg1280)) ?
                      reg1268[(4'h9):(3'h5)] : $signed((~|reg1266))) ?
                  (reg1267[(5'h12):(1'h0)] ^~ {({wire1161} ?
                          $signed(reg1270) : $unsigned(wire1215))}) : reg1274[(4'h9):(2'h2)]);
              reg1284 <= (($unsigned(reg1262) ?
                      {((&(8'hbe)) ?
                              {reg1261,
                                  reg1281} : reg1281)} : $unsigned((8'ha5))) ?
                  (~^$unsigned((~^(reg1267 ? wire1257 : reg1280)))) : wire1158);
            end
        end
      else
        begin
          reg1276 <= (reg1270 ?
              $signed($unsigned(wire1215[(3'h4):(3'h4)])) : wire1260);
        end
      reg1285 <= (^$unsigned(wire1157[(4'hd):(4'hb)]));
    end
  assign wire1286 = (((^~({(8'hbc), reg1270} ?
                            $unsigned(wire1160) : $unsigned(reg1271))) + (reg1279 ?
                            {$unsigned(reg1281), (^reg1219)} : (!(reg1263 ?
                                wire1259 : (8'hb6))))) ?
                        ({reg1282,
                                ($unsigned(reg1272) ?
                                    (-reg1269) : (reg1269 ^ wire1259))} ?
                            wire1257 : $unsigned(wire1215)) : $unsigned((~&reg1279)));
  assign wire1287 = $signed($signed((wire1259 ?
                        wire1260 : reg1274[(3'h5):(3'h4)])));
  assign wire1288 = (~^wire1259);
  always
    @(posedge clk) begin
      if (($signed({(reg1282[(4'h9):(3'h6)] ?
                  (wire1160 ? reg1262 : reg1281) : $unsigned(wire1257))}) ?
          reg1274[(1'h1):(1'h0)] : reg1285))
        begin
          reg1289 <= {reg1264[(2'h3):(2'h2)]};
          reg1290 <= reg1266;
          reg1291 <= $unsigned($unsigned($signed(reg1273)));
        end
      else
        begin
          reg1289 <= $signed(wire1159[(3'h6):(2'h2)]);
          if (({(($signed(reg1270) == {(8'haa)}) ?
                  ((8'ha0) + ((8'ha1) >>> wire1218)) : (8'hba)),
              $unsigned(($unsigned(reg1276) ?
                  (8'hbc) : (+reg1272)))} >> (-((+wire1161) || wire1160[(1'h1):(1'h1)]))))
            begin
              reg1290 <= (~|$unsigned($signed($unsigned($signed(reg1278)))));
            end
          else
            begin
              reg1290 <= (+$signed((reg1266[(4'h9):(1'h1)] ?
                  $unsigned(reg1274[(4'h9):(4'h8)]) : reg1290)));
            end
          if (reg1269)
            begin
              reg1291 <= wire1287[(4'hc):(3'h4)];
              reg1292 <= (~|(+{(^{reg1276}),
                  (reg1262 ? (~wire1257) : {(8'hbd)})}));
            end
          else
            begin
              reg1291 <= $unsigned($signed($signed(reg1290[(2'h3):(1'h1)])));
              reg1292 <= ({(((wire1158 ?
                              wire1217 : reg1276) <<< $unsigned(reg1262)) ?
                          reg1261[(2'h3):(1'h1)] : (wire1160[(3'h4):(1'h1)] <<< (reg1273 ?
                              wire1260 : (8'ha7)))),
                      ($signed(reg1270) ?
                          $signed($unsigned(reg1285)) : reg1278)} ?
                  ((reg1272[(2'h3):(1'h1)] ^ $unsigned({reg1280})) <= reg1269) : ((reg1289[(4'hb):(1'h1)] >>> reg1277[(1'h0):(1'h0)]) ?
                      $signed(reg1271) : (^~$signed(reg1281))));
            end
          reg1293 <= {$signed($signed($signed({(8'had)})))};
          reg1294 <= $unsigned((~^reg1219[(1'h0):(1'h0)]));
        end
      reg1295 <= wire1159[(3'h6):(2'h2)];
      reg1296 <= (^(^~wire1286[(2'h3):(1'h1)]));
      reg1297 <= ((({(reg1284 ? wire1286 : reg1274)} ?
                  $signed($unsigned(reg1219)) : ({(8'hac),
                      (8'hba)} > (wire1288 ? reg1266 : reg1293))) ?
              {wire1257} : (((8'had) ? reg1290 : reg1220[(2'h3):(2'h3)]) ?
                  reg1295[(4'ha):(4'h9)] : reg1280[(4'ha):(3'h6)])) ?
          ($unsigned(reg1290) ?
              $signed($signed($unsigned(reg1273))) : wire1257[(4'he):(2'h3)]) : (8'hac));
      reg1298 <= {($signed((wire1157[(2'h3):(2'h2)] ?
              reg1292 : (8'h9f))) >= {reg1264[(2'h2):(2'h2)]}),
          {(~&wire1161[(1'h1):(1'h1)])}};
    end
  assign wire1299 = wire1286[(2'h3):(2'h3)];
  assign wire1300 = ($signed((8'hb5)) ? wire1259 : reg1282[(4'ha):(3'h6)]);
  assign wire1301 = reg1283;
  assign wire1302 = ($unsigned(wire1160[(4'h8):(2'h3)]) <<< reg1281[(3'h4):(1'h0)]);
  assign wire1303 = $unsigned(((8'h9d) ?
                        (~(&{reg1273, wire1158})) : wire1158[(3'h4):(1'h1)]));
  assign wire1304 = (wire1301[(3'h6):(1'h1)] ?
                        reg1272 : $signed(((reg1292[(1'h1):(1'h0)] ?
                                $unsigned((8'hb5)) : (reg1261 <= reg1296)) ?
                            reg1261 : ($unsigned(wire1299) >>> reg1283[(3'h4):(2'h2)]))));
  assign wire1305 = $unsigned({{((&reg1278) >= $unsigned(wire1257)),
                            ((reg1291 << wire1161) ?
                                $signed(reg1274) : (|reg1285))},
                        ($unsigned($signed(reg1264)) ?
                            reg1270 : reg1277[(1'h0):(1'h0)])});
  assign wire1306 = wire1300;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1140
#( parameter param1151 = {(~|(^(((8'hb2) < (8'hbb)) | ((8'ha9) ? (8'h9f) : (8'hbd))))), (~|(^(~(8'hb2))))}
, parameter param1152 = (-param1151) )
(y, clk, wire1144, wire1143, wire1142, wire1141);
  output wire [(32'h43):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire1144;
  input wire signed [(2'h3):(1'h0)] wire1143;
  input wire [(4'h8):(1'h0)] wire1142;
  input wire signed [(3'h6):(1'h0)] wire1141;
  wire signed [(3'h6):(1'h0)] wire1150;
  wire signed [(4'hd):(1'h0)] wire1149;
  wire signed [(4'hf):(1'h0)] wire1148;
  wire [(5'h15):(1'h0)] wire1147;
  wire [(4'h9):(1'h0)] wire1146;
  wire [(2'h2):(1'h0)] wire1145;
  assign y = {wire1150,
                 wire1149,
                 wire1148,
                 wire1147,
                 wire1146,
                 wire1145,
                 (1'h0)};
  assign wire1145 = {$signed((({wire1142} >> wire1142[(4'h8):(3'h5)]) ?
                            (8'hb5) : wire1141[(1'h0):(1'h0)]))};
  assign wire1146 = (~&(-(wire1142[(3'h5):(3'h5)] + ($signed(wire1143) + (&wire1144)))));
  assign wire1147 = $unsigned({$signed((+$unsigned(wire1144)))});
  assign wire1148 = (~wire1147[(3'h5):(3'h4)]);
  assign wire1149 = wire1145;
  assign wire1150 = $signed(wire1147[(5'h10):(4'h8)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1068
#( parameter param1134 = (((~{((8'h9e) >> (8'hb0)), {(8'hba), (8'h9f)}}) ? ((((8'haa) ? (7'h43) : (8'hbe)) - ((8'ha6) | (8'had))) + ((~(7'h42)) ? (&(8'hb5)) : (~^(8'hb3)))) : {(((7'h44) ? (7'h40) : (8'hb2)) << ((7'h40) ? (8'ha4) : (8'hb4)))}) <= (^((((8'h9e) > (8'ha1)) ? ((8'ha8) ? (8'hbd) : (8'hb1)) : ((8'haf) ^~ (8'hac))) ? (!((8'haf) ? (8'hb8) : (8'ha9))) : (8'hbd))))
, parameter param1135 = ((((~^{param1134}) << {{(8'hab)}}) ^ param1134) ? (param1134 ? (&((param1134 ? param1134 : param1134) && param1134)) : param1134) : ((((param1134 != param1134) && param1134) ? (&{param1134, param1134}) : ({(8'hb3)} ^ (param1134 == param1134))) ^ {{param1134}})) )
(y, clk, wire1069, wire1070, wire1071, wire1072);
  output wire [(32'h162):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire1069;
  input wire signed [(5'h13):(1'h0)] wire1070;
  input wire [(5'h14):(1'h0)] wire1071;
  input wire [(4'ha):(1'h0)] wire1072;
  wire [(3'h5):(1'h0)] wire1133;
  wire [(5'h10):(1'h0)] wire1132;
  reg signed [(4'he):(1'h0)] reg1131 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1130 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire1129;
  wire signed [(3'h7):(1'h0)] wire1128;
  wire signed [(4'h8):(1'h0)] wire1127;
  wire signed [(3'h4):(1'h0)] wire1126;
  wire signed [(4'ha):(1'h0)] wire1125;
  wire [(4'hf):(1'h0)] wire1124;
  wire signed [(4'h9):(1'h0)] wire1123;
  wire [(5'h11):(1'h0)] wire1122;
  wire signed [(2'h2):(1'h0)] wire1121;
  wire [(5'h13):(1'h0)] wire1120;
  reg signed [(3'h4):(1'h0)] reg1119 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1118 = (1'h0);
  reg [(5'h11):(1'h0)] reg1117 = (1'h0);
  reg [(4'ha):(1'h0)] reg1116 = (1'h0);
  wire [(4'h9):(1'h0)] wire1115;
  wire signed [(3'h7):(1'h0)] wire1114;
  reg signed [(2'h3):(1'h0)] reg1113 = (1'h0);
  reg [(2'h3):(1'h0)] reg1073 = (1'h0);
  reg [(4'ha):(1'h0)] reg1074 = (1'h0);
  reg [(4'h9):(1'h0)] reg1075 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1076 = (1'h0);
  reg [(4'hc):(1'h0)] reg1077 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1078 = (1'h0);
  reg [(5'h10):(1'h0)] reg1079 = (1'h0);
  reg [(2'h3):(1'h0)] reg1080 = (1'h0);
  reg [(4'h8):(1'h0)] reg1081 = (1'h0);
  reg [(3'h4):(1'h0)] reg1082 = (1'h0);
  reg [(5'h11):(1'h0)] reg1083 = (1'h0);
  wire [(5'h14):(1'h0)] wire1111;
  assign y = {wire1133,
                 wire1132,
                 reg1131,
                 reg1130,
                 wire1129,
                 wire1128,
                 wire1127,
                 wire1126,
                 wire1125,
                 wire1124,
                 wire1123,
                 wire1122,
                 wire1121,
                 wire1120,
                 reg1119,
                 reg1118,
                 reg1117,
                 reg1116,
                 wire1115,
                 wire1114,
                 reg1113,
                 reg1073,
                 reg1074,
                 reg1075,
                 reg1076,
                 reg1077,
                 reg1078,
                 reg1079,
                 reg1080,
                 reg1081,
                 reg1082,
                 reg1083,
                 wire1111,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire1069[(1'h1):(1'h0)])
        begin
          reg1073 <= wire1070;
          reg1074 <= wire1072;
          if ((wire1071[(3'h6):(3'h5)] != $signed($signed(($unsigned(wire1069) > wire1071[(4'h9):(4'h9)])))))
            begin
              reg1075 <= ($signed(wire1069[(1'h0):(1'h0)]) ?
                  {(wire1072[(4'ha):(3'h7)] && (8'hbf)),
                      {$signed((reg1074 | wire1069))}} : ({$signed((wire1071 ?
                          reg1074 : wire1072))} > (8'hbd)));
              reg1076 <= reg1075;
              reg1077 <= $signed((~^reg1075));
              reg1078 <= reg1074[(4'h8):(3'h6)];
            end
          else
            begin
              reg1075 <= $unsigned((~(({(8'haf), wire1071} ?
                  $signed(wire1071) : (reg1075 ?
                      wire1072 : reg1074)) != reg1075[(4'h8):(3'h4)])));
              reg1076 <= reg1075[(3'h5):(3'h4)];
              reg1077 <= {$signed((wire1069[(1'h1):(1'h0)] ?
                      $signed(((8'hb9) <= wire1069)) : reg1078))};
              reg1078 <= {{($unsigned((wire1071 <<< reg1075)) && {{wire1072,
                              wire1069},
                          reg1075[(1'h1):(1'h1)]})}};
              reg1079 <= wire1069;
            end
          reg1080 <= $unsigned(wire1071[(4'ha):(3'h4)]);
          reg1081 <= {($signed(((reg1077 >> reg1078) >= (|reg1073))) ?
                  (7'h41) : {(~$signed(wire1071)), (^~$unsigned(reg1074))}),
              wire1072};
        end
      else
        begin
          reg1073 <= (reg1073[(2'h2):(2'h2)] ?
              (~&wire1072[(1'h0):(1'h0)]) : reg1073[(2'h2):(2'h2)]);
          if ((~&$unsigned((!(wire1071 ? (wire1070 >= reg1081) : wire1072)))))
            begin
              reg1074 <= $unsigned(((reg1080 ?
                      ($signed(wire1072) <<< (!wire1072)) : wire1071[(4'hc):(4'h9)]) ?
                  $unsigned(($unsigned(reg1080) << $unsigned(wire1069))) : $signed(reg1078)));
              reg1075 <= (((($signed(reg1076) ?
                              ((8'ha1) ? reg1077 : reg1073) : reg1074) ?
                          $unsigned($signed(reg1079)) : $signed((reg1078 ^~ reg1073))) ?
                      {((+wire1069) < $signed(reg1081)),
                          (^(~wire1069))} : ($unsigned((&wire1071)) ?
                          {(8'h9c),
                              (~reg1077)} : $unsigned($unsigned(reg1081)))) ?
                  (reg1080[(2'h3):(2'h3)] + ({reg1075[(3'h5):(1'h1)]} >> reg1078[(4'ha):(3'h7)])) : ($signed(reg1074[(4'h9):(1'h0)]) ?
                      (8'ha3) : reg1073[(2'h2):(2'h2)]));
              reg1076 <= (((^reg1075[(2'h3):(1'h1)]) ?
                  wire1071 : (^$unsigned((-wire1071)))) >= (8'ha0));
              reg1077 <= {$signed(wire1070)};
            end
          else
            begin
              reg1074 <= {(reg1077 ?
                      (~($unsigned((8'ha7)) > reg1079)) : {(~^(~reg1079))}),
                  $signed(reg1074[(2'h3):(1'h1)])};
              reg1075 <= (reg1074 ?
                  $unsigned($signed(((wire1072 ?
                      wire1070 : reg1073) ~^ $signed(reg1073)))) : $signed(wire1072));
            end
          if ((({$unsigned(wire1071[(4'h9):(3'h7)]),
              $signed((8'hb0))} || (|$unsigned(reg1075))) <= reg1077))
            begin
              reg1078 <= ($signed(({$unsigned(wire1069)} ?
                  ($unsigned(reg1080) ^ (reg1078 ?
                      reg1076 : reg1080)) : (8'ha7))) ^ {((8'ha8) & $signed(reg1080))});
              reg1079 <= $unsigned(reg1078);
              reg1080 <= reg1073[(1'h1):(1'h1)];
              reg1081 <= (((reg1077 || (8'ha8)) ?
                      {wire1072[(4'ha):(3'h6)],
                          reg1080[(2'h3):(2'h3)]} : $signed(reg1076[(2'h2):(1'h1)])) ?
                  $unsigned(($unsigned((8'ha6)) ?
                      reg1081 : (+wire1069[(2'h3):(1'h1)]))) : ({$signed((wire1071 ?
                          reg1081 : reg1074)),
                      ($signed((8'hab)) ?
                          (|reg1077) : $unsigned(wire1072))} >>> $signed($signed($unsigned((8'ha6))))));
            end
          else
            begin
              reg1078 <= {({((wire1072 ?
                          wire1071 : (8'hb7)) ^ $unsigned(wire1069)),
                      reg1081} - $signed((^~$signed(reg1081))))};
              reg1079 <= $unsigned((~{(|(-reg1079))}));
              reg1080 <= $signed($signed(((~&$signed(reg1073)) ?
                  reg1081[(2'h3):(1'h1)] : wire1071[(1'h1):(1'h1)])));
              reg1081 <= reg1081[(3'h4):(1'h0)];
            end
          reg1082 <= (((reg1075 ?
                  (8'hb7) : $signed(wire1072[(2'h2):(1'h1)])) <<< $signed({$signed((8'ha7))})) ?
              (^~($signed(reg1074) < ((reg1078 ?
                  reg1081 : reg1080) - (wire1070 ?
                  (8'hb8) : reg1073)))) : ((7'h43) ?
                  (~|$signed($signed(reg1080))) : (~$signed($unsigned(reg1078)))));
        end
      reg1083 <= (+reg1074);
    end
  module1084 modinst1112 (wire1111, clk, reg1075, reg1083, wire1070, wire1071, reg1082);
  always
    @(posedge clk) begin
      reg1113 <= $signed($signed($unsigned($unsigned($signed(reg1074)))));
    end
  assign wire1114 = $signed($signed(($signed($unsigned(reg1080)) > (|$signed(reg1078)))));
  assign wire1115 = reg1080[(2'h3):(2'h2)];
  always
    @(posedge clk) begin
      if ((&$unsigned($signed($unsigned((reg1078 ? reg1078 : wire1072))))))
        begin
          reg1116 <= (reg1113[(2'h3):(1'h1)] | $signed($unsigned(reg1073[(2'h2):(1'h0)])));
          reg1117 <= reg1079[(2'h3):(2'h3)];
          reg1118 <= (^$unsigned(reg1080));
        end
      else
        begin
          reg1116 <= reg1116;
          reg1117 <= (&reg1116[(1'h0):(1'h0)]);
          reg1118 <= {$unsigned(reg1082[(1'h1):(1'h1)])};
        end
      reg1119 <= (+$signed(wire1069));
    end
  assign wire1120 = wire1111;
  assign wire1121 = wire1120[(3'h7):(1'h0)];
  assign wire1122 = $signed($signed((8'ha0)));
  assign wire1123 = $unsigned((8'hb4));
  assign wire1124 = (reg1083[(2'h2):(2'h2)] != reg1081);
  assign wire1125 = $signed(reg1074[(4'ha):(3'h6)]);
  assign wire1126 = (wire1115 <<< ($signed(reg1118[(3'h4):(3'h4)]) || reg1078[(1'h1):(1'h1)]));
  assign wire1127 = ((~|$unsigned(reg1078[(1'h0):(1'h0)])) > $unsigned(reg1080));
  assign wire1128 = reg1118;
  assign wire1129 = reg1077[(4'h8):(3'h5)];
  always
    @(posedge clk) begin
      reg1130 <= (8'ha6);
      reg1131 <= ((8'haa) ?
          $unsigned($signed($unsigned(wire1111[(1'h0):(1'h0)]))) : {($signed($signed(reg1074)) <<< ((reg1116 > reg1116) + wire1069[(2'h3):(1'h1)]))});
    end
  assign wire1132 = ((+$signed({wire1115[(1'h0):(1'h0)]})) ?
                        ((+wire1072[(4'ha):(4'ha)]) + {(~|wire1115)}) : $signed($unsigned(reg1131)));
  assign wire1133 = $signed(reg1118[(4'hb):(1'h1)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1013  (y, clk, wire1014, wire1015, wire1016, wire1017);
  output wire [(32'h107):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire1014;
  input wire [(3'h6):(1'h0)] wire1015;
  input wire [(5'h11):(1'h0)] wire1016;
  input wire signed [(4'ha):(1'h0)] wire1017;
  reg signed [(2'h3):(1'h0)] reg1063 = (1'h0);
  reg [(4'hd):(1'h0)] reg1062 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire1018;
  wire [(3'h5):(1'h0)] wire1019;
  wire [(4'h9):(1'h0)] wire1020;
  reg [(3'h4):(1'h0)] reg1021 = (1'h0);
  reg [(4'hd):(1'h0)] reg1022 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1023 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1024 = (1'h0);
  reg [(5'h14):(1'h0)] reg1025 = (1'h0);
  reg [(4'hf):(1'h0)] reg1026 = (1'h0);
  reg [(5'h12):(1'h0)] reg1027 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1028 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1029 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1030 = (1'h0);
  reg [(4'h9):(1'h0)] reg1031 = (1'h0);
  reg [(5'h13):(1'h0)] reg1032 = (1'h0);
  reg [(3'h4):(1'h0)] reg1033 = (1'h0);
  wire [(5'h14):(1'h0)] wire1034;
  wire [(3'h6):(1'h0)] wire1035;
  wire signed [(4'hf):(1'h0)] wire1036;
  wire signed [(3'h4):(1'h0)] wire1037;
  wire [(4'hf):(1'h0)] wire1060;
  assign y = {reg1063,
                 reg1062,
                 wire1018,
                 wire1019,
                 wire1020,
                 reg1021,
                 reg1022,
                 reg1023,
                 reg1024,
                 reg1025,
                 reg1026,
                 reg1027,
                 reg1028,
                 reg1029,
                 reg1030,
                 reg1031,
                 reg1032,
                 reg1033,
                 wire1034,
                 wire1035,
                 wire1036,
                 wire1037,
                 wire1060,
                 (1'h0)};
  assign wire1018 = ($signed({wire1015[(3'h5):(2'h2)]}) ?
                        wire1016 : wire1016[(5'h11):(4'hf)]);
  assign wire1019 = wire1016[(4'h9):(3'h4)];
  assign wire1020 = $signed($unsigned({(8'ha8), wire1015[(2'h2):(1'h1)]}));
  always
    @(posedge clk) begin
      reg1021 <= (((({wire1017, wire1020} || {wire1017, wire1014}) ?
              ((wire1020 ?
                  (8'ha5) : wire1017) ^ (!wire1015)) : {$signed(wire1018)}) ~^ (wire1014 ?
              $signed((wire1019 ?
                  wire1015 : wire1016)) : (wire1017[(3'h6):(1'h1)] ?
                  (wire1018 >= wire1019) : $unsigned((8'hb1))))) ?
          wire1020[(1'h1):(1'h0)] : ($unsigned(wire1016) ?
              (~^((^wire1018) ?
                  $unsigned(wire1019) : wire1014[(3'h6):(3'h4)])) : (-(~|$signed(wire1017)))));
      if (wire1020)
        begin
          reg1022 <= (($unsigned({((8'ha4) || wire1019),
                      (wire1018 ? wire1019 : wire1017)}) ?
                  (wire1018 >>> {(~&wire1019)}) : $unsigned((^{reg1021,
                      reg1021}))) ?
              $signed(wire1017[(3'h5):(3'h4)]) : wire1019[(2'h2):(1'h1)]);
          if (($unsigned((wire1019 ?
                  $unsigned($signed(wire1020)) : (~|(wire1018 * (8'hb4))))) ?
              $unsigned(wire1019[(1'h1):(1'h0)]) : reg1022))
            begin
              reg1023 <= $unsigned(((~&$unsigned($unsigned(wire1014))) ^~ $signed(wire1017)));
              reg1024 <= reg1022;
            end
          else
            begin
              reg1023 <= (^~((8'hac) ?
                  wire1015 : $signed(reg1024[(4'hb):(4'h9)])));
              reg1024 <= wire1016;
              reg1025 <= (8'hb4);
              reg1026 <= (((8'ha6) && $unsigned($signed((!wire1014)))) ?
                  (reg1021[(2'h2):(1'h1)] ?
                      reg1021 : ((((8'h9e) - wire1017) ? reg1021 : (8'h9e)) ?
                          reg1022[(1'h1):(1'h1)] : {(reg1021 << wire1019)})) : reg1024[(4'he):(4'hb)]);
              reg1027 <= wire1017[(1'h1):(1'h0)];
            end
          if ((~(reg1024 > wire1014)))
            begin
              reg1028 <= $unsigned((reg1023 ?
                  wire1019[(1'h0):(1'h0)] : $unsigned($signed(reg1023))));
              reg1029 <= ((8'hb1) ?
                  $unsigned(wire1015) : $unsigned($unsigned($signed((reg1026 != reg1023)))));
              reg1030 <= (($signed($unsigned($signed(wire1020))) | wire1019) || wire1016[(3'h4):(1'h0)]);
              reg1031 <= $unsigned(wire1015);
            end
          else
            begin
              reg1028 <= ((+(~^($unsigned(reg1031) ?
                  $signed(wire1015) : $signed(reg1022)))) >>> reg1024[(4'h9):(3'h7)]);
              reg1029 <= reg1024;
            end
          reg1032 <= (($signed(($signed(reg1031) >>> $signed((8'ha2)))) ?
              (wire1015 <= (^(!wire1014))) : reg1022) & $signed($signed($signed({wire1018,
              wire1019}))));
        end
      else
        begin
          if (($signed(($signed(reg1028) ?
                  ($signed(reg1027) != $unsigned(reg1031)) : reg1024)) ?
              reg1031[(1'h0):(1'h0)] : ($unsigned(((reg1027 ?
                          wire1015 : reg1032) ?
                      reg1028[(3'h7):(3'h6)] : reg1022)) ?
                  ($signed((wire1017 >>> wire1014)) * (^$signed(reg1021))) : $unsigned(reg1032))))
            begin
              reg1022 <= $unsigned(reg1023);
              reg1023 <= {$unsigned((-$unsigned((reg1027 <<< (7'h40)))))};
              reg1024 <= $signed(($unsigned(reg1028) ?
                  reg1026 : $unsigned(reg1021[(2'h2):(1'h1)])));
              reg1025 <= wire1017[(1'h1):(1'h0)];
            end
          else
            begin
              reg1022 <= $signed($unsigned(($unsigned($signed(reg1024)) != (!((7'h42) ?
                  (8'hb2) : reg1032)))));
              reg1023 <= wire1014[(3'h4):(1'h0)];
              reg1024 <= reg1030[(2'h2):(1'h0)];
              reg1025 <= (^~(^~reg1030));
            end
          if ($signed(reg1024))
            begin
              reg1026 <= ((($unsigned((~^(8'h9e))) ?
                          $unsigned(reg1021) : reg1026) ?
                      reg1026 : wire1015) ?
                  wire1014[(1'h1):(1'h0)] : $unsigned(reg1022[(3'h7):(2'h2)]));
            end
          else
            begin
              reg1026 <= (~^($signed(wire1014[(4'hd):(3'h4)]) ?
                  {((reg1023 | wire1019) ?
                          $signed(reg1028) : (reg1023 ? (8'had) : wire1015)),
                      (8'ha0)} : $unsigned(((reg1023 ^ (7'h44)) + reg1031[(4'h8):(3'h4)]))));
              reg1027 <= reg1029[(1'h0):(1'h0)];
            end
        end
      reg1033 <= $unsigned({(+reg1027),
          (|(((8'hb9) ? wire1019 : reg1022) ?
              (reg1026 ? reg1021 : wire1020) : reg1030[(4'he):(2'h2)]))});
    end
  assign wire1034 = (!reg1032);
  assign wire1035 = reg1029[(2'h2):(2'h2)];
  assign wire1036 = $unsigned((($unsigned((wire1019 ? wire1016 : reg1031)) ?
                        $unsigned($signed(wire1017)) : (reg1030 != $signed(reg1023))) ^~ reg1024[(3'h4):(2'h2)]));
  assign wire1037 = ((+$signed(reg1023)) + $unsigned($unsigned({(8'hb2)})));
  module1038 modinst1061 (.wire1043(wire1036), .clk(clk), .wire1040(wire1014), .y(wire1060), .wire1039(wire1019), .wire1042(wire1037), .wire1041(wire1018));
  always
    @(posedge clk) begin
      reg1062 <= wire1020;
      reg1063 <= $signed((-reg1030[(2'h2):(2'h2)]));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1038
#( parameter param1058 = ((~|({((7'h40) >= (8'hbc)), {(8'hb3)}} ? {(^~(8'hb1)), {(8'hb5), (8'hb1)}} : {((8'ha7) ? (8'hae) : (7'h42)), ((8'ha6) != (8'ha0))})) ? (~{((8'h9e) == (~|(7'h42)))}) : {(((~(8'hb6)) ? ((8'hb0) << (8'h9f)) : (^~(8'ha9))) ? (((8'hb3) <<< (8'hb4)) ? ((8'hbf) ? (8'hb4) : (7'h41)) : ((7'h42) ? (7'h42) : (8'ha1))) : (((8'h9c) <<< (8'hbb)) > ((8'ha5) ? (8'ha6) : (8'hae)))), ({((8'ha9) ~^ (8'hb0))} & ({(7'h44)} || ((8'h9f) ? (8'hbd) : (8'hb9))))})
, parameter param1059 = (^param1058) )
(y, clk, wire1043, wire1042, wire1041, wire1040, wire1039);
  output wire [(32'hbc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire1043;
  input wire [(3'h4):(1'h0)] wire1042;
  input wire [(3'h6):(1'h0)] wire1041;
  input wire signed [(4'hb):(1'h0)] wire1040;
  input wire signed [(3'h5):(1'h0)] wire1039;
  wire [(4'hb):(1'h0)] wire1057;
  wire signed [(5'h15):(1'h0)] wire1056;
  wire [(4'he):(1'h0)] wire1055;
  wire [(4'h9):(1'h0)] wire1054;
  wire [(3'h7):(1'h0)] wire1053;
  wire [(5'h15):(1'h0)] wire1052;
  wire signed [(5'h12):(1'h0)] wire1051;
  wire signed [(3'h6):(1'h0)] wire1050;
  wire signed [(5'h11):(1'h0)] wire1049;
  wire [(5'h13):(1'h0)] wire1048;
  wire signed [(2'h2):(1'h0)] wire1047;
  wire [(5'h12):(1'h0)] wire1046;
  wire signed [(2'h3):(1'h0)] wire1045;
  reg [(5'h15):(1'h0)] reg1044 = (1'h0);
  assign y = {wire1057,
                 wire1056,
                 wire1055,
                 wire1054,
                 wire1053,
                 wire1052,
                 wire1051,
                 wire1050,
                 wire1049,
                 wire1048,
                 wire1047,
                 wire1046,
                 wire1045,
                 reg1044,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1044 <= wire1039[(1'h1):(1'h0)];
    end
  assign wire1045 = $unsigned(wire1039[(3'h4):(1'h1)]);
  assign wire1046 = wire1040[(3'h4):(2'h3)];
  assign wire1047 = {(wire1045[(2'h3):(1'h1)] ?
                            $unsigned($unsigned({wire1042})) : {wire1043[(4'hc):(4'ha)]}),
                        (+($signed((wire1043 <= wire1043)) ?
                            $signed((wire1046 ?
                                wire1039 : wire1042)) : $signed($unsigned(wire1042))))};
  assign wire1048 = $unsigned(((wire1042[(1'h1):(1'h0)] ?
                        $unsigned({wire1046,
                            (8'hb4)}) : ($unsigned(wire1046) ^ $signed((7'h43)))) + (~|(8'hb6))));
  assign wire1049 = wire1042;
  assign wire1050 = $unsigned((({(8'hbb)} || $signed((~^wire1042))) < $signed(wire1039[(2'h3):(1'h1)])));
  assign wire1051 = wire1042[(3'h4):(1'h0)];
  assign wire1052 = ($signed((((|wire1041) <= {wire1051}) ?
                        wire1051[(1'h0):(1'h0)] : (wire1043[(1'h1):(1'h1)] ?
                            (wire1042 + wire1049) : {wire1045,
                                wire1039}))) + (~(~&wire1045[(2'h3):(2'h2)])));
  assign wire1053 = (($unsigned((-(8'hb7))) ?
                            ((wire1041 ?
                                    $unsigned(wire1045) : $unsigned(wire1040)) ?
                                (~|(wire1045 ?
                                    wire1042 : wire1042)) : wire1039) : wire1039) ?
                        (($unsigned($unsigned(reg1044)) ?
                            (wire1047 >> wire1052) : $signed({wire1052,
                                (8'ha8)})) * (~(8'hb2))) : $signed($signed($signed((^wire1048)))));
  assign wire1054 = $unsigned($unsigned($unsigned(((~^wire1046) >> wire1051[(3'h5):(3'h5)]))));
  assign wire1055 = $signed(wire1052[(1'h1):(1'h1)]);
  assign wire1056 = wire1054[(3'h7):(3'h6)];
  assign wire1057 = wire1041;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1084  (y, clk, wire1089, wire1088, wire1087, wire1086, wire1085);
  output wire [(32'hd1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire1089;
  input wire [(5'h11):(1'h0)] wire1088;
  input wire signed [(5'h13):(1'h0)] wire1087;
  input wire signed [(5'h14):(1'h0)] wire1086;
  input wire signed [(3'h4):(1'h0)] wire1085;
  wire [(4'he):(1'h0)] wire1110;
  wire signed [(4'hc):(1'h0)] wire1109;
  reg [(4'h8):(1'h0)] reg1108 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1107 = (1'h0);
  reg [(5'h12):(1'h0)] reg1106 = (1'h0);
  wire [(3'h6):(1'h0)] wire1105;
  reg [(3'h5):(1'h0)] reg1104 = (1'h0);
  reg [(4'hb):(1'h0)] reg1103 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1102 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1101 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1100 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1099 = (1'h0);
  reg [(4'h8):(1'h0)] reg1098 = (1'h0);
  reg [(3'h4):(1'h0)] reg1097 = (1'h0);
  reg [(3'h6):(1'h0)] reg1096 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1095 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1094;
  wire signed [(4'hb):(1'h0)] wire1093;
  wire [(4'ha):(1'h0)] wire1092;
  wire [(2'h3):(1'h0)] wire1091;
  wire signed [(4'h9):(1'h0)] wire1090;
  assign y = {wire1110,
                 wire1109,
                 reg1108,
                 reg1107,
                 reg1106,
                 wire1105,
                 reg1104,
                 reg1103,
                 reg1102,
                 reg1101,
                 reg1100,
                 reg1099,
                 reg1098,
                 reg1097,
                 reg1096,
                 reg1095,
                 wire1094,
                 wire1093,
                 wire1092,
                 wire1091,
                 wire1090,
                 (1'h0)};
  assign wire1090 = (~&wire1089[(1'h1):(1'h0)]);
  assign wire1091 = (~^$signed($signed($signed($signed(wire1089)))));
  assign wire1092 = (wire1090[(1'h1):(1'h1)] ^~ $unsigned(wire1089));
  assign wire1093 = (-{wire1086});
  assign wire1094 = $signed(wire1087);
  always
    @(posedge clk) begin
      if ((^$signed({wire1090, wire1087[(4'h8):(3'h4)]})))
        begin
          if (((|$unsigned(wire1091[(1'h0):(1'h0)])) != wire1091[(2'h2):(2'h2)]))
            begin
              reg1095 <= $signed($unsigned((~|wire1089[(1'h1):(1'h1)])));
            end
          else
            begin
              reg1095 <= wire1085;
              reg1096 <= (({{(-wire1093)}} ?
                  reg1095[(4'ha):(4'h9)] : (|wire1091)) <= (~|wire1087));
              reg1097 <= reg1095;
            end
          reg1098 <= (((-($signed(wire1085) ?
                      (reg1095 << reg1096) : (!wire1088))) ?
                  (&wire1085[(1'h0):(1'h0)]) : wire1088) ?
              (~|{wire1089[(3'h4):(2'h2)]}) : (reg1097[(1'h1):(1'h1)] ?
                  $signed(wire1085[(1'h0):(1'h0)]) : $signed($unsigned(reg1095[(3'h4):(3'h4)]))));
          if (($signed(wire1092[(4'h9):(4'h9)]) ?
              reg1097 : ($unsigned(reg1096) != $signed(wire1093[(4'ha):(3'h4)]))))
            begin
              reg1099 <= {((~$unsigned((reg1095 > wire1090))) && (~^(wire1093 ?
                      (wire1087 ? wire1087 : reg1095) : (|reg1096))))};
              reg1100 <= (((wire1089[(3'h4):(1'h1)] ?
                          ($signed(wire1088) >>> reg1096[(2'h2):(1'h0)]) : ($unsigned(reg1096) == {reg1098})) ?
                      $unsigned((!$unsigned(wire1086))) : (((&wire1088) << (reg1096 ?
                              reg1096 : wire1094)) ?
                          (~^(wire1089 ? wire1093 : wire1092)) : wire1088)) ?
                  ($signed((((8'ha2) | wire1093) <= (~reg1096))) >>> ((((8'hba) ?
                          wire1092 : reg1098) | wire1089[(3'h7):(3'h7)]) ?
                      (wire1090 ~^ $unsigned(wire1089)) : ((wire1087 ?
                              (8'hb9) : wire1090) ?
                          $unsigned(reg1099) : $signed(wire1088)))) : (-(({wire1090} ^~ $unsigned(wire1085)) ?
                      (wire1085[(1'h1):(1'h0)] ?
                          (wire1086 ~^ wire1091) : (wire1088 ?
                              wire1087 : wire1092)) : wire1085)));
              reg1101 <= $signed(((^({wire1087, wire1093} ?
                  $signed(wire1085) : (&reg1099))) * wire1086));
            end
          else
            begin
              reg1099 <= (~$signed($unsigned($signed($signed(reg1099)))));
              reg1100 <= $unsigned($unsigned(($signed(wire1087) * $signed($signed((8'hb3))))));
            end
          reg1102 <= $signed({reg1100[(3'h6):(3'h6)]});
        end
      else
        begin
          reg1095 <= (wire1089 ?
              (wire1086[(5'h10):(4'hd)] >> wire1090[(3'h5):(1'h0)]) : ((~(~|$unsigned(wire1089))) ^ $signed(((+(8'ha0)) ?
                  (~|reg1098) : $unsigned(wire1091)))));
          reg1096 <= ((!((^~(+reg1102)) >> reg1095)) ? wire1093 : (8'hb0));
          reg1097 <= $unsigned($signed((reg1095[(4'he):(1'h1)] ?
              $unsigned(wire1091) : wire1093)));
          if ($unsigned((wire1085 <= $signed(reg1095))))
            begin
              reg1098 <= ($signed((wire1094[(4'hd):(3'h5)] ?
                      (wire1090 != wire1087[(4'ha):(2'h3)]) : ($signed((8'hb2)) ?
                          $unsigned(reg1099) : reg1098[(1'h0):(1'h0)]))) ?
                  (7'h42) : $unsigned($signed($unsigned(((8'hb8) - reg1100)))));
              reg1099 <= reg1101[(4'h9):(2'h3)];
            end
          else
            begin
              reg1098 <= $unsigned(reg1098[(1'h1):(1'h1)]);
              reg1099 <= reg1100;
              reg1100 <= ($signed({$signed($unsigned(wire1087))}) ^~ $signed(((-(|wire1092)) ?
                  {(wire1089 ? (8'hb0) : wire1088)} : $signed((8'ha8)))));
              reg1101 <= $signed(reg1099[(1'h1):(1'h0)]);
            end
          if ({(+(-$unsigned(reg1100))), {wire1085[(2'h3):(1'h1)], reg1101}})
            begin
              reg1102 <= $signed(wire1085[(2'h2):(1'h1)]);
              reg1103 <= $signed($signed(reg1098[(2'h3):(2'h2)]));
            end
          else
            begin
              reg1102 <= (reg1103 ? reg1097 : {reg1097, wire1086});
              reg1103 <= $signed(({wire1089,
                      {{reg1102, reg1101}, (reg1095 ? wire1088 : wire1094)}} ?
                  $signed(reg1098[(4'h8):(2'h3)]) : $signed(({(8'ha7),
                      wire1089} & reg1103[(2'h3):(2'h2)]))));
            end
        end
      reg1104 <= (!wire1086);
    end
  assign wire1105 = (((($signed(wire1089) ?
                        reg1097[(2'h2):(1'h1)] : reg1104[(3'h4):(1'h1)]) && (!$signed(wire1094))) ^ (8'ha3)) >> {$signed($signed($signed(wire1085)))});
  always
    @(posedge clk) begin
      if ($signed((((~^(wire1085 ~^ (8'haf))) ?
              ((^(8'hb2)) || (reg1096 == reg1101)) : reg1098) ?
          reg1099[(1'h1):(1'h0)] : $unsigned(reg1099))))
        begin
          if (($signed({(^~wire1090)}) ? $unsigned(reg1100) : wire1092))
            begin
              reg1106 <= $signed(wire1091[(1'h1):(1'h1)]);
            end
          else
            begin
              reg1106 <= ((-wire1090) ?
                  wire1091[(1'h0):(1'h0)] : ($unsigned($unsigned((~|reg1100))) ?
                      (reg1102 ?
                          (~&$signed(wire1091)) : $signed($unsigned((8'hb8)))) : (~^{(wire1085 ^~ reg1096)})));
            end
        end
      else
        begin
          reg1106 <= ($signed(reg1098) ?
              $signed($signed(((reg1097 & reg1098) ?
                  (reg1100 ?
                      wire1089 : wire1093) : ((8'hb7) >> wire1088)))) : ({{wire1092,
                          (reg1098 ? reg1101 : reg1101)},
                      $unsigned($unsigned(reg1096))} ?
                  ($unsigned($unsigned(wire1091)) ^ $unsigned((reg1097 <= (8'hb2)))) : $signed(reg1102[(4'hf):(4'hc)])));
          reg1107 <= (-$signed(wire1088[(5'h10):(4'ha)]));
          reg1108 <= wire1085[(2'h3):(1'h0)];
        end
    end
  assign wire1109 = reg1097[(3'h4):(2'h3)];
  assign wire1110 = reg1107[(4'h9):(4'h9)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1221
#( parameter param1256 = ((((+(+(8'hb0))) ^~ {{(8'hb2), (8'haf)}}) << (~|(8'hb0))) ? (8'ha6) : (!(7'h41))) )
(y, clk, wire1225, wire1224, wire1223, wire1222);
  output wire [(32'h17a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire1225;
  input wire [(3'h5):(1'h0)] wire1224;
  input wire signed [(4'hd):(1'h0)] wire1223;
  input wire [(5'h14):(1'h0)] wire1222;
  wire [(5'h11):(1'h0)] wire1255;
  reg signed [(4'he):(1'h0)] reg1254 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1253 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1252 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1251 = (1'h0);
  reg [(4'hb):(1'h0)] reg1250 = (1'h0);
  reg [(4'hf):(1'h0)] reg1249 = (1'h0);
  reg [(5'h11):(1'h0)] reg1248 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1247 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1246 = (1'h0);
  wire [(3'h7):(1'h0)] wire1245;
  wire [(5'h11):(1'h0)] wire1244;
  wire signed [(4'hc):(1'h0)] wire1243;
  wire [(3'h6):(1'h0)] wire1242;
  wire [(5'h10):(1'h0)] wire1241;
  reg signed [(5'h10):(1'h0)] reg1240 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1239 = (1'h0);
  reg [(5'h11):(1'h0)] reg1238 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1237 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1236 = (1'h0);
  reg [(2'h2):(1'h0)] reg1235 = (1'h0);
  reg [(4'hd):(1'h0)] reg1234 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1233 = (1'h0);
  reg [(4'h8):(1'h0)] reg1232 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1231 = (1'h0);
  reg [(5'h13):(1'h0)] reg1230 = (1'h0);
  wire [(5'h11):(1'h0)] wire1229;
  wire signed [(2'h3):(1'h0)] wire1228;
  wire signed [(4'hb):(1'h0)] wire1227;
  wire [(5'h10):(1'h0)] wire1226;
  assign y = {wire1255,
                 reg1254,
                 reg1253,
                 reg1252,
                 reg1251,
                 reg1250,
                 reg1249,
                 reg1248,
                 reg1247,
                 reg1246,
                 wire1245,
                 wire1244,
                 wire1243,
                 wire1242,
                 wire1241,
                 reg1240,
                 reg1239,
                 reg1238,
                 reg1237,
                 reg1236,
                 reg1235,
                 reg1234,
                 reg1233,
                 reg1232,
                 reg1231,
                 reg1230,
                 wire1229,
                 wire1228,
                 wire1227,
                 wire1226,
                 (1'h0)};
  assign wire1226 = (wire1224[(2'h3):(2'h3)] ?
                        (~&wire1223[(4'hc):(4'h9)]) : wire1223);
  assign wire1227 = (~&$unsigned(wire1222));
  assign wire1228 = ($signed(((wire1222[(4'ha):(3'h7)] ?
                                wire1222[(3'h6):(3'h6)] : $unsigned(wire1227)) ?
                            (~|$unsigned(wire1224)) : $unsigned({wire1227,
                                wire1222}))) ?
                        {(((wire1226 < wire1222) ?
                                (+wire1223) : wire1224) - (~|$signed(wire1227))),
                            $signed(wire1226[(1'h1):(1'h1)])} : (wire1224 ?
                            (!wire1225) : (((wire1223 ? wire1223 : wire1225) ?
                                wire1224[(2'h3):(1'h0)] : wire1223[(3'h5):(1'h1)]) << {$unsigned(wire1223),
                                wire1222})));
  assign wire1229 = $unsigned(wire1223);
  always
    @(posedge clk) begin
      if ($unsigned($signed((~&({wire1224} ?
          (wire1227 ? wire1225 : wire1229) : (wire1228 >= (8'hae)))))))
        begin
          reg1230 <= wire1228;
          reg1231 <= wire1227[(4'hb):(3'h5)];
          if ($signed(({wire1227,
              (wire1227 * $signed(wire1227))} + wire1224[(3'h4):(2'h2)])))
            begin
              reg1232 <= (8'hb5);
              reg1233 <= $signed($unsigned(($unsigned((reg1232 ?
                      reg1231 : wire1228)) ?
                  $signed(wire1225) : $unsigned(wire1223[(1'h1):(1'h1)]))));
              reg1234 <= reg1230;
              reg1235 <= ((~|wire1223[(4'ha):(4'ha)]) ?
                  $unsigned($signed((^(|wire1224)))) : $unsigned($unsigned(reg1232[(1'h1):(1'h1)])));
              reg1236 <= $signed(($signed($signed({reg1230})) ?
                  wire1226[(3'h5):(2'h2)] : ((8'hb7) ?
                      wire1222[(3'h4):(2'h2)] : $signed({(8'ha9), wire1229}))));
            end
          else
            begin
              reg1232 <= $unsigned($unsigned($unsigned(reg1236)));
              reg1233 <= (~|$signed(wire1228));
              reg1234 <= $unsigned((~^reg1235));
            end
        end
      else
        begin
          if ($unsigned((reg1231[(3'h4):(2'h3)] ?
              {($unsigned((8'h9d)) ?
                      (wire1227 ? wire1225 : reg1236) : {reg1231}),
                  reg1233} : ($unsigned($signed(wire1225)) >> ((^~reg1230) ?
                  {reg1235} : (|wire1227))))))
            begin
              reg1230 <= ($unsigned((~^$signed((reg1230 ?
                  reg1234 : wire1228)))) == (^reg1230));
              reg1231 <= $unsigned((~&(&{$unsigned(wire1222)})));
              reg1232 <= ($unsigned(wire1222) ?
                  (reg1233[(5'h13):(4'h8)] || $signed((wire1229[(4'hf):(3'h5)] >= (wire1225 ?
                      reg1233 : reg1230)))) : $unsigned($unsigned(wire1223)));
              reg1233 <= (((wire1227 ?
                      (^~$unsigned((8'hbd))) : $signed({(8'hb9), wire1222})) ?
                  (wire1227[(1'h1):(1'h0)] ?
                      ($unsigned(wire1228) ?
                          (wire1227 & reg1236) : (reg1236 ?
                              (8'h9c) : wire1229)) : $unsigned($unsigned(reg1230))) : (8'hbd)) * ($signed((((8'ha9) <<< reg1235) ?
                      $unsigned(wire1224) : (reg1233 > reg1231))) ?
                  {reg1232} : reg1232));
            end
          else
            begin
              reg1230 <= wire1227[(3'h7):(2'h3)];
              reg1231 <= reg1230[(4'hc):(2'h3)];
              reg1232 <= (wire1225[(1'h0):(1'h0)] <<< (wire1225 * ($signed($unsigned(reg1230)) < (~(wire1227 ?
                  wire1226 : wire1228)))));
            end
          reg1234 <= reg1232;
          reg1235 <= ((($unsigned({(8'hb9), reg1230}) ?
              (7'h44) : (reg1235[(1'h0):(1'h0)] ?
                  $signed(wire1228) : $signed(wire1225))) < (^~(!reg1234))) >> ($signed(($unsigned(reg1230) ?
              reg1235[(2'h2):(1'h1)] : wire1227)) >> $signed(($signed(reg1231) < $signed(reg1233)))));
        end
      reg1237 <= $signed((reg1233 ?
          (8'hae) : $unsigned($unsigned({reg1233, (8'hb1)}))));
      reg1238 <= (^(7'h43));
      reg1239 <= ((&$unsigned((wire1224 + reg1230))) | (wire1222[(5'h13):(3'h7)] ?
          ({((8'ha1) <<< wire1227), ((8'h9c) ? reg1233 : wire1227)} ?
              ((!reg1237) & $unsigned((8'h9c))) : {(reg1230 ?
                      wire1224 : wire1223)}) : reg1232));
      reg1240 <= ($signed($unsigned(reg1235)) != (+$signed($unsigned(reg1235))));
    end
  assign wire1241 = wire1222;
  assign wire1242 = (|(((!(wire1225 ? (8'h9f) : reg1235)) ?
                            $unsigned(wire1226[(1'h0):(1'h0)]) : reg1234[(4'ha):(3'h5)]) ?
                        {(!$unsigned(reg1232)),
                            $signed($signed(reg1238))} : reg1235[(1'h0):(1'h0)]));
  assign wire1243 = {((+($unsigned(reg1233) <= $unsigned(reg1231))) ?
                            (~$unsigned((reg1231 ?
                                wire1225 : wire1222))) : $signed($unsigned((^wire1228))))};
  assign wire1244 = (wire1222[(4'ha):(1'h0)] || wire1227);
  assign wire1245 = ($unsigned(wire1224[(1'h1):(1'h1)]) ?
                        ({wire1224[(2'h3):(1'h0)],
                            {reg1235, (~(8'had))}} > {reg1231[(3'h7):(3'h7)],
                            reg1236[(5'h12):(5'h12)]}) : (~&(|wire1228[(2'h2):(1'h0)])));
  always
    @(posedge clk) begin
      if ((~^(($unsigned((~reg1233)) ?
          $unsigned($unsigned(reg1236)) : $unsigned(wire1223[(1'h1):(1'h1)])) || (~&(8'hb4)))))
        begin
          reg1246 <= (~^({reg1238} ?
              (wire1242[(3'h5):(1'h1)] ^ {(wire1243 ?
                      wire1229 : reg1235)}) : reg1232));
          if (wire1229)
            begin
              reg1247 <= {wire1242[(1'h1):(1'h1)]};
            end
          else
            begin
              reg1247 <= $unsigned((~^$unsigned(wire1241)));
              reg1248 <= (wire1223[(1'h1):(1'h1)] ?
                  ({reg1230} ?
                      reg1234 : (($signed((8'hbf)) ?
                          $unsigned(reg1232) : (!reg1233)) == $unsigned(reg1247[(2'h2):(2'h2)]))) : wire1242[(1'h1):(1'h1)]);
            end
          if (wire1227[(3'h7):(1'h1)])
            begin
              reg1249 <= (wire1224[(1'h0):(1'h0)] ?
                  $unsigned(wire1241[(4'hc):(2'h3)]) : ({((+reg1233) ?
                          reg1231[(2'h3):(1'h0)] : (wire1242 ?
                              wire1241 : wire1241)),
                      ((reg1234 <<< wire1222) >>> (wire1244 + reg1237))} - (~^$unsigned(wire1227))));
              reg1250 <= $signed(((+($unsigned((7'h41)) != (8'hb4))) ?
                  $signed((!(reg1233 * wire1243))) : reg1236));
              reg1251 <= $unsigned(($signed((7'h43)) != $signed(wire1226)));
            end
          else
            begin
              reg1249 <= (reg1248 != $unsigned(wire1226));
              reg1250 <= wire1229;
              reg1251 <= reg1234;
              reg1252 <= reg1248;
            end
          reg1253 <= $unsigned($unsigned(reg1249[(2'h3):(1'h1)]));
        end
      else
        begin
          reg1246 <= $signed((reg1251 ^~ (^~$signed((reg1249 ?
              reg1232 : (8'had))))));
          reg1247 <= reg1238[(3'h7):(3'h7)];
          reg1248 <= ((~&$unsigned($signed(wire1242))) ?
              (reg1250[(4'h9):(3'h4)] ?
                  wire1222[(4'h9):(2'h3)] : wire1242) : (^$unsigned($unsigned(wire1224))));
          reg1249 <= (wire1223 + (wire1223[(3'h6):(2'h2)] != reg1233[(2'h2):(1'h0)]));
          if (reg1248)
            begin
              reg1250 <= (+((reg1232[(2'h2):(1'h0)] - $unsigned(wire1227)) >>> $unsigned(reg1235)));
              reg1251 <= wire1242;
            end
          else
            begin
              reg1250 <= (|(+reg1252[(3'h7):(2'h3)]));
            end
        end
      reg1254 <= ($unsigned((~|$unsigned($signed(wire1245)))) * wire1241[(1'h1):(1'h0)]);
    end
  assign wire1255 = reg1240;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1162  (y, clk, wire1166, wire1165, wire1164, wire1163);
  output wire [(32'h22a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire1166;
  input wire [(3'h6):(1'h0)] wire1165;
  input wire [(5'h13):(1'h0)] wire1164;
  input wire signed [(4'hc):(1'h0)] wire1163;
  wire [(2'h2):(1'h0)] wire1214;
  wire signed [(5'h10):(1'h0)] wire1213;
  wire [(4'h8):(1'h0)] wire1212;
  reg [(3'h4):(1'h0)] reg1211 = (1'h0);
  reg [(3'h6):(1'h0)] reg1210 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1209 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1208 = (1'h0);
  reg [(5'h11):(1'h0)] reg1207 = (1'h0);
  reg [(4'h8):(1'h0)] reg1206 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1205 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1204 = (1'h0);
  reg [(4'h8):(1'h0)] reg1203 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1202 = (1'h0);
  reg [(3'h6):(1'h0)] reg1201 = (1'h0);
  reg [(2'h2):(1'h0)] reg1200 = (1'h0);
  reg [(5'h12):(1'h0)] reg1199 = (1'h0);
  reg [(5'h14):(1'h0)] reg1198 = (1'h0);
  reg [(5'h13):(1'h0)] reg1197 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1196 = (1'h0);
  reg [(2'h2):(1'h0)] reg1195 = (1'h0);
  reg [(5'h10):(1'h0)] reg1194 = (1'h0);
  reg [(4'hc):(1'h0)] reg1193 = (1'h0);
  reg [(5'h12):(1'h0)] reg1192 = (1'h0);
  reg [(3'h4):(1'h0)] reg1191 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1190 = (1'h0);
  reg [(4'hc):(1'h0)] reg1189 = (1'h0);
  reg [(4'ha):(1'h0)] reg1188 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire1187;
  wire [(5'h13):(1'h0)] wire1186;
  wire [(3'h4):(1'h0)] wire1185;
  reg [(4'h8):(1'h0)] reg1184 = (1'h0);
  reg [(4'hc):(1'h0)] reg1183 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1182 = (1'h0);
  reg [(4'h8):(1'h0)] reg1181 = (1'h0);
  reg [(5'h11):(1'h0)] reg1180 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1179 = (1'h0);
  reg [(4'hc):(1'h0)] reg1178 = (1'h0);
  reg [(5'h13):(1'h0)] reg1177 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1176 = (1'h0);
  reg [(5'h13):(1'h0)] reg1175 = (1'h0);
  reg [(5'h15):(1'h0)] reg1174 = (1'h0);
  reg [(4'h9):(1'h0)] reg1173 = (1'h0);
  reg [(5'h15):(1'h0)] reg1172 = (1'h0);
  wire [(3'h6):(1'h0)] wire1171;
  wire [(5'h10):(1'h0)] wire1170;
  wire [(5'h12):(1'h0)] wire1169;
  wire signed [(3'h6):(1'h0)] wire1168;
  wire signed [(5'h14):(1'h0)] wire1167;
  assign y = {wire1214,
                 wire1213,
                 wire1212,
                 reg1211,
                 reg1210,
                 reg1209,
                 reg1208,
                 reg1207,
                 reg1206,
                 reg1205,
                 reg1204,
                 reg1203,
                 reg1202,
                 reg1201,
                 reg1200,
                 reg1199,
                 reg1198,
                 reg1197,
                 reg1196,
                 reg1195,
                 reg1194,
                 reg1193,
                 reg1192,
                 reg1191,
                 reg1190,
                 reg1189,
                 reg1188,
                 wire1187,
                 wire1186,
                 wire1185,
                 reg1184,
                 reg1183,
                 reg1182,
                 reg1181,
                 reg1180,
                 reg1179,
                 reg1178,
                 reg1177,
                 reg1176,
                 reg1175,
                 reg1174,
                 reg1173,
                 reg1172,
                 wire1171,
                 wire1170,
                 wire1169,
                 wire1168,
                 wire1167,
                 (1'h0)};
  assign wire1167 = wire1164;
  assign wire1168 = (wire1165[(1'h1):(1'h0)] == (!wire1164[(4'hc):(1'h0)]));
  assign wire1169 = ($signed($signed($unsigned(wire1165[(3'h5):(3'h5)]))) > ($signed(wire1164[(4'hb):(4'h8)]) ^~ wire1168[(2'h2):(2'h2)]));
  assign wire1170 = ((8'hb6) ?
                        {(|($signed((8'hb9)) || (wire1166 != wire1164))),
                            wire1165} : $signed((^~wire1168[(2'h2):(2'h2)])));
  assign wire1171 = ((wire1165[(1'h1):(1'h0)] && (($unsigned(wire1165) && $signed(wire1165)) >> $unsigned(wire1170))) << $unsigned(((^(8'hb4)) & $signed((|wire1163)))));
  always
    @(posedge clk) begin
      reg1172 <= (+wire1169);
      if (($signed(({$unsigned(wire1170)} ?
          wire1167 : $signed((^~wire1169)))) ^~ (8'ha1)))
        begin
          reg1173 <= $unsigned(wire1164[(4'h9):(1'h1)]);
          if (wire1165)
            begin
              reg1174 <= ((wire1165 ?
                  (!$unsigned(reg1172[(4'h9):(3'h6)])) : wire1163) + $unsigned((wire1165 ?
                  ($unsigned((8'hb7)) <<< $signed(wire1168)) : (+(wire1169 ?
                      reg1173 : wire1163)))));
              reg1175 <= (!{$unsigned(((^~wire1169) ?
                      wire1167[(1'h0):(1'h0)] : $signed(wire1165))),
                  (wire1166 ?
                      $signed(((8'ha7) ~^ reg1172)) : $unsigned((!reg1173)))});
              reg1176 <= $signed(wire1166);
              reg1177 <= (~|($unsigned(wire1163) > $unsigned(wire1168[(3'h5):(3'h5)])));
              reg1178 <= $signed({wire1164});
            end
          else
            begin
              reg1174 <= (~((reg1176[(4'hc):(1'h0)] ?
                      (wire1171 >= reg1173) : $unsigned((^wire1165))) ?
                  ($signed($unsigned(wire1170)) ?
                      (wire1170[(1'h1):(1'h0)] ^~ $signed(wire1165)) : reg1172[(3'h5):(3'h4)]) : wire1166[(2'h3):(1'h1)]));
            end
          reg1179 <= (8'hbf);
        end
      else
        begin
          reg1173 <= wire1171;
          reg1174 <= reg1173;
          reg1175 <= (((wire1163 * reg1176) ?
                  (^{wire1164[(2'h3):(1'h0)],
                      $signed(wire1169)}) : ($signed((reg1179 ?
                          (8'ha0) : reg1178)) ?
                      (-reg1174) : ($unsigned((8'hbd)) ?
                          ((8'ha8) ?
                              wire1170 : wire1170) : wire1166[(4'h8):(3'h6)]))) ?
              wire1163 : (wire1171 ?
                  (wire1163 < (~^(8'hbc))) : (^~{(&reg1176),
                      $signed(wire1167)})));
          reg1176 <= $unsigned(reg1177);
          if ({{($unsigned($unsigned(reg1175)) == $signed(wire1167[(5'h14):(5'h14)]))}})
            begin
              reg1177 <= (($signed(({(8'ha9)} <= ((8'hb0) - wire1163))) != ($unsigned($signed((8'ha0))) << wire1171[(3'h6):(2'h3)])) ?
                  {$unsigned($signed($unsigned(wire1163)))} : reg1173);
              reg1178 <= $signed($unsigned(reg1176));
              reg1179 <= (reg1175 < wire1170);
              reg1180 <= $signed(((reg1177 ?
                  ({reg1174} ?
                      reg1175[(3'h7):(2'h2)] : (8'hac)) : $unsigned($signed(wire1169))) ~^ (~&(7'h41))));
            end
          else
            begin
              reg1177 <= (~|{(+($unsigned(wire1164) >>> wire1171))});
              reg1178 <= ((~|$unsigned((reg1172 ?
                  reg1176[(4'hf):(1'h1)] : wire1168))) >= ((wire1170 ?
                      reg1177[(4'hf):(4'he)] : {(~|(8'h9e)),
                          reg1180[(4'hf):(4'he)]}) ?
                  {(^$signed(reg1172)),
                      (((8'hbd) >>> wire1163) ?
                          (wire1171 >= (8'hb7)) : $unsigned(wire1163))} : wire1171));
              reg1179 <= ($unsigned(wire1163) ?
                  ({(reg1178[(3'h7):(2'h3)] & $unsigned((8'hb0)))} <= $signed(((wire1169 ^~ reg1180) >>> reg1180))) : $unsigned((8'ha2)));
              reg1180 <= (|reg1177);
              reg1181 <= (~&(~|$unsigned({(~|wire1164),
                  (reg1176 ? reg1180 : reg1175)})));
            end
        end
      if ((|reg1174[(5'h12):(4'hb)]))
        begin
          reg1182 <= {($unsigned(($unsigned(reg1173) ?
                  wire1168[(1'h0):(1'h0)] : wire1164[(3'h7):(2'h3)])) & (7'h42))};
        end
      else
        begin
          reg1182 <= ((reg1172[(5'h13):(4'h8)] ? reg1180 : reg1173) ?
              reg1176 : ($signed(reg1180) ^~ $signed($signed(wire1168[(1'h0):(1'h0)]))));
          reg1183 <= $signed($unsigned({reg1172[(2'h2):(1'h0)],
              ((wire1168 ? wire1170 : reg1177) ?
                  $signed(wire1164) : (~reg1176))}));
          reg1184 <= $signed((|{$signed((wire1171 <<< wire1170)), reg1181}));
        end
    end
  assign wire1185 = (&wire1169[(1'h1):(1'h1)]);
  assign wire1186 = $signed(reg1181);
  assign wire1187 = (8'ha0);
  always
    @(posedge clk) begin
      reg1188 <= (8'hb9);
      if ((reg1176 ?
          wire1164[(5'h12):(3'h4)] : $signed($unsigned(wire1163[(1'h1):(1'h1)]))))
        begin
          reg1189 <= (reg1182 <<< $unsigned((({wire1186, reg1174} ?
                  (~reg1178) : $signed(wire1168)) ?
              $signed(wire1164[(5'h10):(2'h2)]) : $unsigned((reg1182 || reg1179)))));
          if ((((wire1167 ?
                      (&wire1166) : {reg1181[(3'h5):(2'h2)],
                          (wire1170 ? wire1163 : wire1165)}) ?
                  $unsigned((~^(~|reg1184))) : reg1174[(4'hd):(3'h6)]) ?
              $unsigned($signed((wire1169[(3'h4):(2'h3)] ?
                  $unsigned(wire1169) : $signed(wire1171)))) : (-reg1175[(1'h0):(1'h0)])))
            begin
              reg1190 <= $unsigned({($signed($unsigned(wire1187)) == wire1185),
                  (8'ha2)});
              reg1191 <= (7'h44);
            end
          else
            begin
              reg1190 <= $signed(reg1182[(3'h4):(3'h4)]);
            end
          if (reg1178)
            begin
              reg1192 <= reg1189[(3'h6):(1'h0)];
              reg1193 <= (|{((reg1173[(4'h8):(2'h2)] ?
                          {reg1182, reg1184} : $signed(reg1189)) ?
                      $signed(reg1181) : reg1180[(4'he):(4'hb)])});
            end
          else
            begin
              reg1192 <= {(~wire1185), wire1167[(2'h3):(1'h0)]};
            end
          if ((+(|wire1168[(3'h6):(1'h0)])))
            begin
              reg1194 <= {(($unsigned(reg1175) ?
                      (-$unsigned(reg1189)) : (8'haf)) || $signed({(reg1178 ?
                          wire1170 : wire1171),
                      (wire1166 ? wire1164 : wire1164)})),
                  {{wire1187, reg1177}}};
              reg1195 <= {{$signed(((|wire1171) ?
                          $signed(wire1186) : wire1171[(3'h6):(3'h6)])),
                      reg1177}};
            end
          else
            begin
              reg1194 <= $signed((wire1163[(1'h0):(1'h0)] ?
                  reg1193 : wire1171));
              reg1195 <= wire1167;
              reg1196 <= {(((|wire1169) ? reg1182 : (8'had)) || (8'hb7)),
                  $signed($unsigned(reg1176[(4'h8):(1'h0)]))};
              reg1197 <= (^~$unsigned((!(8'hb1))));
            end
          reg1198 <= wire1167;
        end
      else
        begin
          reg1189 <= ((!(+{$signed(reg1178)})) <= $signed(((^~{wire1164}) ?
              wire1168[(2'h2):(2'h2)] : {(|wire1187)})));
          if (($unsigned((8'hb2)) ?
              $signed((~^(~&reg1177[(1'h0):(1'h0)]))) : reg1181))
            begin
              reg1190 <= wire1185[(1'h1):(1'h0)];
            end
          else
            begin
              reg1190 <= (~|$unsigned(wire1167[(3'h4):(1'h0)]));
              reg1191 <= (reg1183 || $unsigned($unsigned(($signed(reg1178) >= $signed(wire1169)))));
              reg1192 <= reg1197;
              reg1193 <= $unsigned(reg1194);
              reg1194 <= $unsigned(wire1166);
            end
        end
      if (({(|reg1194)} ? (8'haf) : reg1174))
        begin
          reg1199 <= $unsigned($signed($signed(((|wire1169) & {reg1173,
              (8'hb3)}))));
          reg1200 <= $unsigned(reg1194[(4'ha):(2'h3)]);
          if ($unsigned((~&$signed((reg1198 & $signed(wire1171))))))
            begin
              reg1201 <= $unsigned(reg1194);
              reg1202 <= (((((^~reg1198) ? (^(8'h9d)) : {wire1163}) ?
                      (!(reg1192 > reg1195)) : ($signed(wire1167) < (reg1173 | wire1185))) ?
                  $unsigned(wire1169) : $signed(reg1198[(5'h13):(2'h2)])) == ({(-$unsigned(reg1180)),
                      $signed((reg1199 != wire1166))} ?
                  (reg1182[(2'h3):(2'h2)] ?
                      ((^~wire1166) ?
                          reg1198[(2'h2):(2'h2)] : {wire1186}) : {reg1195[(1'h0):(1'h0)]}) : (|(~reg1197))));
              reg1203 <= $signed((~&$signed(reg1172)));
            end
          else
            begin
              reg1201 <= (^~(reg1191 >>> (wire1167 ^~ reg1197)));
              reg1202 <= reg1184;
              reg1203 <= ($unsigned({reg1198[(2'h3):(2'h3)]}) ^~ $unsigned(reg1200));
            end
          reg1204 <= $unsigned((|$signed(reg1179[(3'h4):(1'h1)])));
          reg1205 <= $unsigned(reg1189[(4'hb):(4'h9)]);
        end
      else
        begin
          if ({(-reg1182[(4'he):(4'h9)]), (~reg1199[(3'h7):(2'h3)])})
            begin
              reg1199 <= ((7'h40) <<< ($signed($signed($signed(reg1173))) - ({$signed(wire1185)} * reg1180)));
            end
          else
            begin
              reg1199 <= {$unsigned(wire1169), (~|wire1166)};
              reg1200 <= (reg1179 ?
                  ({{{reg1190}, $unsigned(wire1168)}} ?
                      ({wire1187} ?
                          $signed((reg1196 ?
                              reg1176 : reg1175)) : ($unsigned(reg1179) ?
                              $unsigned(reg1175) : $unsigned(reg1191))) : reg1194) : $signed((~^((reg1182 ?
                          reg1205 : reg1194) ?
                      (reg1172 >= reg1204) : {reg1177}))));
              reg1201 <= (8'hb5);
            end
          if ((reg1192[(4'hf):(3'h5)] ?
              reg1182[(3'h4):(2'h3)] : reg1193[(4'hc):(1'h0)]))
            begin
              reg1202 <= ($signed(reg1184[(3'h6):(1'h1)]) > ($signed(reg1190) - (({wire1168,
                          reg1173} ?
                      $signed((7'h44)) : (~^(8'hb9))) ?
                  $unsigned((wire1164 ? (8'hbc) : reg1188)) : {(8'h9d),
                      wire1164[(4'hb):(1'h1)]})));
              reg1203 <= reg1184[(3'h4):(3'h4)];
              reg1204 <= (wire1170[(2'h2):(1'h1)] ^ ((-(~^$signed(wire1166))) ?
                  ((-((8'haf) ? wire1170 : reg1201)) ?
                      {reg1193,
                          (~^reg1199)} : (reg1188 ^ reg1181)) : (((~|reg1196) ?
                      $unsigned(reg1184) : (wire1186 ?
                          wire1168 : (8'ha4))) >= ($signed(reg1177) * (reg1194 ?
                      reg1205 : wire1187)))));
              reg1205 <= ((~|$signed(wire1165)) <= reg1188);
              reg1206 <= (wire1167 ?
                  (reg1197 ? reg1176 : wire1167) : reg1191[(2'h3):(1'h1)]);
            end
          else
            begin
              reg1202 <= wire1185[(1'h1):(1'h0)];
              reg1203 <= $unsigned(reg1203[(3'h5):(1'h0)]);
            end
          reg1207 <= reg1204[(3'h5):(2'h3)];
          reg1208 <= wire1165;
          reg1209 <= (~reg1176);
        end
      reg1210 <= (~reg1197);
      reg1211 <= reg1176[(3'h7):(1'h0)];
    end
  assign wire1212 = ((reg1177[(4'ha):(3'h7)] ?
                            (($signed(reg1177) || reg1180) & $signed(reg1203[(3'h6):(3'h6)])) : (|(+wire1163))) ?
                        $signed($unsigned((~reg1178))) : $signed({$signed((reg1210 ?
                                (8'hb3) : reg1198)),
                            ((^~reg1211) * $unsigned(reg1193))}));
  assign wire1213 = ($unsigned(($unsigned((|reg1206)) ?
                            ((~&reg1199) ?
                                (wire1212 ?
                                    reg1188 : reg1211) : (reg1176 && (8'ha8))) : wire1164)) ?
                        reg1188[(4'h8):(3'h4)] : wire1165[(1'h1):(1'h0)]);
  assign wire1214 = (wire1166 ?
                        ((^~$unsigned(((8'hb2) ? (8'hb2) : reg1199))) ?
                            $unsigned(((reg1179 >>> reg1193) >>> (reg1204 != wire1168))) : (+$signed((^~(8'ha7))))) : $unsigned($signed(($unsigned(wire1167) ?
                            wire1168 : (~&wire1169)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1580  (y, clk, wire1585, wire1584, wire1583, wire1582, wire1581);
  output wire [(32'h26f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire1585;
  input wire [(2'h2):(1'h0)] wire1584;
  input wire signed [(4'hd):(1'h0)] wire1583;
  input wire signed [(4'hf):(1'h0)] wire1582;
  input wire signed [(5'h15):(1'h0)] wire1581;
  reg signed [(4'hf):(1'h0)] reg1637 = (1'h0);
  reg [(4'hc):(1'h0)] reg1636 = (1'h0);
  reg [(3'h6):(1'h0)] reg1635 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1634 = (1'h0);
  reg [(4'hb):(1'h0)] reg1633 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1632 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1631 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1630 = (1'h0);
  reg [(4'h9):(1'h0)] reg1629 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1628 = (1'h0);
  reg [(4'hc):(1'h0)] reg1627 = (1'h0);
  reg [(3'h7):(1'h0)] reg1626 = (1'h0);
  reg [(5'h14):(1'h0)] reg1625 = (1'h0);
  reg [(2'h3):(1'h0)] reg1624 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1623 = (1'h0);
  reg [(4'hb):(1'h0)] reg1622 = (1'h0);
  wire [(5'h14):(1'h0)] wire1621;
  wire [(4'h8):(1'h0)] wire1620;
  wire signed [(4'hc):(1'h0)] wire1619;
  wire [(3'h5):(1'h0)] wire1618;
  wire signed [(5'h13):(1'h0)] wire1617;
  reg signed [(4'ha):(1'h0)] reg1616 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1615 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1614 = (1'h0);
  reg [(4'he):(1'h0)] reg1613 = (1'h0);
  reg [(5'h10):(1'h0)] reg1612 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1611 = (1'h0);
  reg [(3'h5):(1'h0)] reg1610 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1609 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1608 = (1'h0);
  reg [(5'h13):(1'h0)] reg1607 = (1'h0);
  reg [(3'h7):(1'h0)] reg1606 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1605 = (1'h0);
  reg [(4'hb):(1'h0)] reg1604 = (1'h0);
  reg [(3'h5):(1'h0)] reg1603 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1602 = (1'h0);
  reg [(4'hb):(1'h0)] reg1601 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1600 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1599 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1598 = (1'h0);
  reg [(3'h6):(1'h0)] reg1597 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1596;
  wire [(5'h15):(1'h0)] wire1595;
  wire signed [(4'ha):(1'h0)] wire1594;
  wire [(4'hc):(1'h0)] wire1593;
  wire signed [(2'h2):(1'h0)] wire1592;
  wire signed [(4'he):(1'h0)] wire1591;
  wire signed [(4'he):(1'h0)] wire1590;
  wire signed [(5'h15):(1'h0)] wire1589;
  wire [(4'hd):(1'h0)] wire1588;
  wire [(4'he):(1'h0)] wire1587;
  wire signed [(5'h15):(1'h0)] wire1586;
  assign y = {reg1637,
                 reg1636,
                 reg1635,
                 reg1634,
                 reg1633,
                 reg1632,
                 reg1631,
                 reg1630,
                 reg1629,
                 reg1628,
                 reg1627,
                 reg1626,
                 reg1625,
                 reg1624,
                 reg1623,
                 reg1622,
                 wire1621,
                 wire1620,
                 wire1619,
                 wire1618,
                 wire1617,
                 reg1616,
                 reg1615,
                 reg1614,
                 reg1613,
                 reg1612,
                 reg1611,
                 reg1610,
                 reg1609,
                 reg1608,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1604,
                 reg1603,
                 reg1602,
                 reg1601,
                 reg1600,
                 reg1599,
                 reg1598,
                 reg1597,
                 wire1596,
                 wire1595,
                 wire1594,
                 wire1593,
                 wire1592,
                 wire1591,
                 wire1590,
                 wire1589,
                 wire1588,
                 wire1587,
                 wire1586,
                 (1'h0)};
  assign wire1586 = $unsigned($signed(((wire1581 & $signed(wire1583)) ?
                        (wire1583[(2'h3):(2'h2)] < ((8'hb7) ?
                            wire1584 : wire1582)) : $signed((|wire1584)))));
  assign wire1587 = {(($signed($unsigned(wire1583)) << wire1585[(2'h2):(1'h1)]) ?
                            (8'hab) : (~|{wire1585[(1'h1):(1'h0)],
                                (wire1584 >>> wire1584)}))};
  assign wire1588 = $unsigned(wire1583);
  assign wire1589 = wire1588[(1'h0):(1'h0)];
  assign wire1590 = wire1581[(4'ha):(3'h4)];
  assign wire1591 = {{(^~(wire1589 > (~&wire1582))),
                            ((+(!wire1587)) >>> wire1584)}};
  assign wire1592 = (wire1583[(1'h0):(1'h0)] ^ $signed((wire1582[(1'h0):(1'h0)] << wire1586)));
  assign wire1593 = (wire1583[(2'h3):(1'h0)] >> (~|$unsigned(((wire1587 ?
                        wire1588 : wire1581) || wire1581))));
  assign wire1594 = (~^$signed($signed($unsigned(wire1593))));
  assign wire1595 = wire1587;
  assign wire1596 = ($unsigned(wire1591[(4'ha):(4'h9)]) ?
                        wire1590[(3'h6):(2'h3)] : $unsigned((~^{$unsigned(wire1595),
                            wire1588[(2'h3):(2'h2)]})));
  always
    @(posedge clk) begin
      if (wire1590[(4'hd):(3'h4)])
        begin
          if ({$unsigned((+wire1593)),
              $unsigned((($unsigned(wire1592) ? $signed(wire1594) : wire1595) ?
                  $signed(wire1584[(1'h0):(1'h0)]) : (wire1589[(4'hc):(4'h9)] ^ wire1581)))})
            begin
              reg1597 <= $unsigned($signed(wire1583));
              reg1598 <= ($signed(({wire1591,
                      (reg1597 | wire1588)} & (((8'ha3) | wire1591) ?
                      wire1592[(2'h2):(2'h2)] : $signed((8'ha7))))) ?
                  ($signed($unsigned($unsigned(wire1591))) >> wire1582[(4'hf):(2'h2)]) : $signed((reg1597 ?
                      (~&(wire1596 ?
                          wire1585 : wire1592)) : ($unsigned((8'hb3)) << wire1591[(4'h8):(3'h7)]))));
              reg1599 <= {$unsigned((-(^(wire1589 ~^ wire1594))))};
            end
          else
            begin
              reg1597 <= ((((~reg1597) + (wire1594[(3'h7):(3'h6)] != (^wire1582))) >>> $signed((8'hbd))) || (reg1599[(5'h13):(4'hd)] > (8'h9f)));
            end
          if ((($signed($unsigned((wire1593 | wire1587))) ?
              $signed(reg1597[(2'h3):(1'h1)]) : $signed(wire1581[(5'h13):(5'h12)])) ^~ ({(wire1593[(4'h9):(4'h8)] == (wire1582 ?
                  wire1581 : wire1593))} + $unsigned(($signed(wire1592) ~^ wire1583)))))
            begin
              reg1600 <= (&{wire1594[(3'h4):(1'h0)]});
            end
          else
            begin
              reg1600 <= wire1588;
              reg1601 <= $signed($unsigned((~&$unsigned((wire1583 >= wire1585)))));
              reg1602 <= $signed(wire1593);
            end
          reg1603 <= wire1591[(4'hd):(4'hb)];
          reg1604 <= wire1585[(2'h2):(2'h2)];
        end
      else
        begin
          reg1597 <= ($signed((((reg1597 << (8'hb0)) << (wire1595 && wire1589)) ?
              $signed(wire1586) : $signed({wire1583,
                  wire1583}))) * (($signed({reg1602}) == {wire1582[(1'h0):(1'h0)],
              wire1586[(4'h9):(2'h3)]}) | wire1593[(4'h8):(2'h2)]));
          if ((~^{wire1590}))
            begin
              reg1598 <= $signed(wire1581[(2'h2):(1'h0)]);
              reg1599 <= {$signed(($unsigned((reg1598 ?
                      wire1591 : wire1583)) | wire1586))};
              reg1600 <= ((~wire1587) ? wire1593[(1'h1):(1'h1)] : wire1581);
              reg1601 <= wire1588[(4'h9):(1'h0)];
              reg1602 <= wire1588[(4'h9):(3'h4)];
            end
          else
            begin
              reg1598 <= $signed(((($signed(reg1601) > (~^(8'ha7))) != reg1602) != {wire1589,
                  wire1585}));
              reg1599 <= (wire1583 * {$signed({(~wire1591)}),
                  reg1598[(2'h2):(1'h1)]});
              reg1600 <= ({$unsigned($unsigned((!wire1581)))} ?
                  wire1592[(2'h2):(1'h1)] : ($unsigned($unsigned((wire1591 >>> reg1602))) >> $signed({(wire1588 ?
                          wire1588 : wire1594)})));
              reg1601 <= $signed($unsigned(reg1603[(2'h2):(1'h1)]));
            end
          reg1603 <= $signed((8'ha4));
          if ($unsigned(reg1602[(3'h7):(3'h7)]))
            begin
              reg1604 <= (($unsigned((|(~^wire1593))) ^~ ((reg1599 && (~^wire1581)) <= reg1600)) ?
                  (^($unsigned(reg1597[(3'h4):(2'h2)]) ?
                      (^wire1585[(3'h4):(2'h2)]) : wire1593)) : (($unsigned((^wire1594)) <<< (wire1589 ?
                      $signed(wire1587) : $signed(reg1603))) > wire1594[(4'h9):(3'h4)]));
            end
          else
            begin
              reg1604 <= wire1584;
              reg1605 <= (wire1596[(3'h5):(2'h2)] < (-wire1595[(4'hc):(4'ha)]));
              reg1606 <= {$signed(($signed(wire1596[(1'h1):(1'h0)]) ?
                      wire1584[(2'h2):(2'h2)] : wire1582[(4'hc):(2'h2)])),
                  (((~^reg1605[(1'h1):(1'h1)]) ?
                      (!$signed(wire1593)) : wire1584[(2'h2):(1'h0)]) << $signed(wire1595))};
            end
        end
    end
  always
    @(posedge clk) begin
      if (wire1582[(3'h4):(3'h4)])
        begin
          if ({{(reg1603 ?
                      ($signed(reg1600) >>> reg1600[(4'h8):(3'h6)]) : $unsigned(wire1591)),
                  (wire1593[(3'h6):(3'h6)] ?
                      wire1595[(1'h0):(1'h0)] : wire1587[(3'h4):(2'h3)])},
              (&(wire1585[(4'h9):(1'h0)] || wire1583[(4'hc):(1'h1)]))})
            begin
              reg1607 <= wire1589;
              reg1608 <= (reg1605 ?
                  (^~((-(wire1590 + wire1591)) ?
                      ((^wire1588) >= $unsigned(reg1605)) : $unsigned($signed(wire1589)))) : $unsigned($signed({$unsigned(wire1590)})));
              reg1609 <= ({(reg1598[(3'h5):(2'h3)] ?
                      wire1588[(4'hd):(1'h1)] : ($signed(reg1605) - wire1593[(1'h0):(1'h0)])),
                  ((-(reg1602 ? wire1583 : wire1581)) ?
                      ($signed(reg1603) | $unsigned(reg1605)) : reg1598)} ~^ ($signed($unsigned(wire1590)) + ($unsigned($unsigned(wire1594)) ?
                  wire1591[(3'h4):(2'h2)] : (((8'ha4) | wire1584) + reg1607))));
            end
          else
            begin
              reg1607 <= (($signed(reg1598) ?
                      {wire1593[(1'h1):(1'h1)]} : ({{wire1595, (8'hac)}} ?
                          $unsigned((7'h43)) : ((wire1594 ?
                              reg1608 : (8'hb3)) <<< (reg1602 ?
                              (8'had) : reg1600)))) ?
                  {reg1598, reg1605} : $unsigned((&(8'hbc))));
              reg1608 <= wire1594[(1'h0):(1'h0)];
              reg1609 <= ((wire1595[(4'he):(4'h8)] ?
                      $signed(reg1598[(3'h4):(2'h2)]) : {(((8'hae) >>> reg1597) ?
                              $unsigned(wire1584) : wire1584[(2'h2):(1'h0)])}) ?
                  (^~reg1609) : ({$unsigned((+reg1597)),
                      (~&(|reg1603))} | $unsigned($signed(wire1595[(2'h2):(1'h1)]))));
              reg1610 <= wire1595[(1'h0):(1'h0)];
              reg1611 <= (8'h9e);
            end
          reg1612 <= $signed(wire1593);
          reg1613 <= reg1608;
          reg1614 <= (8'hba);
          reg1615 <= wire1588[(4'hb):(3'h4)];
        end
      else
        begin
          reg1607 <= wire1596;
        end
      reg1616 <= {$signed(wire1596[(3'h4):(2'h3)]), (8'hba)};
    end
  assign wire1617 = wire1581[(5'h12):(5'h12)];
  assign wire1618 = reg1600;
  assign wire1619 = (~|reg1608);
  assign wire1620 = $unsigned($signed(wire1588));
  assign wire1621 = ((wire1593[(4'hc):(3'h5)] ^ {wire1589[(4'h8):(3'h6)],
                            ((wire1620 ?
                                wire1587 : reg1614) || $signed(wire1586))}) ?
                        {$signed(wire1595[(2'h3):(1'h0)]),
                            $signed({$unsigned((8'ha4))})} : $unsigned(wire1583[(3'h7):(3'h6)]));
  always
    @(posedge clk) begin
      reg1622 <= wire1590;
      if ($signed($unsigned($signed((&(~&wire1596))))))
        begin
          reg1623 <= ($signed(reg1599[(1'h1):(1'h0)]) - $signed((&reg1603)));
          if (reg1616)
            begin
              reg1624 <= wire1584;
            end
          else
            begin
              reg1624 <= (~(($signed({wire1619}) ? (8'hb1) : wire1587) ?
                  $unsigned($unsigned(reg1599[(4'hd):(4'hd)])) : reg1600[(2'h3):(2'h3)]));
              reg1625 <= ((8'hbd) ?
                  (wire1621 ?
                      ($signed($signed(reg1598)) == $unsigned(wire1585[(2'h3):(2'h2)])) : (~|reg1614[(1'h0):(1'h0)])) : wire1583[(4'hb):(3'h5)]);
              reg1626 <= reg1605;
              reg1627 <= (~|$signed($signed(((reg1606 ? wire1590 : wire1586) ?
                  $unsigned(reg1607) : $signed(reg1623)))));
            end
        end
      else
        begin
          reg1623 <= ((&(^wire1584)) | $signed(reg1624));
          reg1624 <= $unsigned($signed($signed($unsigned(wire1588[(3'h4):(3'h4)]))));
          reg1625 <= {$signed((8'h9c))};
        end
      if ((!$unsigned(reg1616)))
        begin
          reg1628 <= reg1597[(2'h3):(1'h0)];
          if (reg1625[(4'ha):(3'h7)])
            begin
              reg1629 <= $unsigned($unsigned(($unsigned({reg1625,
                  (8'hb7)}) | $unsigned(reg1599[(4'hc):(1'h1)]))));
              reg1630 <= $signed($signed(reg1624[(2'h2):(2'h2)]));
              reg1631 <= {((reg1599[(4'h8):(4'h8)] ?
                      {(wire1593 ^~ reg1616)} : ($signed(reg1600) & (~^reg1610))) * (8'haf))};
              reg1632 <= (reg1598[(4'h9):(3'h6)] ?
                  $unsigned((reg1614 ?
                      {(wire1596 < reg1616)} : (-$signed(wire1583)))) : $signed($unsigned({(wire1588 ?
                          reg1597 : reg1613)})));
              reg1633 <= $unsigned({$unsigned((~&(wire1617 >> wire1596))),
                  (+((~^wire1585) & reg1629[(3'h6):(3'h6)]))});
            end
          else
            begin
              reg1629 <= (|{({(!reg1632), reg1612[(4'hd):(4'h9)]} + wire1583)});
              reg1630 <= (($unsigned(((&(7'h43)) && (reg1623 > reg1606))) ?
                      {(reg1630 >= {reg1603})} : $signed($signed(reg1607[(5'h12):(1'h1)]))) ?
                  reg1610[(1'h1):(1'h1)] : ((reg1615[(1'h1):(1'h0)] ?
                          wire1587[(3'h5):(3'h5)] : $signed($unsigned(wire1590))) ?
                      wire1594[(1'h0):(1'h0)] : reg1604[(4'ha):(3'h6)]));
              reg1631 <= {(((^~(reg1603 | reg1600)) ?
                      (!reg1607[(5'h13):(4'he)]) : reg1603[(2'h3):(2'h3)]) * wire1618),
                  wire1594};
              reg1632 <= reg1622[(3'h6):(2'h3)];
              reg1633 <= reg1599;
            end
          if (reg1628)
            begin
              reg1634 <= {(($unsigned((7'h43)) ?
                          $unsigned((^~reg1612)) : wire1620) ?
                      (((^reg1606) ? reg1602 : (wire1592 ? reg1612 : (8'h9d))) ?
                          (^$signed((8'h9d))) : reg1626) : {reg1616[(4'ha):(3'h6)],
                          $unsigned(wire1595[(5'h10):(3'h4)])})};
            end
          else
            begin
              reg1634 <= (8'hae);
            end
          reg1635 <= (^(wire1619 >>> ($unsigned({wire1617,
              wire1620}) ^~ ((wire1586 == reg1609) != reg1627[(1'h1):(1'h1)]))));
          reg1636 <= reg1609[(3'h6):(2'h2)];
        end
      else
        begin
          reg1628 <= reg1624;
        end
      if ((^~((($signed(wire1618) > (~(8'hb1))) ?
              (+(wire1585 ? reg1600 : reg1625)) : reg1636[(4'h8):(2'h3)]) ?
          (+reg1601[(3'h7):(3'h6)]) : reg1631[(4'he):(4'hc)])))
        begin
          reg1637 <= {reg1625};
        end
      else
        begin
          reg1637 <= $unsigned({$signed({$unsigned(wire1590),
                  $signed(reg1601)}),
              $unsigned(((~&wire1587) * {wire1587, reg1628}))});
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1545
#( parameter param1569 = ({(-{((8'hb4) ? (8'hb5) : (8'hb5)), (+(8'hb3))}), ((~&{(8'haf)}) ? {(~^(8'hb3))} : (((8'haf) < (8'had)) + {(8'hab), (7'h40)}))} ~^ {(8'h9f)}) )
(y, clk, wire1550, wire1549, wire1548, wire1547, wire1546);
  output wire [(32'hb8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire1550;
  input wire [(5'h10):(1'h0)] wire1549;
  input wire [(5'h11):(1'h0)] wire1548;
  input wire [(2'h2):(1'h0)] wire1547;
  input wire signed [(3'h4):(1'h0)] wire1546;
  wire [(2'h3):(1'h0)] wire1568;
  reg signed [(4'he):(1'h0)] reg1567 = (1'h0);
  reg [(4'he):(1'h0)] reg1566 = (1'h0);
  reg [(4'hb):(1'h0)] reg1565 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1564 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1563 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1562 = (1'h0);
  reg [(2'h2):(1'h0)] reg1561 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1560 = (1'h0);
  reg [(4'h9):(1'h0)] reg1559 = (1'h0);
  reg [(2'h2):(1'h0)] reg1558 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1557 = (1'h0);
  reg [(4'h8):(1'h0)] reg1556 = (1'h0);
  wire [(5'h12):(1'h0)] wire1555;
  wire signed [(5'h14):(1'h0)] wire1554;
  wire [(4'hc):(1'h0)] wire1553;
  wire signed [(2'h3):(1'h0)] wire1552;
  wire signed [(2'h2):(1'h0)] wire1551;
  assign y = {wire1568,
                 reg1567,
                 reg1566,
                 reg1565,
                 reg1564,
                 reg1563,
                 reg1562,
                 reg1561,
                 reg1560,
                 reg1559,
                 reg1558,
                 reg1557,
                 reg1556,
                 wire1555,
                 wire1554,
                 wire1553,
                 wire1552,
                 wire1551,
                 (1'h0)};
  assign wire1551 = (wire1549[(4'hd):(1'h1)] ?
                        (8'ha7) : (&wire1548[(3'h4):(2'h2)]));
  assign wire1552 = wire1546;
  assign wire1553 = wire1550[(4'hc):(4'ha)];
  assign wire1554 = wire1547[(1'h0):(1'h0)];
  assign wire1555 = wire1548;
  always
    @(posedge clk) begin
      reg1556 <= ({(|$unsigned(((8'hb6) ? wire1554 : wire1549))),
          wire1546[(2'h2):(1'h1)]} || wire1553);
      if (((~&(|wire1548)) != (!(~($unsigned((8'hbe)) ?
          $unsigned(wire1550) : (wire1547 ~^ (8'ha1)))))))
        begin
          reg1557 <= {($unsigned({(~&wire1551)}) ?
                  {(~^reg1556), (~^(wire1546 <= wire1551))} : wire1550)};
        end
      else
        begin
          reg1557 <= (8'hb0);
          reg1558 <= {$unsigned($unsigned($unsigned(reg1557[(3'h7):(1'h0)]))),
              (wire1552[(2'h2):(1'h1)] ?
                  $unsigned(wire1548) : ((8'hb0) ?
                      (8'haa) : $unsigned(wire1554[(4'hc):(1'h0)])))};
        end
      if (((+$unsigned($unsigned({reg1557,
          (7'h40)}))) ^ $signed($unsigned((&(wire1550 >>> reg1557))))))
        begin
          if ({wire1549, $unsigned(wire1554[(3'h7):(3'h6)])})
            begin
              reg1559 <= (($unsigned({$signed((8'ha1))}) ?
                      wire1547[(2'h2):(1'h0)] : $unsigned(($signed(reg1558) ?
                          $signed(wire1554) : $unsigned(wire1555)))) ?
                  reg1556 : (($signed({wire1546,
                          (8'hbd)}) | (-$unsigned(wire1555))) ?
                      (-($signed(reg1556) ?
                          (^wire1548) : (^wire1548))) : wire1546[(1'h0):(1'h0)]));
              reg1560 <= ((wire1546 ?
                  reg1556 : {wire1548}) | $unsigned(($signed({wire1551}) <= ({(7'h40)} ^~ (~|reg1558)))));
              reg1561 <= wire1551[(1'h1):(1'h1)];
              reg1562 <= (($unsigned((reg1559 > $signed(reg1557))) ?
                      reg1561[(1'h1):(1'h1)] : $signed($unsigned((reg1557 ~^ wire1553)))) ?
                  $signed({$unsigned((wire1555 ? reg1557 : wire1548)),
                      reg1561}) : reg1556[(2'h3):(1'h0)]);
              reg1563 <= (($signed(($unsigned((7'h44)) ?
                      (&wire1552) : ((8'h9f) ? wire1549 : reg1557))) ?
                  $signed($signed((|reg1561))) : $unsigned(reg1561)) > $unsigned(reg1562[(1'h1):(1'h1)]));
            end
          else
            begin
              reg1559 <= wire1555;
              reg1560 <= $signed(wire1549[(2'h3):(1'h1)]);
              reg1561 <= ($signed((((reg1558 == reg1563) ^ (~^reg1557)) >>> $unsigned({wire1552}))) ?
                  (+wire1546[(2'h3):(2'h3)]) : (8'hb9));
              reg1562 <= {(^(!(reg1560 || (~reg1559))))};
              reg1563 <= ((($signed((~|wire1547)) <<< ((wire1551 > reg1558) ?
                      {reg1559, (7'h43)} : wire1550)) ?
                  (+$unsigned($unsigned(wire1554))) : $signed(wire1546[(1'h1):(1'h1)])) ^~ wire1552);
            end
          reg1564 <= reg1559[(3'h4):(1'h1)];
          reg1565 <= ((|reg1561[(2'h2):(1'h1)]) ? reg1556 : reg1561);
        end
      else
        begin
          if ($signed({($signed($signed(reg1563)) ?
                  ((8'hbf) != (reg1559 ?
                      wire1549 : (8'h9e))) : $unsigned(reg1560)),
              reg1563[(2'h3):(1'h0)]}))
            begin
              reg1559 <= wire1554[(4'hc):(3'h5)];
              reg1560 <= ($unsigned($unsigned({wire1555[(4'ha):(3'h6)],
                  ((8'h9f) & wire1549)})) >>> ($signed((^~wire1549)) == (^$signed(reg1558[(2'h2):(2'h2)]))));
              reg1561 <= reg1563[(4'hb):(4'ha)];
              reg1562 <= $signed((($signed((8'ha8)) ?
                      (-$signed(wire1549)) : wire1550[(1'h0):(1'h0)]) ?
                  ($unsigned(wire1552[(1'h0):(1'h0)]) ?
                      $signed((wire1550 ?
                          (8'hbf) : reg1565)) : wire1551[(1'h1):(1'h1)]) : (-((wire1552 ?
                          wire1551 : reg1565) ?
                      {reg1562, wire1552} : $unsigned(reg1558)))));
              reg1563 <= $signed(reg1563);
            end
          else
            begin
              reg1559 <= ((|wire1555) ?
                  ($unsigned(reg1564[(4'hb):(2'h2)]) ?
                      wire1546[(3'h4):(2'h3)] : $unsigned($unsigned($unsigned(wire1548)))) : $unsigned($unsigned($signed(reg1556))));
            end
          if (($signed(($unsigned(wire1547[(2'h2):(1'h1)]) < reg1565[(3'h6):(2'h2)])) ?
              $signed((reg1561[(2'h2):(1'h1)] >>> ($unsigned(wire1549) << ((8'hb4) <= reg1565)))) : wire1550))
            begin
              reg1564 <= wire1547[(2'h2):(1'h1)];
              reg1565 <= (-$unsigned($unsigned(wire1546)));
              reg1566 <= $unsigned(({($signed(reg1565) ?
                          (~^reg1561) : wire1552)} ?
                  ($unsigned(reg1562) ?
                      ($unsigned(wire1555) > wire1553[(3'h4):(1'h0)]) : (((8'hba) >> wire1555) ?
                          ((8'hb2) ?
                              (8'hbe) : reg1561) : $unsigned(reg1564))) : $unsigned($signed(wire1553))));
            end
          else
            begin
              reg1564 <= (wire1547 <<< $unsigned($signed($unsigned((|reg1566)))));
              reg1565 <= (^(~&$signed(((reg1563 ? reg1561 : reg1560) ?
                  $unsigned(reg1559) : $signed(wire1551)))));
              reg1566 <= reg1560;
              reg1567 <= ((~&((wire1546[(1'h0):(1'h0)] <<< (|wire1552)) * wire1547[(2'h2):(1'h1)])) ^~ ((wire1550[(5'h13):(1'h0)] ?
                  (~(wire1555 ^~ reg1557)) : (+reg1563[(3'h6):(3'h6)])) >> $unsigned((reg1557 ?
                  (reg1558 <= (8'h9d)) : (~&wire1552)))));
            end
        end
    end
  assign wire1568 = (wire1546 ?
                        reg1561 : $unsigned($signed((&(reg1567 ?
                            reg1562 : wire1549)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1508  (y, clk, wire1513, wire1512, wire1511, wire1510, wire1509);
  output wire [(32'h13b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire1513;
  input wire [(3'h6):(1'h0)] wire1512;
  input wire signed [(4'hf):(1'h0)] wire1511;
  input wire [(5'h15):(1'h0)] wire1510;
  input wire [(3'h5):(1'h0)] wire1509;
  wire signed [(2'h3):(1'h0)] wire1542;
  reg [(5'h13):(1'h0)] reg1541 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1540 = (1'h0);
  reg [(3'h4):(1'h0)] reg1539 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1538 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1537 = (1'h0);
  reg [(4'h8):(1'h0)] reg1536 = (1'h0);
  reg [(4'ha):(1'h0)] reg1535 = (1'h0);
  reg [(4'hc):(1'h0)] reg1534 = (1'h0);
  reg [(3'h6):(1'h0)] reg1533 = (1'h0);
  wire [(4'ha):(1'h0)] wire1532;
  wire [(4'hc):(1'h0)] wire1531;
  reg [(3'h5):(1'h0)] reg1530 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1529 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1528 = (1'h0);
  reg [(4'h8):(1'h0)] reg1527 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1526 = (1'h0);
  reg [(4'hc):(1'h0)] reg1525 = (1'h0);
  reg [(3'h6):(1'h0)] reg1524 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1523 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1522 = (1'h0);
  reg [(4'h9):(1'h0)] reg1521 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1520 = (1'h0);
  reg [(4'hc):(1'h0)] reg1519 = (1'h0);
  reg [(3'h4):(1'h0)] reg1518 = (1'h0);
  reg [(5'h11):(1'h0)] reg1517 = (1'h0);
  reg [(5'h15):(1'h0)] reg1516 = (1'h0);
  reg [(4'hb):(1'h0)] reg1515 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire1514;
  assign y = {wire1542,
                 reg1541,
                 reg1540,
                 reg1539,
                 reg1538,
                 reg1537,
                 reg1536,
                 reg1535,
                 reg1534,
                 reg1533,
                 wire1532,
                 wire1531,
                 reg1530,
                 reg1529,
                 reg1528,
                 reg1527,
                 reg1526,
                 reg1525,
                 reg1524,
                 reg1523,
                 reg1522,
                 reg1521,
                 reg1520,
                 reg1519,
                 reg1518,
                 reg1517,
                 reg1516,
                 reg1515,
                 wire1514,
                 (1'h0)};
  assign wire1514 = wire1510[(2'h3):(1'h1)];
  always
    @(posedge clk) begin
      if ((|wire1511))
        begin
          if ($unsigned(wire1513))
            begin
              reg1515 <= ({wire1509[(3'h5):(3'h4)]} ^~ ($signed($unsigned(wire1513)) + $signed($signed(((8'hb1) ?
                  wire1513 : wire1511)))));
            end
          else
            begin
              reg1515 <= ({(($unsigned(reg1515) ^~ $signed(wire1514)) ?
                      (reg1515[(3'h4):(2'h2)] ^~ (reg1515 ?
                          wire1511 : (8'ha9))) : $signed((wire1513 ?
                          wire1511 : (8'hbb))))} ^ $unsigned(wire1513));
              reg1516 <= ((((wire1512 + (reg1515 <= wire1512)) ?
                  (~|(wire1511 ~^ (8'ha7))) : (wire1513 ?
                      wire1512[(2'h2):(1'h0)] : $unsigned(wire1511))) <= ($signed(wire1514) <= (7'h44))) & (-({$signed((8'hb4)),
                  (wire1513 ? wire1511 : (7'h42))} <<< (^~{(7'h44),
                  (8'had)}))));
              reg1517 <= wire1512;
              reg1518 <= ($signed(wire1514) * {$signed((wire1510[(3'h6):(1'h0)] >> (-reg1517)))});
              reg1519 <= wire1509;
            end
          reg1520 <= {wire1514};
          reg1521 <= ({(($signed(reg1519) ?
                      $unsigned((8'ha5)) : ((8'ha6) ?
                          wire1514 : reg1517)) >>> (^(wire1513 << (8'hbd))))} ?
              wire1511 : $unsigned($unsigned(((+reg1520) ^ reg1515[(2'h2):(1'h1)]))));
        end
      else
        begin
          if ($signed($signed(((~&(reg1520 + reg1519)) ?
              reg1520[(4'h9):(3'h5)] : $unsigned((!reg1521))))))
            begin
              reg1515 <= ((wire1513 || (~&wire1510[(4'he):(4'hb)])) ?
                  reg1521[(1'h0):(1'h0)] : (8'ha7));
              reg1516 <= (reg1519 && (~&{(((8'h9d) >= reg1515) ?
                      (reg1519 <= wire1512) : $signed((8'ha1))),
                  (wire1509[(1'h0):(1'h0)] == {wire1512})}));
            end
          else
            begin
              reg1515 <= $unsigned(($signed({(~|wire1511)}) ?
                  reg1517[(4'h8):(3'h7)] : wire1513));
              reg1516 <= reg1519[(1'h1):(1'h0)];
              reg1517 <= wire1510[(4'hf):(4'h9)];
              reg1518 <= (reg1518[(2'h3):(1'h1)] >> reg1520[(1'h1):(1'h1)]);
            end
          reg1519 <= {(~^$unsigned((~^$unsigned(wire1513)))),
              $unsigned($signed(({wire1514, reg1520} ?
                  reg1516 : $signed(wire1509))))};
          reg1520 <= reg1521[(4'h9):(1'h1)];
          reg1521 <= {$signed(reg1516)};
          reg1522 <= $signed($unsigned(reg1521));
        end
      if ((^~$signed(reg1520[(1'h0):(1'h0)])))
        begin
          reg1523 <= ($unsigned(reg1521) ^ reg1516);
          reg1524 <= $signed($unsigned($signed($signed({reg1515, reg1520}))));
          reg1525 <= $unsigned(reg1524[(2'h3):(2'h3)]);
          reg1526 <= wire1513[(4'h8):(1'h1)];
          reg1527 <= ($unsigned((($unsigned(wire1514) >= wire1513[(1'h0):(1'h0)]) ?
                  $unsigned($signed(wire1512)) : {$unsigned(reg1524),
                      (reg1519 <<< (8'ha5))})) ?
              (~^($unsigned($unsigned(wire1510)) ?
                  reg1519 : $unsigned($signed((8'ha8))))) : {(8'ha6), (8'ha9)});
        end
      else
        begin
          if ((~|{({wire1509[(1'h1):(1'h1)], $signed(reg1527)} ?
                  $unsigned(reg1519) : {(+reg1519), (reg1523 | reg1523)}),
              reg1521}))
            begin
              reg1523 <= {wire1509[(3'h4):(1'h1)],
                  $unsigned((reg1524 ?
                      $unsigned(reg1525[(4'hb):(3'h5)]) : (~^(8'hb7))))};
              reg1524 <= (~|(|$signed($signed($unsigned(reg1517)))));
              reg1525 <= $signed($unsigned((~&$unsigned($unsigned(reg1523)))));
              reg1526 <= wire1509;
            end
          else
            begin
              reg1523 <= $unsigned((~$unsigned((^~$unsigned((8'hb7))))));
            end
          if ({(^~wire1509[(3'h5):(2'h3)]),
              ($unsigned((!$signed(reg1522))) ?
                  (8'hb6) : $unsigned($unsigned((reg1525 ?
                      wire1513 : reg1520))))})
            begin
              reg1527 <= {($signed({reg1521}) <<< wire1513[(1'h1):(1'h1)])};
              reg1528 <= ((+$unsigned(((+wire1510) ?
                      ((8'h9d) ? reg1518 : reg1516) : $signed(wire1511)))) ?
                  (^$signed((8'hbf))) : $signed({$signed({reg1521}),
                      wire1512[(1'h0):(1'h0)]}));
            end
          else
            begin
              reg1527 <= wire1511;
              reg1528 <= ((!(reg1522[(4'hc):(1'h0)] ?
                  ($signed(reg1520) >> wire1510[(4'ha):(3'h7)]) : ($unsigned(reg1528) ?
                      (wire1513 ?
                          reg1525 : reg1523) : (reg1519 <= reg1519)))) <= reg1526);
            end
          reg1529 <= $signed($unsigned($unsigned(((reg1518 && reg1516) >> reg1528[(2'h3):(1'h0)]))));
          reg1530 <= {$signed(reg1528),
              {(~&reg1520), (reg1529 <<< {$unsigned(reg1526)})}};
        end
    end
  assign wire1531 = wire1509;
  assign wire1532 = reg1527;
  always
    @(posedge clk) begin
      reg1533 <= $unsigned({(8'hbb)});
      reg1534 <= (~^$signed($unsigned(({wire1511} ?
          (wire1511 & wire1511) : reg1530[(3'h5):(2'h2)]))));
      reg1535 <= (wire1510[(3'h7):(3'h4)] ?
          reg1519[(4'h9):(3'h7)] : $signed((~&((reg1530 - (8'hbc)) & $signed(reg1517)))));
      if (($unsigned(reg1515[(2'h2):(1'h1)]) ?
          (reg1516[(5'h12):(4'he)] ?
              $signed($signed(((7'h43) ?
                  reg1524 : wire1510))) : reg1521) : (reg1516[(5'h13):(4'he)] ?
              ((reg1522[(4'h8):(1'h0)] ? (~|wire1513) : (^reg1529)) ?
                  {(reg1535 <<< reg1522)} : $signed($signed((8'hbd)))) : (wire1509[(3'h5):(2'h3)] == reg1517[(1'h1):(1'h0)]))))
        begin
          reg1536 <= reg1523[(3'h4):(2'h3)];
        end
      else
        begin
          if ({wire1532, $signed((wire1532[(1'h1):(1'h0)] > (8'h9d)))})
            begin
              reg1536 <= {(~^reg1530)};
            end
          else
            begin
              reg1536 <= reg1515;
              reg1537 <= {$unsigned((~(^~(reg1527 ? wire1514 : reg1519)))),
                  {$signed(((-reg1520) << $signed(reg1524))),
                      (!$signed((reg1526 <= (8'hb6))))}};
              reg1538 <= (^~(wire1509 ?
                  {(~^(^~reg1536)),
                      (reg1530 ?
                          {wire1531} : (reg1529 & reg1530))} : $unsigned($signed($unsigned(reg1536)))));
              reg1539 <= reg1530[(3'h5):(1'h1)];
            end
          reg1540 <= reg1519[(1'h1):(1'h1)];
          reg1541 <= {reg1521[(2'h3):(2'h2)]};
        end
    end
  assign wire1542 = ($signed($unsigned((~(~|wire1532)))) ?
                        wire1509[(3'h5):(1'h1)] : $unsigned($unsigned(wire1509)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1374
#( parameter param1504 = (!(^((~((8'hb3) ? (8'hbb) : (8'hb9))) | (|(~^(8'ha0))))))
, parameter param1505 = (({(~^(param1504 >>> param1504))} ^ (&{(param1504 > (8'ha6)), ((7'h40) ? param1504 : param1504)})) > param1504) )
(y, clk, wire1379, wire1378, wire1377, wire1376, wire1375);
  output wire [(32'h541):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire1379;
  input wire [(4'hc):(1'h0)] wire1378;
  input wire signed [(5'h11):(1'h0)] wire1377;
  input wire signed [(4'hf):(1'h0)] wire1376;
  input wire signed [(3'h4):(1'h0)] wire1375;
  wire signed [(3'h6):(1'h0)] wire1503;
  wire signed [(5'h12):(1'h0)] wire1502;
  wire signed [(5'h11):(1'h0)] wire1501;
  wire [(4'hf):(1'h0)] wire1500;
  wire [(3'h5):(1'h0)] wire1499;
  wire [(4'hf):(1'h0)] wire1498;
  reg signed [(4'ha):(1'h0)] reg1497 = (1'h0);
  reg [(4'he):(1'h0)] reg1496 = (1'h0);
  reg [(4'he):(1'h0)] reg1495 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire1494;
  wire [(5'h12):(1'h0)] wire1493;
  wire [(5'h13):(1'h0)] wire1492;
  reg signed [(2'h3):(1'h0)] reg1491 = (1'h0);
  reg [(2'h3):(1'h0)] reg1490 = (1'h0);
  reg [(2'h3):(1'h0)] reg1489 = (1'h0);
  reg [(5'h13):(1'h0)] reg1488 = (1'h0);
  reg [(3'h7):(1'h0)] reg1487 = (1'h0);
  reg [(2'h2):(1'h0)] reg1486 = (1'h0);
  reg [(5'h15):(1'h0)] reg1485 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1484 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1483 = (1'h0);
  reg [(3'h6):(1'h0)] reg1482 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1481 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire1480;
  wire signed [(4'hd):(1'h0)] wire1479;
  reg signed [(3'h6):(1'h0)] reg1478 = (1'h0);
  reg [(4'hc):(1'h0)] reg1477 = (1'h0);
  reg [(4'ha):(1'h0)] reg1476 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1475 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1474 = (1'h0);
  reg [(4'hc):(1'h0)] reg1473 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1472 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1471 = (1'h0);
  reg [(4'hb):(1'h0)] reg1470 = (1'h0);
  reg [(4'hc):(1'h0)] reg1469 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1468 = (1'h0);
  reg [(5'h12):(1'h0)] reg1467 = (1'h0);
  reg [(3'h5):(1'h0)] reg1466 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1465 = (1'h0);
  reg [(4'h8):(1'h0)] reg1464 = (1'h0);
  reg [(3'h6):(1'h0)] reg1463 = (1'h0);
  reg [(4'hc):(1'h0)] reg1462 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1461 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1460 = (1'h0);
  reg [(5'h11):(1'h0)] reg1459 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire1458;
  reg [(2'h2):(1'h0)] reg1457 = (1'h0);
  reg [(2'h3):(1'h0)] reg1456 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1455 = (1'h0);
  reg [(4'h8):(1'h0)] reg1454 = (1'h0);
  reg [(5'h15):(1'h0)] reg1453 = (1'h0);
  reg [(5'h14):(1'h0)] reg1452 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1451 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1450 = (1'h0);
  reg [(4'h9):(1'h0)] reg1449 = (1'h0);
  reg [(3'h4):(1'h0)] reg1448 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1447 = (1'h0);
  reg [(4'ha):(1'h0)] reg1446 = (1'h0);
  reg [(4'ha):(1'h0)] reg1445 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1444 = (1'h0);
  reg [(2'h2):(1'h0)] reg1443 = (1'h0);
  reg [(3'h5):(1'h0)] reg1442 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1441 = (1'h0);
  reg [(4'h8):(1'h0)] reg1440 = (1'h0);
  reg [(5'h15):(1'h0)] reg1439 = (1'h0);
  reg [(2'h2):(1'h0)] reg1438 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1437 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1436 = (1'h0);
  reg [(4'hc):(1'h0)] reg1435 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1434 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1433 = (1'h0);
  reg [(4'he):(1'h0)] reg1432 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1431 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1430 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1429 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1428 = (1'h0);
  reg [(5'h11):(1'h0)] reg1427 = (1'h0);
  reg [(4'hc):(1'h0)] reg1426 = (1'h0);
  reg [(3'h6):(1'h0)] reg1425 = (1'h0);
  reg [(5'h10):(1'h0)] reg1424 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1423 = (1'h0);
  reg [(3'h4):(1'h0)] reg1422 = (1'h0);
  reg [(5'h12):(1'h0)] reg1421 = (1'h0);
  reg [(4'he):(1'h0)] reg1420 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1419 = (1'h0);
  reg [(4'ha):(1'h0)] reg1418 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1417 = (1'h0);
  wire [(5'h14):(1'h0)] wire1416;
  wire signed [(5'h13):(1'h0)] wire1415;
  reg signed [(3'h4):(1'h0)] reg1414 = (1'h0);
  reg [(4'hc):(1'h0)] reg1413 = (1'h0);
  reg [(4'hf):(1'h0)] reg1412 = (1'h0);
  reg [(3'h4):(1'h0)] reg1411 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1410 = (1'h0);
  reg [(5'h10):(1'h0)] reg1409 = (1'h0);
  reg [(4'hd):(1'h0)] reg1408 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1407 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1406 = (1'h0);
  reg [(3'h5):(1'h0)] reg1405 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1404 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1403 = (1'h0);
  reg [(5'h11):(1'h0)] reg1402 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1401 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1400 = (1'h0);
  reg [(3'h6):(1'h0)] reg1399 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1398 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1397 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1396 = (1'h0);
  reg [(5'h11):(1'h0)] reg1395 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1394 = (1'h0);
  reg [(3'h7):(1'h0)] reg1393 = (1'h0);
  reg [(3'h4):(1'h0)] reg1392 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1391 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1390 = (1'h0);
  reg [(4'h9):(1'h0)] reg1389 = (1'h0);
  reg [(5'h14):(1'h0)] reg1388 = (1'h0);
  reg [(3'h6):(1'h0)] reg1387 = (1'h0);
  reg [(5'h10):(1'h0)] reg1386 = (1'h0);
  reg [(4'ha):(1'h0)] reg1385 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1384 = (1'h0);
  reg [(4'h8):(1'h0)] reg1383 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1382 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire1381;
  wire [(3'h4):(1'h0)] wire1380;
  assign y = {wire1503,
                 wire1502,
                 wire1501,
                 wire1500,
                 wire1499,
                 wire1498,
                 reg1497,
                 reg1496,
                 reg1495,
                 wire1494,
                 wire1493,
                 wire1492,
                 reg1491,
                 reg1490,
                 reg1489,
                 reg1488,
                 reg1487,
                 reg1486,
                 reg1485,
                 reg1484,
                 reg1483,
                 reg1482,
                 reg1481,
                 wire1480,
                 wire1479,
                 reg1478,
                 reg1477,
                 reg1476,
                 reg1475,
                 reg1474,
                 reg1473,
                 reg1472,
                 reg1471,
                 reg1470,
                 reg1469,
                 reg1468,
                 reg1467,
                 reg1466,
                 reg1465,
                 reg1464,
                 reg1463,
                 reg1462,
                 reg1461,
                 reg1460,
                 reg1459,
                 wire1458,
                 reg1457,
                 reg1456,
                 reg1455,
                 reg1454,
                 reg1453,
                 reg1452,
                 reg1451,
                 reg1450,
                 reg1449,
                 reg1448,
                 reg1447,
                 reg1446,
                 reg1445,
                 reg1444,
                 reg1443,
                 reg1442,
                 reg1441,
                 reg1440,
                 reg1439,
                 reg1438,
                 reg1437,
                 reg1436,
                 reg1435,
                 reg1434,
                 reg1433,
                 reg1432,
                 reg1431,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1427,
                 reg1426,
                 reg1425,
                 reg1424,
                 reg1423,
                 reg1422,
                 reg1421,
                 reg1420,
                 reg1419,
                 reg1418,
                 reg1417,
                 wire1416,
                 wire1415,
                 reg1414,
                 reg1413,
                 reg1412,
                 reg1411,
                 reg1410,
                 reg1409,
                 reg1408,
                 reg1407,
                 reg1406,
                 reg1405,
                 reg1404,
                 reg1403,
                 reg1402,
                 reg1401,
                 reg1400,
                 reg1399,
                 reg1398,
                 reg1397,
                 reg1396,
                 reg1395,
                 reg1394,
                 reg1393,
                 reg1392,
                 reg1391,
                 reg1390,
                 reg1389,
                 reg1388,
                 reg1387,
                 reg1386,
                 reg1385,
                 reg1384,
                 reg1383,
                 reg1382,
                 wire1381,
                 wire1380,
                 (1'h0)};
  assign wire1380 = ($unsigned((wire1379[(4'h8):(2'h3)] < wire1378[(2'h2):(2'h2)])) ~^ wire1377);
  assign wire1381 = $unsigned($signed(($unsigned((wire1377 << wire1376)) - $unsigned(((8'ha3) & wire1379)))));
  always
    @(posedge clk) begin
      if ($signed(((($signed(wire1378) ?
          wire1379 : $signed((8'hbf))) << (~^$unsigned(wire1381))) != $unsigned(wire1376))))
        begin
          reg1382 <= wire1375;
          if ($unsigned(reg1382))
            begin
              reg1383 <= (wire1378[(4'h9):(3'h5)] ?
                  (^(&(wire1380 & wire1378[(4'h8):(3'h7)]))) : $unsigned((($signed(wire1379) ?
                      reg1382[(1'h1):(1'h1)] : $signed(wire1381)) <= (|(|wire1380)))));
              reg1384 <= wire1378[(1'h1):(1'h0)];
              reg1385 <= wire1378;
            end
          else
            begin
              reg1383 <= {$signed(wire1381[(2'h2):(1'h0)]),
                  (reg1384 ?
                      wire1378[(4'h9):(1'h1)] : (wire1375 - (+wire1376)))};
              reg1384 <= ((wire1379[(1'h1):(1'h1)] != $signed((8'hb8))) >= wire1380[(1'h1):(1'h0)]);
            end
          if (($unsigned({(reg1384[(2'h2):(1'h1)] ^ (+wire1380))}) ?
              wire1380 : ({{$signed(wire1378)}} <<< (reg1384 <<< {(reg1384 ?
                      reg1385 : wire1381)}))))
            begin
              reg1386 <= wire1377;
              reg1387 <= reg1384;
              reg1388 <= ((({$unsigned(wire1378)} ?
                          $signed($unsigned((8'ha8))) : $signed($unsigned(reg1384))) ?
                      ($signed($signed(wire1377)) ^ ($unsigned(wire1379) && (wire1381 && wire1378))) : (wire1375[(1'h0):(1'h0)] != {(!reg1383)})) ?
                  ((~^{((8'hab) - wire1377)}) <= $signed(reg1385)) : (~(reg1383 ?
                      wire1378[(4'hc):(3'h4)] : {wire1377[(4'he):(3'h4)],
                          $signed(wire1381)})));
              reg1389 <= ({$signed(((wire1376 ?
                      reg1384 : reg1388) << wire1375))} ~^ (wire1379[(1'h0):(1'h0)] ?
                  ((reg1383 ?
                      (reg1388 ? (8'ha8) : reg1383) : ((8'hbf) ?
                          wire1375 : reg1382)) & reg1386) : (reg1388[(3'h6):(3'h5)] + (^$unsigned(reg1382)))));
            end
          else
            begin
              reg1386 <= ((+((^~$unsigned(wire1381)) >>> $unsigned($signed(wire1376)))) & ({(^~reg1389[(1'h1):(1'h1)])} & $unsigned($signed(reg1383))));
            end
          if ((8'hb4))
            begin
              reg1390 <= reg1388[(4'h9):(2'h2)];
              reg1391 <= ((-(~|wire1379[(3'h5):(3'h4)])) ?
                  wire1377[(2'h3):(2'h3)] : (!$unsigned(((&wire1376) + $unsigned(reg1386)))));
              reg1392 <= {(wire1375 == {((wire1381 ? wire1375 : reg1383) ?
                          {reg1391, reg1384} : (wire1376 == reg1383)),
                      reg1386[(2'h3):(2'h2)]}),
                  reg1384[(2'h2):(1'h1)]};
              reg1393 <= ($signed(wire1377) ?
                  wire1376[(4'hd):(3'h6)] : reg1384);
              reg1394 <= ((&($signed(reg1383) ?
                      ($unsigned((7'h44)) ~^ $unsigned(reg1383)) : (8'hba))) ?
                  {(wire1381 ?
                          wire1376 : $signed(wire1377))} : (|$signed(wire1379)));
            end
          else
            begin
              reg1390 <= $signed((!(^((reg1389 < reg1390) ?
                  (&reg1392) : (8'ha2)))));
              reg1391 <= (|reg1394[(3'h4):(2'h3)]);
              reg1392 <= reg1384[(1'h1):(1'h0)];
            end
          reg1395 <= reg1388[(5'h11):(4'h9)];
        end
      else
        begin
          reg1382 <= (^~$signed((!(reg1387 ?
              $unsigned((7'h40)) : reg1391[(2'h2):(1'h1)]))));
          if ((wire1381[(1'h0):(1'h0)] ?
              reg1393[(1'h1):(1'h0)] : $unsigned($signed($signed($unsigned(reg1388))))))
            begin
              reg1383 <= (~^reg1390);
              reg1384 <= (reg1382 ?
                  (-$signed((((8'hb5) ? reg1385 : wire1379) ?
                      reg1395 : $unsigned(reg1383)))) : (8'ha6));
              reg1385 <= reg1386;
            end
          else
            begin
              reg1383 <= (wire1376[(3'h6):(2'h3)] ^~ ({reg1391[(2'h3):(1'h1)],
                      {reg1389, $signed(reg1390)}} ?
                  $signed($unsigned($unsigned(reg1392))) : (|(|(reg1392 ?
                      reg1390 : wire1380)))));
              reg1384 <= wire1377;
              reg1385 <= $signed(wire1377);
              reg1386 <= (+({reg1391[(1'h0):(1'h0)]} & {(~reg1392[(3'h4):(3'h4)])}));
              reg1387 <= ((~|wire1380) ?
                  reg1389[(3'h7):(2'h2)] : $unsigned((^(reg1394[(1'h1):(1'h1)] ?
                      (reg1392 ? reg1385 : wire1378) : (^(8'hba))))));
            end
          if (reg1395)
            begin
              reg1388 <= $signed({$signed(((reg1384 ? reg1389 : wire1378) ?
                      ((8'ha2) ~^ reg1393) : ((8'hac) ? reg1388 : reg1395)))});
              reg1389 <= {reg1395[(3'h5):(1'h0)]};
            end
          else
            begin
              reg1388 <= wire1380[(3'h4):(2'h3)];
              reg1389 <= {(reg1384 ?
                      $signed(wire1379) : $signed((reg1393 > (reg1384 ?
                          reg1387 : (7'h42)))))};
              reg1390 <= ($unsigned((+reg1388[(4'hd):(3'h4)])) ?
                  reg1393[(1'h1):(1'h0)] : (~|$signed(({wire1380,
                      wire1376} == (+reg1384)))));
            end
          reg1391 <= $unsigned($unsigned((reg1382[(2'h2):(1'h1)] ?
              $signed(reg1383) : ($signed(reg1385) >> (reg1395 ~^ reg1387)))));
          reg1392 <= (($signed(($unsigned(reg1391) ?
                  $unsigned(reg1384) : {reg1388})) > (~^(reg1383[(4'h8):(2'h3)] ?
                  ((8'haa) ? wire1378 : reg1388) : $signed((8'haf))))) ?
              reg1384[(1'h1):(1'h0)] : ($signed(((&wire1379) << wire1378)) ?
                  $signed(wire1377[(3'h4):(1'h0)]) : reg1386[(1'h0):(1'h0)]));
        end
      reg1396 <= (~|(~&((((8'hb6) ^ (8'ha4)) ^~ wire1377[(4'ha):(2'h3)]) ?
          (8'ha3) : reg1388)));
      reg1397 <= {$unsigned(($signed((+reg1396)) == $signed((~reg1390))))};
      if ({(+{(reg1384[(2'h2):(1'h1)] | (wire1375 != wire1376)),
              (reg1395 ^~ reg1396)}),
          reg1382[(1'h0):(1'h0)]})
        begin
          reg1398 <= reg1391;
          reg1399 <= reg1384;
          reg1400 <= (~&(reg1395[(2'h2):(1'h1)] ?
              {$signed(reg1397), (8'ha3)} : $signed(reg1392[(1'h0):(1'h0)])));
          if ((^(~|$unsigned(wire1376[(4'ha):(3'h6)]))))
            begin
              reg1401 <= ({($unsigned((wire1379 ?
                      wire1377 : reg1384)) ^~ ($unsigned((8'had)) ~^ (8'hbf))),
                  (~|reg1386)} - $unsigned($unsigned(reg1390)));
              reg1402 <= (8'ha8);
              reg1403 <= reg1401[(4'hf):(3'h6)];
            end
          else
            begin
              reg1401 <= $signed((reg1397 ?
                  reg1390[(4'h8):(3'h4)] : (((^~wire1381) - (wire1378 ?
                          reg1396 : reg1397)) ?
                      reg1398 : ($signed(reg1389) ?
                          $unsigned(reg1392) : (reg1395 ?
                              wire1375 : wire1380)))));
              reg1402 <= $unsigned(((($unsigned((7'h43)) | (+wire1378)) ?
                  (wire1378[(2'h3):(2'h2)] & {wire1381}) : $signed((reg1386 >>> reg1392))) << reg1402[(4'hc):(3'h7)]));
            end
        end
      else
        begin
          reg1398 <= wire1376[(2'h2):(1'h0)];
          reg1399 <= (8'hac);
          reg1400 <= $unsigned((($unsigned((~^wire1376)) ?
                  (reg1391[(1'h1):(1'h1)] * {(8'h9e)}) : {reg1388[(4'h9):(1'h0)],
                      reg1400}) ?
              $signed(reg1386) : wire1378[(3'h5):(3'h5)]));
          reg1401 <= {(wire1378 ?
                  $unsigned((^~(~^wire1380))) : $signed((+$signed((8'hb0))))),
              (($unsigned(reg1384[(2'h2):(2'h2)]) ?
                      ((wire1379 <= wire1378) ?
                          reg1396[(3'h4):(1'h1)] : (reg1384 >>> (8'hb3))) : ($unsigned(reg1388) ?
                          (wire1379 >= reg1389) : (8'ha0))) ?
                  reg1383[(2'h2):(1'h0)] : $signed(((&(8'hb6)) ?
                      $unsigned((7'h42)) : (reg1394 + reg1402))))};
          reg1402 <= (~^$signed({(~^$signed(reg1390))}));
        end
      if ($signed(reg1399[(3'h5):(2'h3)]))
        begin
          reg1404 <= ($unsigned($unsigned(((wire1376 ?
                  reg1399 : (8'hba)) * (reg1393 && reg1390)))) ?
              wire1375 : (&{($signed(wire1379) ?
                      $unsigned(reg1392) : $unsigned(reg1383))}));
          if ((|(8'hbe)))
            begin
              reg1405 <= (~(reg1404[(1'h0):(1'h0)] ?
                  {((&wire1378) ? (~|reg1384) : wire1377[(5'h11):(3'h7)]),
                      $unsigned((~^reg1398))} : (|reg1383)));
              reg1406 <= reg1397[(2'h2):(1'h0)];
            end
          else
            begin
              reg1405 <= (wire1380 ?
                  {($unsigned((reg1394 ?
                          (8'hab) : wire1381)) >= $signed({(7'h43)}))} : (($signed(reg1404[(4'h8):(2'h2)]) ?
                          {(~^reg1386),
                              (reg1388 >= (8'ha3))} : wire1381[(1'h0):(1'h0)]) ?
                      {$signed(reg1406)} : (!(^~$signed(wire1375)))));
              reg1406 <= $unsigned((8'hb3));
              reg1407 <= $signed(($signed($unsigned((wire1381 & (7'h42)))) && reg1402[(4'hb):(2'h3)]));
              reg1408 <= reg1383[(3'h6):(2'h2)];
            end
          reg1409 <= reg1393;
          reg1410 <= $signed({reg1394,
              $unsigned($signed((reg1408 ? (8'ha1) : reg1404)))});
          if (((7'h42) ?
              $unsigned((reg1398 ?
                  (|$unsigned((8'ha6))) : $signed($unsigned(reg1403)))) : reg1401))
            begin
              reg1411 <= $signed($signed($signed(($signed((8'hac)) <= (8'hba)))));
              reg1412 <= ((+reg1385) ?
                  (^~$unsigned(((reg1403 ?
                      reg1396 : reg1410) >>> (^(7'h42))))) : $signed($signed($signed((reg1407 ?
                      (7'h40) : reg1391)))));
              reg1413 <= ((+$unsigned(reg1405)) == wire1377[(1'h1):(1'h1)]);
              reg1414 <= ($signed($signed(($unsigned(reg1395) ^ {reg1412,
                      reg1396}))) ?
                  wire1375[(1'h0):(1'h0)] : $signed((reg1389[(4'h8):(3'h7)] || $unsigned((!reg1386)))));
            end
          else
            begin
              reg1411 <= reg1406[(3'h5):(3'h5)];
              reg1412 <= $signed($signed($signed((~|wire1377))));
              reg1413 <= reg1393[(3'h7):(2'h2)];
              reg1414 <= wire1380;
            end
        end
      else
        begin
          reg1404 <= ($signed(reg1384) ^~ reg1406);
          if (reg1400)
            begin
              reg1405 <= $unsigned(({(&reg1409)} ?
                  (((&reg1413) ?
                      (8'hbb) : wire1381[(1'h1):(1'h1)]) >> ($unsigned(reg1392) ?
                      $unsigned(reg1412) : reg1390)) : wire1380[(2'h2):(2'h2)]));
              reg1406 <= reg1406[(1'h1):(1'h1)];
              reg1407 <= (+$unsigned($unsigned(reg1396)));
              reg1408 <= (((~|wire1380) ? reg1394 : wire1379[(4'hd):(4'hd)]) ?
                  ($unsigned((^(wire1378 ?
                      wire1379 : reg1410))) + reg1386) : (8'had));
            end
          else
            begin
              reg1405 <= reg1400[(1'h0):(1'h0)];
              reg1406 <= (8'hbf);
              reg1407 <= (reg1385[(3'h4):(1'h1)] - (~^(reg1407[(4'hd):(3'h7)] & (reg1413 ?
                  (reg1401 ? reg1388 : wire1379) : (reg1390 <= reg1394)))));
              reg1408 <= reg1413;
              reg1409 <= $unsigned((~$unsigned($signed($signed(reg1391)))));
            end
          reg1410 <= ((^~(~|((~wire1377) ?
                  wire1380 : reg1389[(3'h6):(3'h6)]))) ?
              ((($unsigned(reg1401) >> wire1376) ?
                  reg1402 : ($signed(reg1388) <= $unsigned(reg1386))) >= (|((reg1399 ?
                      (8'hb7) : reg1407) ?
                  {reg1394} : $signed(reg1400)))) : $signed($signed(($signed((8'ha8)) ?
                  reg1384[(1'h1):(1'h1)] : $signed(reg1388)))));
        end
    end
  assign wire1415 = (((reg1403[(2'h2):(1'h0)] <= ({(8'had)} ?
                                (~|reg1404) : $unsigned(reg1405))) ?
                            (reg1391[(1'h1):(1'h1)] - $signed((8'ha6))) : reg1383) ?
                        reg1405 : reg1404);
  assign wire1416 = reg1387;
  always
    @(posedge clk) begin
      if (($unsigned($unsigned($signed((|reg1396)))) > wire1416[(4'h8):(3'h5)]))
        begin
          reg1417 <= reg1398[(4'hb):(3'h5)];
        end
      else
        begin
          if ({$signed(reg1414[(1'h1):(1'h1)]),
              {$signed(reg1407[(1'h0):(1'h0)]),
                  (((reg1414 ? reg1392 : reg1401) ? reg1402 : (~^reg1403)) ?
                      $signed((reg1405 ?
                          reg1391 : reg1411)) : reg1405[(3'h5):(3'h4)])}})
            begin
              reg1417 <= (^~(^((!{reg1387, (8'ha5)}) ?
                  ($signed(reg1417) ?
                      (reg1385 ^ reg1389) : reg1395[(1'h1):(1'h0)]) : (^(reg1385 || reg1396)))));
              reg1418 <= ($signed(reg1402[(4'h9):(3'h5)]) ?
                  $unsigned(($signed(((8'hbe) ? reg1389 : reg1403)) ?
                      (^~(~|reg1404)) : ({reg1411,
                          reg1385} & $signed((8'hbf))))) : reg1384[(2'h2):(1'h1)]);
              reg1419 <= $signed({({{reg1395, wire1381}} ?
                      wire1415[(4'h8):(4'h8)] : wire1380[(2'h3):(2'h2)]),
                  (~$signed((reg1414 | (8'hbf))))});
              reg1420 <= wire1379;
            end
          else
            begin
              reg1417 <= $signed((7'h41));
              reg1418 <= $unsigned((~^(~reg1404)));
              reg1419 <= reg1408[(3'h4):(1'h0)];
              reg1420 <= reg1390;
            end
          reg1421 <= reg1403;
          if ({((~reg1384[(1'h1):(1'h1)]) > ((!(reg1402 ? reg1407 : reg1387)) ?
                  reg1418 : reg1414)),
              ((&(reg1391 >>> $signed(wire1379))) ?
                  reg1408[(4'h8):(3'h7)] : $signed($signed((wire1415 > reg1383))))})
            begin
              reg1422 <= {reg1390[(4'h8):(2'h2)], (^~{reg1418})};
              reg1423 <= {reg1397};
              reg1424 <= reg1387[(1'h0):(1'h0)];
              reg1425 <= $unsigned(((({reg1385, (8'hbb)} ?
                          {wire1416} : (wire1378 & reg1400)) ?
                      reg1405 : $unsigned((-reg1417))) ?
                  (reg1410[(3'h4):(1'h0)] ?
                      (reg1393 && reg1420[(4'ha):(4'h9)]) : $signed(((8'ha1) >>> reg1410))) : reg1385[(4'h8):(3'h7)]));
              reg1426 <= $unsigned(wire1375);
            end
          else
            begin
              reg1422 <= (|(|(+reg1409[(4'hd):(4'hc)])));
              reg1423 <= wire1380;
              reg1424 <= (!reg1387);
            end
          reg1427 <= reg1389[(4'h9):(3'h7)];
          if ($signed({(((wire1416 < reg1390) ?
                  $signed((8'hb8)) : {reg1418, (8'hae)}) ^~ (((8'hbb) ?
                  wire1380 : reg1427) ~^ (~reg1390))),
              (8'ha4)}))
            begin
              reg1428 <= $signed({$unsigned(({reg1419,
                      wire1380} & reg1427[(4'h8):(1'h0)]))});
            end
          else
            begin
              reg1428 <= ((^~$signed({{(8'hb0),
                      reg1390}})) ^~ ($unsigned(((reg1407 ? reg1409 : reg1412) ?
                      (reg1406 ? reg1407 : reg1388) : $signed((8'hb5)))) ?
                  (reg1385[(4'h9):(4'h9)] ^ (~&$unsigned(wire1416))) : reg1424[(1'h1):(1'h1)]));
              reg1429 <= (^((((&reg1395) ? reg1387 : reg1424[(3'h5):(3'h4)]) ?
                  $signed(reg1403) : reg1399[(1'h0):(1'h0)]) * reg1389));
              reg1430 <= wire1416[(2'h2):(2'h2)];
              reg1431 <= (~|reg1408[(4'h8):(3'h7)]);
              reg1432 <= reg1410;
            end
        end
      if (reg1409[(2'h2):(1'h0)])
        begin
          if ({((reg1405[(2'h2):(1'h0)] ?
                  $signed(reg1387[(3'h5):(2'h2)]) : $signed((reg1383 < reg1429))) & reg1419)})
            begin
              reg1433 <= (!((reg1414 << {reg1418[(3'h6):(3'h4)], reg1410}) ?
                  ($signed(reg1426[(4'h9):(4'h8)]) ?
                      ((reg1402 - reg1382) ?
                          (-reg1410) : reg1387[(2'h2):(1'h1)]) : (|{reg1390,
                          reg1418})) : (($unsigned(reg1386) >= (reg1430 ?
                          wire1379 : reg1391)) ?
                      ({reg1431} & (-reg1429)) : ((reg1404 ?
                          reg1385 : reg1404) < (~|wire1376)))));
              reg1434 <= (~|$signed(reg1405));
              reg1435 <= ((+$unsigned((~&$unsigned(reg1433)))) ?
                  $signed((((^~reg1390) ?
                          $unsigned((8'hb3)) : (reg1428 > reg1390)) ?
                      (!{reg1433,
                          reg1417}) : reg1420)) : (+(reg1424[(3'h4):(1'h0)] ?
                      reg1423 : ($signed(reg1413) >>> {(8'hb0), (8'hb4)}))));
              reg1436 <= ((~reg1435) ?
                  (~|reg1389[(3'h6):(2'h2)]) : (reg1408[(4'ha):(3'h5)] ?
                      reg1435[(4'hb):(4'ha)] : $unsigned($signed($unsigned(reg1399)))));
            end
          else
            begin
              reg1433 <= $unsigned(wire1381);
            end
          reg1437 <= $signed(((~&($unsigned(reg1413) ?
                  (~|reg1434) : (reg1417 << reg1418))) ?
              reg1394[(1'h0):(1'h0)] : $signed(($unsigned(reg1434) ^~ ((7'h40) && reg1387)))));
          reg1438 <= {$signed((~wire1381[(1'h0):(1'h0)])),
              $unsigned((reg1427[(4'he):(4'hc)] >= reg1387[(1'h0):(1'h0)]))};
          if ($unsigned((reg1435[(2'h3):(1'h1)] ?
              reg1398 : $signed(((reg1393 ?
                  reg1414 : reg1393) && $unsigned((8'ha6)))))))
            begin
              reg1439 <= wire1380;
              reg1440 <= reg1423[(3'h6):(3'h4)];
              reg1441 <= (&reg1433[(4'hc):(2'h2)]);
              reg1442 <= reg1391[(1'h0):(1'h0)];
              reg1443 <= reg1395;
            end
          else
            begin
              reg1439 <= (&reg1412[(4'h8):(3'h7)]);
              reg1440 <= reg1399[(1'h0):(1'h0)];
            end
          if ((reg1424[(4'hd):(3'h5)] + ({(^(~&reg1406))} >>> $unsigned(wire1375[(1'h0):(1'h0)]))))
            begin
              reg1444 <= (reg1443[(2'h2):(1'h0)] == $unsigned($signed((!$unsigned(reg1411)))));
              reg1445 <= $signed((($unsigned($signed((8'haa))) << ((reg1405 << (8'hb4)) ?
                  $signed(reg1397) : $signed(reg1441))) - reg1390[(3'h6):(2'h2)]));
              reg1446 <= (reg1411[(3'h4):(1'h1)] - $signed($signed($unsigned(reg1389[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg1444 <= $unsigned($unsigned((-reg1420)));
              reg1445 <= reg1445[(4'ha):(3'h5)];
              reg1446 <= (~|(~^$unsigned((~^reg1426))));
              reg1447 <= $signed(((+reg1446) ?
                  $signed(reg1443[(1'h0):(1'h0)]) : $signed({{reg1435}})));
            end
        end
      else
        begin
          reg1433 <= (7'h44);
        end
      reg1448 <= ({($signed((^~reg1423)) << reg1422[(2'h3):(2'h3)]),
              $signed(((+reg1384) && $unsigned(reg1406)))} ?
          $signed(reg1421) : (wire1375 ?
              $signed($signed((^~(8'hb7)))) : $signed((^~reg1426))));
    end
  always
    @(posedge clk) begin
      reg1449 <= (8'ha7);
      reg1450 <= reg1425[(3'h4):(2'h3)];
      if ((($signed($unsigned(reg1448[(1'h0):(1'h0)])) ?
          (^reg1439[(2'h3):(2'h2)]) : {(reg1400 ?
                  $unsigned(reg1410) : reg1400)}) >= (reg1383 && $signed(($unsigned(reg1409) ?
          $unsigned(reg1449) : (reg1393 & reg1404))))))
        begin
          if ((~&(($signed((reg1394 ? (8'hbc) : (8'hb9))) << ($signed(reg1417) ?
              $unsigned(reg1402) : (&(8'ha9)))) != $signed(((8'hb5) <= reg1435)))))
            begin
              reg1451 <= $unsigned((-reg1419));
            end
          else
            begin
              reg1451 <= reg1401;
              reg1452 <= (reg1410 - $signed(reg1394[(3'h5):(2'h3)]));
              reg1453 <= ((~|$signed($signed(reg1402))) * $unsigned(((reg1452[(5'h14):(5'h12)] << $unsigned(reg1417)) ?
                  (reg1429[(4'he):(4'hd)] ?
                      (reg1411 || reg1408) : reg1427[(5'h11):(2'h2)]) : $signed((~^reg1440)))));
            end
          reg1454 <= (^~({(^~wire1415),
              ({reg1446, reg1424} ?
                  (reg1419 | reg1433) : wire1375[(1'h0):(1'h0)])} >> ($unsigned($signed(wire1381)) ~^ $signed($unsigned(reg1423)))));
          reg1455 <= $signed((reg1406[(2'h2):(1'h0)] ?
              reg1435 : $unsigned((reg1429[(5'h10):(4'hd)] ^~ (reg1391 >= reg1403)))));
        end
      else
        begin
          reg1451 <= $signed((^((~^(reg1450 ?
              reg1449 : reg1394)) >>> ($unsigned(wire1380) <= (reg1400 ~^ wire1415)))));
        end
      reg1456 <= reg1395;
      reg1457 <= $unsigned(reg1428);
    end
  assign wire1458 = reg1390[(3'h7):(2'h3)];
  always
    @(posedge clk) begin
      reg1459 <= $signed((+(~wire1378)));
      if ($signed($signed({$signed(reg1459[(1'h0):(1'h0)])})))
        begin
          reg1460 <= ((((8'ha7) ? $signed($signed((8'hb9))) : (~(~^reg1403))) ?
                  wire1416 : reg1454[(4'h8):(4'h8)]) ?
              wire1458[(5'h14):(5'h13)] : ($signed($unsigned((reg1405 >= reg1420))) ?
                  $signed($unsigned(wire1375[(2'h3):(1'h1)])) : ($signed((~|reg1411)) & $unsigned((^~(8'hb1))))));
          reg1461 <= (!($signed(((wire1380 ?
                  reg1453 : reg1384) <= reg1418[(4'h8):(3'h5)])) ?
              (^~(^~(+reg1441))) : (reg1443 & reg1443)));
          if (($unsigned($unsigned(reg1382[(1'h0):(1'h0)])) ?
              reg1432[(4'hb):(3'h4)] : reg1410))
            begin
              reg1462 <= ((reg1419[(4'hc):(4'ha)] ?
                      ($unsigned($signed(reg1461)) ?
                          ((7'h42) - (reg1411 > reg1402)) : wire1415) : $unsigned($signed({(8'ha6),
                          reg1460}))) ?
                  (!(reg1388 || (((8'h9d) ? wire1458 : reg1398) ?
                      $unsigned(reg1421) : reg1383[(4'h8):(3'h7)]))) : (reg1385 >= $unsigned($signed((&reg1423)))));
              reg1463 <= {{((~&{reg1402}) + {(~&reg1418), $signed(reg1438)})},
                  $unsigned(($unsigned($signed(reg1396)) >> reg1411[(1'h1):(1'h0)]))};
            end
          else
            begin
              reg1462 <= ($unsigned(reg1408) ?
                  (8'had) : (reg1455 ^~ wire1381[(1'h1):(1'h1)]));
              reg1463 <= $unsigned({({(reg1447 ^~ reg1389),
                      $signed(reg1421)} && reg1451),
                  {{reg1406[(3'h6):(3'h5)], $signed(reg1423)}}});
              reg1464 <= $unsigned($signed($unsigned(wire1458)));
            end
          reg1465 <= reg1423;
          reg1466 <= reg1385;
        end
      else
        begin
          reg1460 <= (~&$signed((((reg1447 ? reg1392 : reg1463) ?
              (reg1421 ? reg1399 : wire1415) : (reg1454 ?
                  (8'hb8) : reg1382)) <<< $unsigned((reg1427 - reg1411)))));
          reg1461 <= (^{$signed({(+reg1399), $signed(reg1430)}), reg1429});
          if ($signed($signed(($unsigned((^reg1450)) & ((-reg1404) ?
              $signed(reg1412) : $unsigned((8'hba)))))))
            begin
              reg1462 <= $unsigned(((^wire1416) << $signed(reg1393[(3'h4):(1'h1)])));
              reg1463 <= $signed({(((wire1378 ?
                      (8'hbf) : reg1396) ^~ (reg1452 >= reg1448)) + $unsigned($signed(reg1447)))});
              reg1464 <= {(($unsigned($signed(reg1441)) ?
                          $unsigned($signed(wire1380)) : $unsigned((reg1404 < reg1396))) ?
                      reg1427[(4'hb):(2'h2)] : (reg1434[(4'hb):(3'h6)] - ((reg1456 + reg1442) ?
                          (reg1426 >= wire1380) : reg1386[(4'h8):(4'h8)]))),
                  reg1388[(1'h1):(1'h0)]};
              reg1465 <= reg1445;
            end
          else
            begin
              reg1462 <= $signed(($unsigned((8'hac)) ?
                  {{((8'hbd) || reg1443)}} : (reg1402[(4'ha):(4'h8)] ?
                      $unsigned($unsigned(reg1385)) : (-(+(8'hb5))))));
              reg1463 <= $signed($signed($unsigned($signed((reg1421 || (7'h44))))));
              reg1464 <= $unsigned($signed($unsigned($signed(((8'hb5) ?
                  reg1394 : reg1465)))));
            end
          reg1466 <= (+reg1433);
        end
      if (((-(+(~reg1429))) >= wire1380[(1'h1):(1'h0)]))
        begin
          if (reg1420[(3'h6):(1'h1)])
            begin
              reg1467 <= reg1459[(4'hb):(2'h3)];
              reg1468 <= ((~^reg1424) ^~ $unsigned({((7'h44) << $unsigned((8'haa)))}));
            end
          else
            begin
              reg1467 <= reg1399[(3'h6):(3'h4)];
              reg1468 <= {reg1394, $signed($unsigned(reg1435))};
              reg1469 <= reg1394;
            end
          if ((wire1378[(4'ha):(3'h6)] ?
              {(({reg1403} <<< reg1423[(3'h4):(2'h3)]) >= (reg1459[(4'h8):(2'h2)] ?
                      $signed(reg1403) : reg1465)),
                  $signed($signed({reg1434}))} : ($signed((|reg1436)) ?
                  $signed($unsigned((reg1449 ?
                      wire1378 : reg1456))) : (8'h9c))))
            begin
              reg1470 <= (reg1466[(2'h2):(1'h1)] * (reg1386 >>> (~|{$signed(reg1453),
                  $unsigned(reg1393)})));
            end
          else
            begin
              reg1470 <= ((~|(reg1461 ?
                  ($unsigned(reg1450) ?
                      reg1433[(3'h5):(1'h0)] : (&reg1424)) : (~^(+reg1464)))) << $unsigned($signed($signed(((8'h9c) >>> reg1413)))));
              reg1471 <= (-(+$signed((|(reg1419 < reg1457)))));
              reg1472 <= {$unsigned(reg1439),
                  {reg1410[(4'h9):(2'h2)], reg1448}};
              reg1473 <= $unsigned(($unsigned($unsigned(reg1457)) != {$signed({reg1438}),
                  ({reg1388} ? $signed(reg1385) : (reg1437 != reg1394))}));
              reg1474 <= (~^$signed((((!reg1473) == (wire1376 | reg1459)) ?
                  (reg1465[(3'h4):(1'h0)] + $unsigned(reg1453)) : (~^{reg1429,
                      reg1405}))));
            end
          reg1475 <= ({$signed(((reg1436 ^ reg1462) ?
                      {reg1459} : (~reg1424)))} ?
              (^~reg1447[(2'h2):(1'h0)]) : ($signed(((-wire1377) ?
                      $signed(reg1383) : wire1381)) ?
                  (((reg1413 ? reg1395 : reg1401) ? (~|reg1390) : {(8'ha2)}) ?
                      $signed((+(7'h43))) : (wire1379 ?
                          {reg1417} : $unsigned((7'h40)))) : {(~{(8'hba),
                          reg1384}),
                      (((8'hb4) ? reg1390 : reg1389) | ((8'haa) ?
                          reg1399 : (8'hbf)))}));
        end
      else
        begin
          if (($signed((8'hb1)) ?
              (reg1407[(4'h8):(1'h1)] > (+$signed(reg1396))) : $unsigned((reg1410 ?
                  $signed(reg1437) : {$unsigned(reg1391)}))))
            begin
              reg1467 <= $unsigned((reg1404[(1'h0):(1'h0)] || (({reg1389} >= (reg1402 ?
                  reg1410 : reg1455)) || (~(-reg1417)))));
              reg1468 <= $signed({reg1420[(4'h8):(2'h3)]});
              reg1469 <= {reg1473, (reg1473[(3'h5):(3'h4)] && reg1387)};
              reg1470 <= reg1393;
              reg1471 <= (-((reg1389 ?
                      $signed((-reg1391)) : $signed((reg1462 < reg1409))) ?
                  (((-reg1436) ^ (|reg1457)) >> {(reg1469 <= reg1442)}) : reg1420[(3'h4):(2'h3)]));
            end
          else
            begin
              reg1467 <= reg1390[(1'h0):(1'h0)];
              reg1468 <= {(^{((reg1423 ^~ reg1403) << reg1452),
                      reg1452[(4'hd):(1'h0)]}),
                  $signed($signed(($unsigned(wire1415) ?
                      (reg1435 & (8'hbb)) : $unsigned(reg1422))))};
              reg1469 <= $unsigned($signed(wire1376[(2'h2):(1'h0)]));
            end
          if ($signed(reg1472[(3'h6):(3'h4)]))
            begin
              reg1472 <= (~^$unsigned(wire1379[(1'h0):(1'h0)]));
              reg1473 <= {{(({reg1453} ? reg1459 : reg1472[(3'h5):(1'h1)]) ?
                          (^reg1461) : $unsigned(reg1399))}};
            end
          else
            begin
              reg1472 <= $unsigned($unsigned(wire1378[(2'h2):(1'h0)]));
              reg1473 <= (~|reg1461);
              reg1474 <= {wire1377,
                  ((reg1429[(3'h5):(1'h0)] ?
                      $signed($signed((7'h42))) : reg1467) + $signed(($unsigned(reg1406) ?
                      {wire1377, reg1447} : (^~reg1396))))};
              reg1475 <= (~^{((8'h9d) ?
                      (reg1391[(2'h3):(1'h0)] > $signed(reg1425)) : $unsigned(((8'hb4) >> reg1422)))});
              reg1476 <= ({$signed($signed((~&wire1415))),
                  $unsigned(($signed(reg1404) ?
                      (~&reg1419) : reg1420[(4'he):(1'h0)]))} || $unsigned(reg1386));
            end
          reg1477 <= (reg1476[(1'h0):(1'h0)] >> ($signed(wire1378) ?
              (({reg1384, reg1391} << reg1405) ?
                  (8'hbd) : ($signed(reg1451) ?
                      (^~reg1430) : $unsigned((8'ha6)))) : ($unsigned({wire1379,
                  reg1403}) << {$unsigned((8'hbe))})));
        end
      reg1478 <= $signed($signed(($unsigned((reg1433 ?
          reg1447 : reg1471)) << ((|reg1473) ? $signed(wire1378) : reg1387))));
    end
  assign wire1479 = (8'hbd);
  assign wire1480 = reg1459[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg1481 <= ((8'ha0) != {($unsigned((-(8'ha2))) >>> (&$signed(reg1455))),
          $signed(reg1448)});
      reg1482 <= $signed($signed(((-$unsigned(reg1481)) < (^reg1446))));
      if ((8'hb5))
        begin
          if (reg1382[(3'h5):(1'h0)])
            begin
              reg1483 <= (-$signed($signed(reg1443)));
              reg1484 <= reg1432;
            end
          else
            begin
              reg1483 <= (~&((~^(~$signed(reg1477))) - (($signed(reg1410) ?
                  {reg1475} : (reg1404 | reg1472)) >> reg1395[(5'h11):(3'h7)])));
              reg1484 <= $unsigned((~|($signed({reg1477}) ?
                  ($unsigned(reg1402) >> (reg1426 ?
                      reg1383 : reg1448)) : (reg1397 ?
                      $signed(reg1404) : ((8'hac) ? reg1451 : wire1479)))));
            end
          if (reg1447[(1'h1):(1'h1)])
            begin
              reg1485 <= (reg1409 * $unsigned(($signed(reg1475) ?
                  reg1447[(1'h0):(1'h0)] : (~|(reg1474 ? reg1473 : reg1421)))));
              reg1486 <= (-reg1419);
            end
          else
            begin
              reg1485 <= $unsigned(wire1416);
              reg1486 <= ($unsigned((reg1408[(4'ha):(1'h1)] ?
                      reg1423 : (reg1413[(2'h3):(2'h3)] || (reg1389 * reg1440)))) ?
                  ({{$unsigned(reg1433), $unsigned(reg1452)}} ?
                      wire1415 : {$signed($unsigned(reg1457))}) : reg1394);
              reg1487 <= wire1379;
            end
        end
      else
        begin
          if ($signed(reg1389[(1'h1):(1'h0)]))
            begin
              reg1483 <= (~|wire1480);
            end
          else
            begin
              reg1483 <= (~reg1455[(2'h3):(2'h2)]);
              reg1484 <= (^~(|($signed((reg1383 ?
                  reg1470 : reg1387)) == ($unsigned(reg1386) ?
                  reg1456 : (^~reg1436)))));
              reg1485 <= $signed(reg1428);
              reg1486 <= (($signed({(~&reg1413), reg1435}) ?
                  $unsigned(reg1429) : $signed((&wire1379[(2'h3):(2'h2)]))) & $signed((~^($signed(reg1411) != (reg1410 * reg1487)))));
            end
        end
      if ($unsigned(reg1414))
        begin
          reg1488 <= reg1431;
          reg1489 <= {(reg1451 ?
                  (reg1469 ?
                      wire1479 : ($unsigned((8'haa)) || ((8'had) ^ reg1476))) : $unsigned(reg1470[(4'ha):(1'h1)]))};
          reg1490 <= $unsigned(reg1435[(2'h3):(2'h2)]);
        end
      else
        begin
          if ($unsigned((reg1488[(2'h3):(1'h1)] || reg1436)))
            begin
              reg1488 <= reg1388;
              reg1489 <= reg1414;
              reg1490 <= reg1438;
            end
          else
            begin
              reg1488 <= $signed((7'h40));
            end
          reg1491 <= (~reg1432);
        end
    end
  assign wire1492 = (~$unsigned($signed((&((8'hb5) ? (8'hbb) : reg1403)))));
  assign wire1493 = ($unsigned(reg1413) ?
                        (reg1490 ?
                            $unsigned({(~|(8'had))}) : (reg1477[(3'h5):(2'h2)] ?
                                reg1482[(2'h3):(2'h2)] : reg1408[(3'h4):(1'h1)])) : $unsigned((|$unsigned(reg1406[(1'h1):(1'h0)]))));
  assign wire1494 = (^~(8'hae));
  always
    @(posedge clk) begin
      reg1495 <= reg1433;
      reg1496 <= $unsigned($unsigned(((+(-reg1461)) ?
          (reg1468[(1'h0):(1'h0)] ?
              $unsigned(reg1488) : $signed((8'hbd))) : ((reg1438 ?
              reg1452 : reg1406) >> (reg1439 && reg1418)))));
      reg1497 <= (($signed(((reg1437 ? reg1426 : reg1406) ?
                  $signed(reg1401) : (reg1429 ? reg1399 : reg1464))) ?
              wire1377 : (((8'hbe) ?
                  wire1480 : reg1434[(1'h0):(1'h0)]) > reg1387[(1'h1):(1'h1)])) ?
          reg1447[(4'h9):(4'h8)] : $unsigned((|$unsigned(reg1484[(5'h10):(4'hf)]))));
    end
  assign wire1498 = (reg1439[(3'h4):(1'h1)] ? reg1385[(4'h9):(1'h1)] : reg1462);
  assign wire1499 = $unsigned({(|reg1486[(1'h1):(1'h1)]),
                        (reg1444[(1'h1):(1'h1)] ~^ {wire1376[(1'h1):(1'h1)]})});
  assign wire1500 = $signed(reg1452);
  assign wire1501 = (-(!reg1434));
  assign wire1502 = $signed(reg1382);
  assign wire1503 = $unsigned($signed((reg1452 != (+reg1467[(3'h7):(1'h0)]))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1333
#( parameter param1370 = (|(({(8'ha3), ((8'ha6) ? (7'h41) : (8'hb6))} && ((^(7'h41)) & ((8'ha1) ? (8'h9d) : (8'hab)))) ? {(((8'hbe) >= (8'hbf)) ? (~(8'hbf)) : {(8'ha6)})} : (^(((7'h41) ? (8'hb1) : (8'h9d)) | ((8'hbc) ? (7'h41) : (8'h9d))))))
, parameter param1371 = param1370 )
(y, clk, wire1337, wire1336, wire1335, wire1334);
  output wire [(32'h15f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire1337;
  input wire signed [(3'h6):(1'h0)] wire1336;
  input wire signed [(5'h11):(1'h0)] wire1335;
  input wire signed [(4'h8):(1'h0)] wire1334;
  reg [(5'h11):(1'h0)] reg1369 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1368 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire1367;
  wire [(3'h4):(1'h0)] wire1366;
  wire signed [(5'h11):(1'h0)] wire1365;
  reg signed [(3'h5):(1'h0)] reg1364 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1363 = (1'h0);
  reg [(2'h2):(1'h0)] reg1362 = (1'h0);
  reg [(2'h3):(1'h0)] reg1361 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1360 = (1'h0);
  reg [(4'h9):(1'h0)] reg1359 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1358 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1357 = (1'h0);
  reg [(5'h12):(1'h0)] reg1356 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1355 = (1'h0);
  reg [(4'hd):(1'h0)] reg1354 = (1'h0);
  reg [(5'h11):(1'h0)] reg1353 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1352 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1351 = (1'h0);
  reg [(4'he):(1'h0)] reg1350 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1349 = (1'h0);
  reg [(4'ha):(1'h0)] reg1348 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1347 = (1'h0);
  reg [(5'h14):(1'h0)] reg1346 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1345 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire1344;
  reg [(4'ha):(1'h0)] reg1343 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1342 = (1'h0);
  reg [(3'h6):(1'h0)] reg1341 = (1'h0);
  reg [(3'h6):(1'h0)] reg1340 = (1'h0);
  reg [(4'hf):(1'h0)] reg1339 = (1'h0);
  reg [(4'hb):(1'h0)] reg1338 = (1'h0);
  assign y = {reg1369,
                 reg1368,
                 wire1367,
                 wire1366,
                 wire1365,
                 reg1364,
                 reg1363,
                 reg1362,
                 reg1361,
                 reg1360,
                 reg1359,
                 reg1358,
                 reg1357,
                 reg1356,
                 reg1355,
                 reg1354,
                 reg1353,
                 reg1352,
                 reg1351,
                 reg1350,
                 reg1349,
                 reg1348,
                 reg1347,
                 reg1346,
                 reg1345,
                 wire1344,
                 reg1343,
                 reg1342,
                 reg1341,
                 reg1340,
                 reg1339,
                 reg1338,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (((^~wire1335) ?
          wire1335 : (^($signed($signed(wire1336)) ?
              $unsigned((wire1337 == wire1335)) : wire1334[(3'h5):(2'h3)]))))
        begin
          reg1338 <= wire1335[(4'hc):(1'h1)];
        end
      else
        begin
          if (wire1335)
            begin
              reg1338 <= ((({(|wire1336)} & {reg1338[(4'ha):(4'ha)]}) << (!wire1334)) ?
                  wire1334 : $unsigned({$unsigned(wire1334[(2'h3):(2'h2)])}));
              reg1339 <= wire1335[(5'h11):(4'hb)];
              reg1340 <= {wire1334[(4'h8):(4'h8)]};
              reg1341 <= (wire1334[(1'h0):(1'h0)] ?
                  wire1334 : $signed($signed(($unsigned(wire1335) ^ (reg1338 ^~ wire1337)))));
              reg1342 <= ({$signed((((8'hae) && (8'hb9)) ?
                          (-reg1341) : $unsigned(reg1338))),
                      reg1339[(3'h4):(2'h2)]} ?
                  ($unsigned((&$unsigned(reg1340))) > (+(8'haa))) : $signed((($unsigned(reg1339) ?
                          $signed(wire1336) : (reg1341 <<< reg1340)) ?
                      (8'hb9) : $unsigned({reg1341}))));
            end
          else
            begin
              reg1338 <= $signed($signed((wire1336[(1'h1):(1'h1)] ?
                  reg1339 : $unsigned({reg1342, wire1334}))));
              reg1339 <= $unsigned(reg1338);
              reg1340 <= reg1342;
              reg1341 <= wire1335[(3'h5):(1'h1)];
              reg1342 <= $unsigned((reg1342 ?
                  wire1337 : reg1341[(2'h2):(1'h0)]));
            end
          reg1343 <= (~reg1339[(4'ha):(3'h5)]);
        end
    end
  assign wire1344 = (~$signed($signed(((wire1334 ? wire1337 : wire1335) ?
                        (reg1342 ~^ reg1342) : (~reg1342)))));
  always
    @(posedge clk) begin
      if ($unsigned((8'ha2)))
        begin
          reg1345 <= reg1339[(4'hf):(4'hd)];
          reg1346 <= ($unsigned(wire1336) & reg1338[(3'h4):(3'h4)]);
          reg1347 <= ($signed((~&((~|reg1338) ?
              $unsigned(reg1346) : (reg1340 ?
                  reg1340 : reg1342)))) | wire1337[(2'h2):(2'h2)]);
          reg1348 <= $unsigned((reg1338[(4'h8):(3'h7)] >> ($unsigned($unsigned(reg1342)) ?
              (wire1337[(2'h3):(1'h1)] ^~ wire1335[(1'h0):(1'h0)]) : $signed({wire1344,
                  reg1345}))));
          if (reg1345[(1'h0):(1'h0)])
            begin
              reg1349 <= (-(wire1335[(4'hd):(3'h7)] >> ($signed(reg1348[(4'h8):(3'h5)]) ?
                  $unsigned($unsigned((8'hb5))) : {reg1340[(3'h6):(2'h3)],
                      $signed((8'hb2))})));
              reg1350 <= (~&(!$unsigned(reg1340)));
            end
          else
            begin
              reg1349 <= ({(($signed(reg1348) ?
                              (!wire1337) : reg1350[(4'hb):(3'h5)]) ?
                          {wire1336,
                              reg1343[(4'h8):(1'h0)]} : $signed(reg1346))} ?
                  (~$signed(reg1347[(3'h6):(1'h0)])) : {{$unsigned(reg1346[(4'h8):(3'h7)])},
                      (reg1346[(2'h3):(2'h3)] + ($signed(wire1335) ?
                          (8'had) : $signed(reg1349)))});
              reg1350 <= $signed((wire1337 ?
                  (8'hb5) : (~^$unsigned(reg1343[(4'ha):(1'h0)]))));
              reg1351 <= {($unsigned($unsigned({wire1334,
                      reg1345})) < $unsigned(reg1345)),
                  reg1350};
              reg1352 <= reg1349[(3'h7):(1'h1)];
            end
        end
      else
        begin
          reg1345 <= wire1344[(2'h2):(1'h0)];
          reg1346 <= (($signed($unsigned((reg1343 ? reg1342 : reg1341))) ?
              reg1352[(2'h2):(1'h1)] : $signed(reg1352[(2'h2):(1'h1)])) | reg1348[(3'h7):(3'h5)]);
        end
      reg1353 <= $unsigned((reg1346[(4'hd):(3'h6)] ?
          ($unsigned(reg1339) ?
              (&reg1340[(2'h2):(1'h0)]) : (~|reg1347[(3'h5):(1'h0)])) : (wire1344 ?
              (!$unsigned(reg1352)) : ((reg1343 >= reg1348) >= (reg1346 | wire1344)))));
      reg1354 <= reg1339;
    end
  always
    @(posedge clk) begin
      reg1355 <= ({(reg1346 <= $unsigned($unsigned(reg1348))),
              $unsigned((~$unsigned(wire1336)))} ?
          (reg1349 ?
              (wire1344[(3'h4):(2'h2)] ?
                  {(reg1340 & reg1340)} : reg1338[(3'h4):(3'h4)]) : (~&wire1336[(3'h6):(2'h3)])) : (!reg1340));
      if ({reg1345[(1'h1):(1'h0)], reg1345})
        begin
          if ((-reg1346))
            begin
              reg1356 <= (~&(!$unsigned(reg1341[(3'h5):(3'h5)])));
              reg1357 <= $signed($signed(reg1348[(4'ha):(3'h7)]));
              reg1358 <= (+{reg1350});
            end
          else
            begin
              reg1356 <= $unsigned(((reg1352[(2'h2):(1'h0)] ?
                      reg1346 : (-reg1350)) ?
                  reg1340[(2'h2):(2'h2)] : reg1356[(1'h1):(1'h0)]));
              reg1357 <= reg1351[(2'h3):(2'h2)];
              reg1358 <= wire1336[(2'h3):(2'h2)];
              reg1359 <= $unsigned({(|wire1336)});
            end
          if ($unsigned($signed((~&(|$signed((8'hab)))))))
            begin
              reg1360 <= $unsigned((!reg1359[(2'h2):(1'h0)]));
              reg1361 <= reg1356[(4'ha):(1'h1)];
              reg1362 <= reg1350;
              reg1363 <= (|reg1343[(1'h0):(1'h0)]);
            end
          else
            begin
              reg1360 <= ((!(|$signed((8'ha1)))) > (+{reg1345[(1'h0):(1'h0)]}));
              reg1361 <= wire1336;
              reg1362 <= (reg1363 || $unsigned(($unsigned(((8'hb8) < wire1344)) == (~^reg1341))));
            end
        end
      else
        begin
          reg1356 <= $signed($signed($signed(reg1362)));
          reg1357 <= (({$signed((reg1345 ? reg1355 : reg1350))} ?
                  (&reg1345) : $signed({$unsigned(reg1348),
                      $unsigned(reg1345)})) ?
              reg1351 : $unsigned((reg1351[(4'ha):(1'h1)] ?
                  wire1337 : ((reg1363 + reg1349) ~^ $signed(reg1356)))));
        end
      reg1364 <= (~&{(+reg1361), (7'h43)});
    end
  assign wire1365 = {reg1350[(3'h7):(2'h2)],
                        ((reg1348[(4'ha):(1'h1)] + ($signed(reg1364) ^ (wire1337 * reg1358))) * $signed(reg1357[(4'hc):(4'h9)]))};
  assign wire1366 = ((~(~&((|wire1334) ?
                        reg1362[(1'h1):(1'h1)] : $unsigned(reg1357)))) ^ (($unsigned($signed((8'hbb))) ~^ (^$signed(reg1346))) ?
                        wire1365[(4'hc):(3'h5)] : ((((8'ha0) ?
                            reg1358 : reg1346) ^~ (reg1363 ?
                            reg1350 : reg1359)) ~^ ((~|reg1342) < (&(8'ha2))))));
  assign wire1367 = (!{(!(reg1350 | (8'ha4)))});
  always
    @(posedge clk) begin
      reg1368 <= (+(+({$unsigned(reg1360),
          (wire1365 ? wire1366 : reg1352)} - (+(wire1337 == (8'hbb))))));
      reg1369 <= $unsigned((~(^~($signed(reg1356) ?
          $unsigned(wire1335) : ((8'ha7) ? reg1357 : reg1338)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1743
#( parameter param1768 = (&(8'ha0))
, parameter param1769 = (((((param1768 ^ (8'hbe)) ? {(8'haf), param1768} : (|param1768)) ~^ ((-param1768) <<< {param1768, (8'haf)})) ? param1768 : param1768) ? ((((param1768 ? param1768 : param1768) | ((7'h41) ? param1768 : param1768)) >> (param1768 > (param1768 | param1768))) ? (|((param1768 ? param1768 : param1768) * (param1768 | (8'hbe)))) : (^~(!{param1768}))) : (((^(|param1768)) ? (param1768 ? (!param1768) : ((7'h40) ? param1768 : param1768)) : {param1768, (param1768 > (8'ha8))}) <<< (8'hb5))) )
(y, clk, wire1748, wire1747, wire1746, wire1745, wire1744);
  output wire [(32'hea):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire1748;
  input wire [(4'hd):(1'h0)] wire1747;
  input wire [(4'hb):(1'h0)] wire1746;
  input wire signed [(5'h14):(1'h0)] wire1745;
  input wire [(4'hc):(1'h0)] wire1744;
  reg signed [(4'h8):(1'h0)] reg1767 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1766 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1765 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1764 = (1'h0);
  reg [(3'h4):(1'h0)] reg1763 = (1'h0);
  reg [(5'h15):(1'h0)] reg1762 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1761 = (1'h0);
  reg [(4'hf):(1'h0)] reg1760 = (1'h0);
  reg [(3'h5):(1'h0)] reg1759 = (1'h0);
  reg [(3'h4):(1'h0)] reg1758 = (1'h0);
  wire [(3'h5):(1'h0)] wire1757;
  wire signed [(4'hf):(1'h0)] wire1756;
  wire signed [(5'h11):(1'h0)] wire1755;
  wire [(4'hc):(1'h0)] wire1754;
  wire [(4'hf):(1'h0)] wire1753;
  wire signed [(3'h7):(1'h0)] wire1752;
  wire signed [(4'h9):(1'h0)] wire1751;
  wire [(5'h14):(1'h0)] wire1750;
  wire signed [(5'h12):(1'h0)] wire1749;
  assign y = {reg1767,
                 reg1766,
                 reg1765,
                 reg1764,
                 reg1763,
                 reg1762,
                 reg1761,
                 reg1760,
                 reg1759,
                 reg1758,
                 wire1757,
                 wire1756,
                 wire1755,
                 wire1754,
                 wire1753,
                 wire1752,
                 wire1751,
                 wire1750,
                 wire1749,
                 (1'h0)};
  assign wire1749 = wire1744[(4'hc):(4'hc)];
  assign wire1750 = wire1749[(1'h0):(1'h0)];
  assign wire1751 = {((wire1749 <= $signed($signed(wire1747))) >= (((|(8'hbf)) >>> $signed(wire1744)) ?
                            $unsigned((wire1746 ?
                                wire1749 : wire1750)) : ($unsigned((8'ha3)) ?
                                wire1748 : wire1750))),
                        wire1746};
  assign wire1752 = wire1748;
  assign wire1753 = $unsigned($signed({(^$signed(wire1748))}));
  assign wire1754 = (wire1745[(3'h4):(3'h4)] ?
                        wire1750[(3'h7):(3'h7)] : $signed((!$signed((wire1750 ?
                            wire1752 : (8'hb3))))));
  assign wire1755 = (wire1751[(3'h4):(1'h0)] <<< wire1749[(1'h1):(1'h1)]);
  assign wire1756 = wire1744[(4'ha):(2'h3)];
  assign wire1757 = (wire1756 ?
                        $signed(($signed((wire1746 != wire1751)) || ($signed(wire1749) ?
                            wire1751[(3'h4):(1'h1)] : $signed(wire1751)))) : $signed($unsigned($unsigned(wire1750[(3'h5):(3'h5)]))));
  always
    @(posedge clk) begin
      if (((($signed($unsigned(wire1751)) ?
          (wire1747 * (wire1757 ?
              wire1748 : wire1756)) : (~|(-wire1751))) ^ wire1756) >> wire1753))
        begin
          if ((&(wire1749[(2'h2):(1'h0)] <= (8'h9c))))
            begin
              reg1758 <= wire1750[(4'he):(4'ha)];
              reg1759 <= wire1746[(2'h2):(1'h1)];
              reg1760 <= wire1748[(1'h1):(1'h1)];
            end
          else
            begin
              reg1758 <= wire1746;
              reg1759 <= $unsigned(((!wire1749) ? wire1747 : wire1753));
              reg1760 <= (wire1757[(3'h5):(1'h1)] - wire1755);
              reg1761 <= $unsigned(($unsigned((!$signed(wire1744))) && wire1753));
              reg1762 <= {(|$signed({wire1747[(4'h8):(2'h3)]}))};
            end
          if (wire1746[(4'hb):(4'h8)])
            begin
              reg1763 <= $unsigned((wire1757[(1'h1):(1'h0)] ?
                  (((reg1760 ? reg1759 : wire1757) ?
                          $signed(wire1745) : (wire1751 ^~ (8'hac))) ?
                      (wire1749 * (reg1758 ?
                          (8'had) : wire1748)) : $unsigned((wire1747 ?
                          wire1750 : wire1748))) : ($signed((wire1750 && reg1761)) != (^~(wire1757 ?
                      (8'hb6) : reg1761)))));
            end
          else
            begin
              reg1763 <= reg1762[(4'hd):(4'ha)];
            end
          reg1764 <= (^(8'hb7));
          reg1765 <= (8'hb1);
          reg1766 <= reg1764;
        end
      else
        begin
          reg1758 <= ((~$unsigned((+{reg1762}))) ?
              (~wire1749) : ((wire1748[(2'h2):(2'h2)] ?
                  $signed({wire1747}) : (-(wire1750 | reg1759))) < (((reg1762 << wire1756) & $signed(wire1751)) < wire1755[(2'h3):(1'h1)])));
          reg1759 <= wire1754[(1'h1):(1'h1)];
        end
      reg1767 <= $signed((&$signed(($signed((8'ha7)) ?
          $unsigned(wire1744) : (-reg1763)))));
    end
endmodule