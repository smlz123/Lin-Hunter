(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param566 = (8'ha4), parameter param567 = (8'haf))
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h270):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire0;
  input wire [(3'h5):(1'h0)] wire1;
  input wire signed [(5'h13):(1'h0)] wire2;
  input wire signed [(3'h6):(1'h0)] wire3;
  input wire [(5'h11):(1'h0)] wire4;
  wire signed [(3'h4):(1'h0)] wire565;
  reg [(5'h13):(1'h0)] reg564 = (1'h0);
  reg [(2'h2):(1'h0)] reg563 = (1'h0);
  reg [(5'h11):(1'h0)] reg562 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg561 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg560 = (1'h0);
  reg [(2'h3):(1'h0)] reg559 = (1'h0);
  reg [(2'h3):(1'h0)] reg558 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg557 = (1'h0);
  reg [(5'h15):(1'h0)] forvar556 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg555 = (1'h0);
  reg [(3'h4):(1'h0)] reg554 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg553 = (1'h0);
  reg [(2'h2):(1'h0)] reg552 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg551 = (1'h0);
  reg [(5'h13):(1'h0)] reg550 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg549 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg548 = (1'h0);
  wire [(4'hf):(1'h0)] wire5;
  reg signed [(4'ha):(1'h0)] reg6 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar7 = (1'h0);
  reg [(4'hb):(1'h0)] reg8 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg9 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg10 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg11 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar12 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg14 = (1'h0);
  reg [(4'h8):(1'h0)] reg15 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg16 = (1'h0);
  reg [(4'hb):(1'h0)] forvar17 = (1'h0);
  reg [(4'hb):(1'h0)] reg18 = (1'h0);
  reg [(4'hb):(1'h0)] reg19 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg20 = (1'h0);
  reg [(4'ha):(1'h0)] reg21 = (1'h0);
  reg [(4'ha):(1'h0)] reg22 = (1'h0);
  wire [(4'h9):(1'h0)] wire23;
  wire signed [(3'h6):(1'h0)] wire24;
  reg signed [(4'ha):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg26 = (1'h0);
  reg [(3'h7):(1'h0)] forvar27 = (1'h0);
  reg [(4'hb):(1'h0)] reg28 = (1'h0);
  reg [(5'h11):(1'h0)] reg29 = (1'h0);
  reg [(4'hd):(1'h0)] reg30 = (1'h0);
  wire [(4'h9):(1'h0)] wire31;
  wire signed [(4'hf):(1'h0)] wire32;
  wire [(5'h15):(1'h0)] wire33;
  wire signed [(3'h5):(1'h0)] wire34;
  reg signed [(3'h6):(1'h0)] reg35 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar36 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg37 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg38 = (1'h0);
  wire [(5'h11):(1'h0)] wire39;
  wire signed [(4'hf):(1'h0)] wire546;
  assign y = {wire565,
                 reg564,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 reg558,
                 reg557,
                 forvar556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 reg549,
                 reg548,
                 wire5,
                 reg6,
                 forvar7,
                 reg8,
                 reg9,
                 reg10,
                 reg11,
                 forvar12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 forvar17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 wire23,
                 wire24,
                 reg25,
                 reg26,
                 forvar27,
                 reg28,
                 reg29,
                 reg30,
                 wire31,
                 wire32,
                 wire33,
                 wire34,
                 reg35,
                 forvar36,
                 reg37,
                 reg38,
                 wire39,
                 wire546,
                 (1'h0)};
  assign wire5 = $unsigned(wire1[(3'h5):(3'h5)]);
  always
    @(posedge clk) begin
      reg6 <= ($unsigned(((wire5 ^ (wire4 >= wire2)) ?
          wire5 : wire0)) >>> (((((8'hbd) ? wire0 : (8'haf)) ?
                  wire1 : (-wire3)) ?
              wire5[(1'h1):(1'h0)] : $signed((~|wire1))) ?
          (({wire5} << $unsigned((8'hb9))) ?
              wire1 : $signed(wire3)) : (^$signed((wire4 ? wire5 : wire1)))));
      for (forvar7 = (1'h0); (forvar7 < (2'h2)); forvar7 = (forvar7 + (1'h1)))
        begin
          reg8 = wire4;
        end
      reg9 <= wire2[(5'h10):(3'h5)];
      reg10 = $signed((~&$unsigned(wire1)));
    end
  always
    @(posedge clk) begin
      reg11 = $unsigned((8'h9c));
      for (forvar12 = (1'h0); (forvar12 < (2'h2)); forvar12 = (forvar12 + (1'h1)))
        begin
          reg13 = (!reg8);
          reg14 <= ((7'h42) != (8'ha3));
          reg15 <= {$unsigned($unsigned(reg6))};
          reg16 <= reg8;
          for (forvar17 = (1'h0); (forvar17 < (1'h1)); forvar17 = (forvar17 + (1'h1)))
            begin
              reg18 <= ($signed({$signed((reg11 ? wire2 : wire0)),
                      $signed(forvar17)}) ?
                  forvar17 : wire5[(1'h0):(1'h0)]);
              reg19 = (+(!$unsigned(wire1)));
            end
        end
      reg20 <= (($signed((-{reg6, reg8})) ^ $signed($unsigned((forvar17 ?
          (8'hb8) : forvar17)))) && $signed({({reg19} ?
              wire5 : $unsigned(wire4))}));
    end
  always
    @(posedge clk) begin
      reg21 <= ($unsigned((~|{$signed(reg19), forvar7})) ?
          $unsigned((reg18 ? (8'hbc) : {(^~reg19)})) : (((wire1 ?
                  $unsigned(reg13) : (~(8'hac))) << (~{(8'hb7), reg15})) ?
              $unsigned(((wire4 >> (7'h41)) < reg19[(4'h9):(3'h4)])) : {$unsigned($signed(forvar12))}));
      reg22 = $unsigned(wire5[(4'hf):(4'ha)]);
    end
  assign wire23 = forvar17[(3'h4):(2'h2)];
  assign wire24 = reg13;
  always
    @(posedge clk) begin
      reg25 <= $unsigned($signed((-(-$signed(reg13)))));
      reg26 = {$signed(reg11)};
      for (forvar27 = (1'h0); (forvar27 < (2'h3)); forvar27 = (forvar27 + (1'h1)))
        begin
          reg28 <= $unsigned((~&reg22[(3'h6):(3'h6)]));
          reg29 <= $unsigned(((+{$unsigned(reg20),
              (~^(8'ha8))}) || {(reg10[(3'h6):(3'h5)] >>> (reg25 ^ reg25)),
              ({reg25} ? (&reg26) : $unsigned(reg26))}));
        end
      reg30 <= $unsigned(((((forvar12 * wire2) <<< {reg16, wire0}) ?
              forvar27 : (!$signed(wire24))) ?
          $signed($unsigned(wire2)) : (wire23[(4'h8):(3'h7)] >>> $signed((^reg11)))));
    end
  assign wire31 = ((+$unsigned((~(forvar17 < wire4)))) & reg8);
  assign wire32 = $unsigned((reg18[(1'h1):(1'h1)] ?
                      ((((8'h9c) <<< wire3) ~^ $unsigned((8'hb0))) ?
                          $unsigned((wire24 ?
                              reg29 : reg26)) : $signed(wire4[(1'h0):(1'h0)])) : reg20[(1'h1):(1'h1)]));
  assign wire33 = reg20;
  assign wire34 = $unsigned(forvar12);
  always
    @(posedge clk) begin
      reg35 <= $signed($signed($unsigned($unsigned({forvar17}))));
      for (forvar36 = (1'h0); (forvar36 < (3'h4)); forvar36 = (forvar36 + (1'h1)))
        begin
          reg37 <= $signed(wire31[(4'h8):(3'h6)]);
          reg38 <= reg35;
        end
    end
  assign wire39 = ($unsigned((($signed(reg38) ?
                          $signed(reg14) : reg13[(1'h0):(1'h0)]) >= (+(reg29 ?
                          reg15 : forvar12)))) ?
                      (reg20 | reg29[(2'h3):(1'h0)]) : (~|(-$unsigned($signed((8'hb1))))));
  module40 modinst547 (.wire41(reg26), .clk(clk), .wire43(wire4), .wire44(reg37), .y(wire546), .wire42(forvar36), .wire45(reg25));
  always
    @(posedge clk) begin
      reg548 <= reg6[(1'h0):(1'h0)];
      reg549 <= (($signed((!wire34)) ?
          $unsigned($signed(reg35)) : reg38[(4'ha):(1'h1)]) << reg8);
      reg550 <= $signed((~&reg26));
      reg551 <= ((-wire4) ?
          $signed({(-$signed(reg548))}) : {wire34,
              {wire4[(4'he):(3'h7)], (8'hb7)}});
    end
  always
    @(posedge clk) begin
      reg552 <= ($signed($unsigned(((wire0 ? reg29 : reg8) ?
          (reg16 + wire0) : {forvar12}))) < (^(8'hb8)));
      reg553 <= forvar7[(5'h11):(3'h7)];
      reg554 <= (wire3[(2'h3):(1'h0)] << ($signed((8'hb5)) | (reg551[(3'h4):(1'h0)] ?
          ((~^(8'ha7)) ? $unsigned((8'hbc)) : (reg548 >> (8'hb7))) : wire3)));
      reg555 = $signed(reg548);
      for (forvar556 = (1'h0); (forvar556 < (1'h0)); forvar556 = (forvar556 + (1'h1)))
        begin
          reg557 = reg25[(4'h9):(1'h0)];
          reg558 = ($signed((~reg16)) ?
              ((&reg554[(2'h2):(1'h0)]) ?
                  wire4 : reg30[(1'h1):(1'h0)]) : {wire33[(2'h2):(1'h1)],
                  ((^~reg28) ? reg550 : reg550[(3'h4):(3'h4)])});
          reg559 <= ($unsigned(wire3[(3'h6):(3'h6)]) - ((8'hba) ?
              $unsigned(((reg8 | wire1) ?
                  {reg25} : wire34[(1'h0):(1'h0)])) : (((^~reg551) ?
                      (wire34 + (8'haa)) : $unsigned(wire31)) ?
                  $unsigned((reg35 ?
                      wire23 : (8'ha7))) : $unsigned($signed((8'hb7))))));
        end
    end
  always
    @(posedge clk) begin
      reg560 <= ((&reg38) <= ({(|$unsigned(forvar12))} >= $unsigned($signed(wire31[(1'h0):(1'h0)]))));
    end
  always
    @(posedge clk) begin
      reg561 <= $signed((^((~{reg552, wire3}) ? reg548 : (8'ha3))));
    end
  always
    @(posedge clk) begin
      reg562 <= $signed({(($unsigned(reg559) ?
              (8'hb9) : (^~reg30)) | $unsigned(forvar27[(3'h7):(1'h0)]))});
    end
  always
    @(posedge clk) begin
      reg563 <= (reg37 | $unsigned(wire23[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg564 <= (!$unsigned((forvar12[(4'hc):(2'h3)] ?
          (wire2 | wire4[(4'ha):(3'h5)]) : (|{wire1, reg554}))));
    end
  assign wire565 = ($signed($signed($signed($unsigned(reg10)))) - ($signed(((&wire24) - (wire33 >= wire23))) ?
                       forvar12[(3'h7):(1'h1)] : $signed(wire39)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module40
#( parameter param544 = (((~|((~(8'hbb)) >>> ((8'hb9) ? (8'h9f) : (7'h40)))) * ((((8'hbe) != (8'hb7)) ? ((8'ha6) > (8'ha7)) : ((8'ha3) >>> (7'h42))) >>> (~|((8'hab) <<< (7'h40))))) ? (((((8'hab) ? (8'ha2) : (7'h41)) ^ ((8'ha5) ? (8'hb2) : (8'ha3))) ? (8'h9e) : (((8'ha6) ~^ (8'ha4)) ? (-(8'hb3)) : ((8'hbc) ? (8'h9d) : (8'h9d)))) >> ((((8'hb4) ? (8'ha4) : (8'ha2)) ? (^(7'h40)) : ((8'hbe) ? (8'ha3) : (7'h40))) || ((+(8'ha1)) ? ((8'ha3) ? (8'ha1) : (8'hb0)) : ((8'ha4) ^~ (8'hae))))) : (((~(^(8'ha1))) >= (|((8'ha8) ? (7'h44) : (8'hbc)))) ~^ (^{(~^(8'hbc)), ((8'h9f) ? (8'had) : (8'hb3))})))
, parameter param545 = ((param544 ? {((param544 ? param544 : param544) ? (^~param544) : param544)} : {param544, (((8'hbe) ? (7'h40) : (8'hb5)) > (param544 <<< param544))}) ? (({((7'h41) ? param544 : param544)} > (param544 ? (param544 ? param544 : param544) : (+param544))) <<< (((param544 <= (8'hb0)) << (param544 ? param544 : param544)) ? param544 : ((~^param544) <<< (param544 ? param544 : param544)))) : ((((param544 ? param544 : param544) * param544) >>> param544) ? (({param544} ? (!param544) : (8'hba)) & ((~&(8'hbb)) ? (param544 >>> param544) : (~&param544))) : ((!param544) > (^param544)))) )
(y, clk, wire41, wire42, wire43, wire44, wire45);
  output wire [(32'h476):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire41;
  input wire signed [(5'h14):(1'h0)] wire42;
  input wire signed [(5'h11):(1'h0)] wire43;
  input wire [(5'h13):(1'h0)] wire44;
  input wire [(4'ha):(1'h0)] wire45;
  wire [(4'h9):(1'h0)] wire543;
  wire [(2'h2):(1'h0)] wire542;
  reg signed [(5'h10):(1'h0)] reg541 = (1'h0);
  reg [(5'h11):(1'h0)] reg540 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg539 = (1'h0);
  reg [(5'h10):(1'h0)] reg538 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar537 = (1'h0);
  reg [(4'hd):(1'h0)] reg536 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg535 = (1'h0);
  reg [(4'hf):(1'h0)] forvar534 = (1'h0);
  reg [(4'hf):(1'h0)] reg533 = (1'h0);
  reg [(5'h10):(1'h0)] reg532 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg531 = (1'h0);
  reg [(4'hf):(1'h0)] reg530 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg529 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg528 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar527 = (1'h0);
  reg [(4'hf):(1'h0)] forvar526 = (1'h0);
  reg [(4'hf):(1'h0)] reg516 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg525 = (1'h0);
  reg [(4'hb):(1'h0)] reg524 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar523 = (1'h0);
  reg [(3'h5):(1'h0)] reg522 = (1'h0);
  reg [(3'h6):(1'h0)] reg521 = (1'h0);
  reg [(4'hf):(1'h0)] reg520 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg519 = (1'h0);
  reg [(4'ha):(1'h0)] reg518 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg517 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar516 = (1'h0);
  reg [(3'h7):(1'h0)] reg515 = (1'h0);
  reg [(4'hf):(1'h0)] reg514 = (1'h0);
  reg [(2'h2):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg47 = (1'h0);
  reg [(2'h3):(1'h0)] reg48 = (1'h0);
  reg [(2'h3):(1'h0)] reg49 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire50;
  reg [(3'h5):(1'h0)] reg51 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar52 = (1'h0);
  reg [(5'h14):(1'h0)] reg53 = (1'h0);
  reg [(4'h8):(1'h0)] reg54 = (1'h0);
  reg [(4'hb):(1'h0)] reg55 = (1'h0);
  reg [(4'hd):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg57 = (1'h0);
  reg [(2'h2):(1'h0)] forvar58 = (1'h0);
  reg [(4'hb):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg60 = (1'h0);
  reg [(3'h7):(1'h0)] reg61 = (1'h0);
  wire [(2'h3):(1'h0)] wire62;
  reg signed [(4'hd):(1'h0)] reg63 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar64 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg65 = (1'h0);
  reg [(4'hc):(1'h0)] reg66 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg67 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire68;
  wire signed [(4'he):(1'h0)] wire69;
  wire signed [(4'h8):(1'h0)] wire70;
  reg signed [(5'h15):(1'h0)] reg71 = (1'h0);
  reg [(4'h9):(1'h0)] reg72 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg73 = (1'h0);
  wire [(5'h13):(1'h0)] wire74;
  reg signed [(3'h7):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar76 = (1'h0);
  reg [(5'h12):(1'h0)] reg77 = (1'h0);
  reg [(3'h5):(1'h0)] reg78 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar79 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg80 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg81 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar82 = (1'h0);
  reg [(4'hb):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg84 = (1'h0);
  reg [(5'h15):(1'h0)] reg85 = (1'h0);
  reg [(5'h14):(1'h0)] reg86 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar87 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg88 = (1'h0);
  reg [(4'h9):(1'h0)] reg89 = (1'h0);
  reg [(4'hb):(1'h0)] reg90 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar91 = (1'h0);
  reg [(4'h8):(1'h0)] reg92 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg93 = (1'h0);
  reg [(4'h9):(1'h0)] reg94 = (1'h0);
  reg [(4'ha):(1'h0)] reg95 = (1'h0);
  reg [(5'h11):(1'h0)] reg96 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar97 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg98 = (1'h0);
  reg [(5'h14):(1'h0)] reg99 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg100 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg101 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar103 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg104 = (1'h0);
  reg [(4'hd):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg106 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg108 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire512;
  assign y = {wire543,
                 wire542,
                 reg541,
                 reg540,
                 reg539,
                 reg538,
                 forvar537,
                 reg536,
                 reg535,
                 forvar534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 forvar527,
                 forvar526,
                 reg516,
                 reg525,
                 reg524,
                 forvar523,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 reg517,
                 forvar516,
                 reg515,
                 reg514,
                 reg46,
                 reg47,
                 reg48,
                 reg49,
                 wire50,
                 reg51,
                 forvar52,
                 reg53,
                 reg54,
                 reg55,
                 reg56,
                 reg57,
                 forvar58,
                 reg59,
                 reg60,
                 reg61,
                 wire62,
                 reg63,
                 forvar64,
                 reg65,
                 reg66,
                 reg67,
                 wire68,
                 wire69,
                 wire70,
                 reg71,
                 reg72,
                 reg73,
                 wire74,
                 reg75,
                 forvar76,
                 reg77,
                 reg78,
                 forvar79,
                 reg80,
                 reg76,
                 reg81,
                 forvar82,
                 reg83,
                 reg84,
                 reg85,
                 reg86,
                 forvar87,
                 reg88,
                 reg89,
                 reg90,
                 forvar91,
                 reg92,
                 reg93,
                 reg94,
                 reg95,
                 reg96,
                 forvar97,
                 reg98,
                 reg99,
                 reg100,
                 reg101,
                 reg102,
                 forvar103,
                 reg104,
                 reg105,
                 reg106,
                 reg107,
                 reg108,
                 wire512,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg46 <= wire44;
      reg47 = ({(&{wire44[(4'h9):(4'h9)]}), $signed({wire43})} ?
          (wire41[(1'h1):(1'h0)] ?
              $signed((!$signed(wire41))) : wire41[(2'h2):(1'h0)]) : (((wire43[(4'he):(4'he)] && $unsigned(wire43)) ?
                  ({reg46} ?
                      $signed(reg46) : {wire45, (8'haa)}) : (^~(~(8'ha9)))) ?
              (|wire43[(1'h1):(1'h1)]) : (wire41 ?
                  (~&(wire45 ? reg46 : wire43)) : ((wire43 ?
                      wire43 : (8'hab)) >> wire45))));
      reg48 <= (~|(((reg46[(1'h0):(1'h0)] ?
              ((7'h40) | (8'hb1)) : reg47) && (~^$unsigned((8'haa)))) ?
          $signed((~&$unsigned(wire41))) : (^(wire41 ?
              reg47[(4'he):(4'ha)] : wire43[(4'hf):(3'h4)]))));
      reg49 = (((~&$unsigned((&(8'hb0)))) ?
              wire42 : (reg46[(1'h1):(1'h0)] | wire44[(3'h6):(1'h0)])) ?
          (!reg46[(2'h2):(1'h0)]) : (!$unsigned(($unsigned((7'h42)) ?
              reg48[(2'h2):(1'h1)] : $unsigned(wire43)))));
    end
  assign wire50 = wire41;
  always
    @(posedge clk) begin
      reg51 = {(~(wire42 ? wire43 : $signed((reg48 || (7'h41)))))};
      for (forvar52 = (1'h0); (forvar52 < (1'h1)); forvar52 = (forvar52 + (1'h1)))
        begin
          reg53 <= {$signed($signed((reg48 ?
                  reg47[(1'h0):(1'h0)] : (wire45 & (8'haf))))),
              wire44[(3'h4):(2'h3)]};
          reg54 <= reg48;
          reg55 = $signed($signed(wire41));
        end
      reg56 <= (|($signed(wire50) <<< $signed($unsigned((reg49 | (8'hb7))))));
      reg57 <= $signed(reg48[(2'h3):(1'h0)]);
      for (forvar58 = (1'h0); (forvar58 < (1'h0)); forvar58 = (forvar58 + (1'h1)))
        begin
          reg59 = forvar52[(3'h6):(2'h2)];
          reg60 <= reg55;
          reg61 <= reg57[(3'h4):(2'h3)];
        end
    end
  assign wire62 = wire41;
  always
    @(posedge clk) begin
      reg63 = {$unsigned(wire43[(4'h8):(3'h7)])};
      for (forvar64 = (1'h0); (forvar64 < (2'h2)); forvar64 = (forvar64 + (1'h1)))
        begin
          reg65 <= $unsigned((($signed({wire42, reg57}) ?
              {{(8'hbf)}, $signed(reg60)} : ($signed(reg47) ?
                  (8'hb1) : $unsigned(reg46))) ^ (!$signed((!reg53)))));
          reg66 <= $unsigned($unsigned({$signed($unsigned(reg63))}));
        end
      reg67 = reg54;
    end
  assign wire68 = (+$unsigned((((wire45 + reg48) ? (^reg54) : reg53) ?
                      ((reg53 <<< reg56) ^ $signed(reg55)) : $signed(reg59[(4'ha):(4'h8)]))));
  assign wire69 = $unsigned($unsigned((8'hb7)));
  assign wire70 = $unsigned(wire45[(3'h6):(2'h2)]);
  always
    @(posedge clk) begin
      reg71 <= {wire41, ((8'hb3) ? wire68 : ((-$unsigned(wire68)) - reg54))};
      reg72 = reg67[(3'h6):(2'h3)];
      reg73 <= ((8'hbf) > (|$unsigned(reg48[(1'h0):(1'h0)])));
    end
  assign wire74 = wire44;
  always
    @(posedge clk) begin
      reg75 <= reg46;
      if ((8'h9f))
        begin
          for (forvar76 = (1'h0); (forvar76 < (2'h3)); forvar76 = (forvar76 + (1'h1)))
            begin
              reg77 <= $unsigned(forvar52);
            end
          reg78 <= ($signed((reg55 ? wire62 : reg77[(4'h9):(1'h0)])) >>> reg59);
          for (forvar79 = (1'h0); (forvar79 < (1'h0)); forvar79 = (forvar79 + (1'h1)))
            begin
              reg80 <= ((reg77 ?
                      reg61[(1'h1):(1'h1)] : $unsigned((~^(^~(8'hb5))))) ?
                  reg67[(3'h6):(3'h4)] : (~^($unsigned(reg56) ?
                      $signed($signed(wire69)) : ({forvar79, wire42} ?
                          $unsigned(wire41) : $unsigned(reg57)))));
            end
        end
      else
        begin
          reg76 = {(wire74[(5'h10):(4'hf)] ?
                  $signed($unsigned((~&reg55))) : ($unsigned(reg51) * ((-reg65) <<< (~&(7'h40)))))};
          reg77 <= ((+($signed({forvar64}) ?
              {$unsigned(reg60)} : ($unsigned(reg56) ?
                  $signed(reg65) : (!wire45)))) <<< reg54);
          reg78 <= ({$unsigned($signed($unsigned(reg53)))} * (((&(wire42 <= wire70)) ?
              $unsigned((reg53 ^~ reg47)) : (reg49[(1'h1):(1'h0)] ?
                  $signed(reg46) : $signed(forvar52))) - (+(+{wire42}))));
        end
      reg81 <= (~&($signed(wire74) ?
          {wire41[(2'h3):(2'h3)]} : $signed($unsigned(((8'hb4) << wire43)))));
      for (forvar82 = (1'h0); (forvar82 < (1'h1)); forvar82 = (forvar82 + (1'h1)))
        begin
          reg83 = reg48[(1'h1):(1'h0)];
          reg84 <= (reg65 ?
              $signed(reg73) : ((reg59[(3'h7):(3'h4)] >= ((8'ha1) >>> ((7'h40) >= reg75))) >> reg46[(1'h1):(1'h0)]));
          reg85 <= (-$unsigned(wire70));
          reg86 <= $signed($unsigned($signed($unsigned($signed(wire41)))));
          for (forvar87 = (1'h0); (forvar87 < (2'h2)); forvar87 = (forvar87 + (1'h1)))
            begin
              reg88 <= reg73;
              reg89 <= (reg84 >= $unsigned(($signed((wire50 ? wire50 : reg49)) ?
                  reg80[(1'h0):(1'h0)] : $signed((forvar64 <<< (8'ha0))))));
              reg90 <= reg77;
            end
        end
      for (forvar91 = (1'h0); (forvar91 < (2'h3)); forvar91 = (forvar91 + (1'h1)))
        begin
          reg92 <= reg81;
          reg93 = $unsigned($unsigned(forvar76[(5'h12):(4'hf)]));
          reg94 <= reg85[(4'hf):(4'hc)];
        end
    end
  always
    @(posedge clk) begin
      reg95 <= (~|$signed(({(reg55 * (8'hb1))} * ($signed(forvar79) << {reg78,
          reg78}))));
      reg96 <= forvar82[(3'h4):(2'h2)];
      for (forvar97 = (1'h0); (forvar97 < (2'h2)); forvar97 = (forvar97 + (1'h1)))
        begin
          reg98 <= ((!$unsigned(($unsigned(wire41) && forvar91[(2'h3):(2'h3)]))) ?
              (+(-(8'hbd))) : {reg46,
                  (wire41 + $signed((reg84 ? reg94 : reg66)))});
          reg99 <= ((!(-$signed($signed((8'hbb))))) ^ $unsigned((reg71 ?
              (8'ha5) : (|(reg75 != reg98)))));
        end
      reg100 <= {(reg65[(4'he):(3'h5)] ^~ reg72[(4'h8):(3'h6)])};
      reg101 = ((reg96 <<< ($signed((reg57 < forvar79)) <= {reg67[(2'h2):(2'h2)],
          $unsigned(reg83)})) <<< $unsigned((7'h42)));
    end
  always
    @(posedge clk) begin
      reg102 <= reg49;
      for (forvar103 = (1'h0); (forvar103 < (1'h0)); forvar103 = (forvar103 + (1'h1)))
        begin
          if (($unsigned($unsigned($signed({(8'hb7),
              (8'haf)}))) <= $signed((($signed(forvar52) ?
              $signed((8'hbb)) : (!forvar97)) > reg54[(1'h1):(1'h0)]))))
            begin
              reg104 = (({($unsigned(reg65) ~^ (forvar91 * reg78)),
                          ((wire62 ? forvar103 : reg101) ?
                              $signed((8'ha6)) : (~|reg51))} ?
                      ($signed($unsigned(reg56)) ?
                          $signed(reg100[(2'h3):(2'h2)]) : $signed(reg98[(3'h5):(2'h2)])) : (|($unsigned(wire70) ?
                          (reg95 ? forvar52 : reg59) : {reg73, reg81}))) ?
                  (($unsigned($unsigned(reg53)) < (+(8'ha8))) * (!forvar97[(3'h6):(2'h3)])) : (($unsigned($signed(reg46)) ?
                          (!$signed(reg56)) : $signed(reg102)) ?
                      $unsigned(({reg49} | $signed(forvar52))) : (($unsigned(forvar103) ?
                          forvar52[(4'hc):(4'hb)] : $unsigned(reg54)) ~^ (forvar82[(3'h7):(1'h1)] ?
                          ((8'hb6) ? wire43 : forvar103) : (^reg46)))));
              reg105 <= $unsigned(((((reg92 >> wire44) - $unsigned(reg63)) ?
                  $signed((reg72 ?
                      reg101 : reg54)) : ((!reg56) <= forvar91)) >> (+($signed(reg51) ?
                  (forvar91 ~^ reg104) : ((8'hb2) <<< reg65)))));
              reg106 <= reg92[(2'h2):(1'h1)];
            end
          else
            begin
              reg104 = (8'ha6);
              reg105 <= $unsigned(forvar64);
            end
          reg107 = reg59;
        end
      reg108 <= reg102;
    end
  module109 modinst513 (.clk(clk), .wire112(reg86), .wire111(forvar79), .wire114(wire68), .y(wire512), .wire113(reg93), .wire110(reg78));
  always
    @(posedge clk) begin
      reg514 <= (reg59 ?
          (^~$signed($unsigned($signed(reg57)))) : $unsigned(wire62[(1'h1):(1'h0)]));
      if ((~$signed($signed({wire44, $signed(reg85)}))))
        begin
          reg515 <= $signed($unsigned(reg59));
          for (forvar516 = (1'h0); (forvar516 < (2'h3)); forvar516 = (forvar516 + (1'h1)))
            begin
              reg517 <= reg515;
              reg518 = $signed(((8'haa) ^~ $unsigned(reg92[(3'h4):(2'h3)])));
              reg519 <= $unsigned(($signed({$signed(reg86)}) ?
                  $unsigned(reg59[(4'ha):(4'h9)]) : {$signed(reg96[(4'hb):(2'h3)])}));
              reg520 <= (reg56[(4'hc):(1'h0)] ? reg92 : $unsigned(reg56));
            end
          reg521 = {((wire69[(3'h4):(3'h4)] ?
                      (-$signed((8'ha7))) : ($signed(reg515) != (~&wire43))) ?
                  $unsigned(forvar64) : $signed(reg61[(3'h4):(2'h2)]))};
          reg522 <= wire62;
          for (forvar523 = (1'h0); (forvar523 < (3'h4)); forvar523 = (forvar523 + (1'h1)))
            begin
              reg524 = forvar516;
              reg525 <= reg88[(4'h8):(3'h6)];
            end
        end
      else
        begin
          reg515 = (8'ha7);
          reg516 <= (+wire512);
          reg517 <= ((|(|reg95[(3'h7):(3'h6)])) ?
              reg54[(3'h6):(3'h6)] : $signed(({wire44[(3'h7):(1'h1)]} | (!(reg73 ?
                  wire44 : reg517)))));
        end
      for (forvar526 = (1'h0); (forvar526 < (1'h0)); forvar526 = (forvar526 + (1'h1)))
        begin
          for (forvar527 = (1'h0); (forvar527 < (3'h4)); forvar527 = (forvar527 + (1'h1)))
            begin
              reg528 <= (-$signed($unsigned($signed($unsigned(wire44)))));
              reg529 <= (7'h44);
              reg530 = reg55[(4'h9):(3'h5)];
              reg531 <= forvar87[(1'h0):(1'h0)];
            end
          reg532 <= ((~&reg46) >>> ({reg65[(2'h3):(2'h3)],
                  wire45[(3'h5):(3'h5)]} ?
              reg51[(1'h1):(1'h1)] : forvar526[(4'he):(3'h6)]));
          reg533 = ((&$unsigned(reg531[(4'ha):(3'h5)])) * {reg94,
              reg48[(1'h1):(1'h1)]});
          for (forvar534 = (1'h0); (forvar534 < (3'h4)); forvar534 = (forvar534 + (1'h1)))
            begin
              reg535 <= reg107[(3'h4):(1'h1)];
            end
        end
      reg536 <= (reg51[(1'h0):(1'h0)] ?
          (reg108 ?
              reg106 : $unsigned(($signed(reg105) ?
                  (7'h40) : $unsigned(forvar82)))) : $signed($unsigned((((8'hbe) >>> reg85) > wire512[(4'h9):(4'h8)]))));
      for (forvar537 = (1'h0); (forvar537 < (2'h2)); forvar537 = (forvar537 + (1'h1)))
        begin
          reg538 = $signed(wire512);
          reg539 <= ($signed(reg94) ?
              ((-((reg72 ? reg76 : forvar82) == (forvar87 > reg57))) ?
                  $unsigned(reg531[(3'h4):(1'h0)]) : $unsigned(reg90[(2'h3):(1'h1)])) : {reg528[(3'h6):(2'h3)]});
          reg540 <= $signed($signed(reg71));
          reg541 <= ({$unsigned($signed(forvar516[(3'h4):(1'h0)]))} ?
              $signed($signed((~|$signed((7'h41))))) : {(8'h9d),
                  {((reg528 ? reg101 : reg81) ?
                          (|reg71) : (forvar523 <<< reg96)),
                      $unsigned((reg95 ? reg78 : reg85))}});
        end
    end
  assign wire542 = (($signed(((8'hb6) != ((8'had) >> reg59))) ?
                           $unsigned($unsigned($signed((8'had)))) : (~^$signed((reg72 && (8'hb6))))) ?
                       $signed({wire69[(4'hd):(2'h2)]}) : $signed(($signed($unsigned(reg46)) == ((reg67 ^~ reg530) ?
                           ((8'ha2) < reg517) : (~reg83)))));
  assign wire543 = {wire44[(5'h13):(3'h7)],
                       ($signed($unsigned((~&forvar537))) && $unsigned((~^$unsigned(reg102))))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module109
#( parameter param511 = ((~|(~^{((7'h43) || (8'hbe))})) ? ((|{(8'hb6)}) ? {(((8'hba) > (8'h9c)) ? ((8'hb7) ^ (8'ha7)) : ((8'ha8) ? (8'haf) : (8'ha3))), (((8'hb5) > (8'hb4)) ? (~(7'h42)) : {(8'hbc)})} : ((+((8'hae) ? (8'had) : (8'ha0))) ? ({(8'hb7)} ? (7'h44) : {(7'h43)}) : (((8'ha2) * (8'ha0)) < (~^(8'hae))))) : ({(+(~&(8'hb3))), (((8'hb3) ? (8'hb8) : (8'hbc)) ? (+(8'hbe)) : {(8'h9e)})} ? ((((8'hb7) && (8'hba)) ? (8'ha2) : ((7'h42) && (8'hbe))) ? (((8'hac) ? (8'hb9) : (8'hba)) <= (~|(8'h9c))) : (((8'hba) || (8'hb5)) ? ((8'hb7) > (8'ha9)) : ((8'hb8) ? (7'h42) : (8'hb9)))) : (!(((8'hae) | (7'h41)) < (~(8'hb8)))))) )
(y, clk, wire110, wire111, wire112, wire113, wire114);
  output wire [(32'h15c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire110;
  input wire signed [(5'h13):(1'h0)] wire111;
  input wire signed [(5'h14):(1'h0)] wire112;
  input wire [(4'ha):(1'h0)] wire113;
  input wire [(4'hb):(1'h0)] wire114;
  reg [(5'h10):(1'h0)] reg510 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire509;
  reg [(5'h14):(1'h0)] reg508 = (1'h0);
  reg [(4'he):(1'h0)] reg507 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg506 = (1'h0);
  wire [(3'h5):(1'h0)] wire115;
  wire signed [(3'h6):(1'h0)] wire116;
  reg signed [(4'h8):(1'h0)] forvar117 = (1'h0);
  reg [(5'h13):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar119 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg120 = (1'h0);
  reg [(5'h11):(1'h0)] reg121 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg122 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg124 = (1'h0);
  reg [(4'h8):(1'h0)] reg125 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg126 = (1'h0);
  reg [(5'h11):(1'h0)] reg127 = (1'h0);
  reg [(5'h10):(1'h0)] reg128 = (1'h0);
  reg [(4'hb):(1'h0)] reg129 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg130 = (1'h0);
  reg [(3'h4):(1'h0)] reg131 = (1'h0);
  reg [(4'ha):(1'h0)] reg132 = (1'h0);
  reg signed [(4'he):(1'h0)] reg133 = (1'h0);
  reg [(5'h10):(1'h0)] reg134 = (1'h0);
  reg [(5'h14):(1'h0)] reg135 = (1'h0);
  wire [(3'h6):(1'h0)] wire504;
  assign y = {reg510,
                 wire509,
                 reg508,
                 reg507,
                 reg506,
                 wire115,
                 wire116,
                 forvar117,
                 reg118,
                 forvar119,
                 reg120,
                 reg121,
                 reg122,
                 reg123,
                 reg124,
                 reg125,
                 reg126,
                 reg127,
                 reg128,
                 reg129,
                 reg130,
                 reg131,
                 reg132,
                 reg133,
                 reg134,
                 reg135,
                 wire504,
                 (1'h0)};
  assign wire115 = wire112[(4'h8):(3'h4)];
  assign wire116 = ($unsigned($unsigned(wire110[(2'h2):(1'h0)])) ?
                       {($signed({(7'h43), wire112}) && $unsigned((wire111 ?
                               wire114 : (8'h9c)))),
                           ($signed((-wire113)) >>> $unsigned((~wire113)))} : ({$unsigned(((8'ha2) ?
                                   wire111 : wire111)),
                               wire111[(3'h7):(3'h5)]} ?
                           ((^~$unsigned(wire110)) ?
                               (wire112[(4'ha):(4'h9)] ?
                                   $unsigned(wire115) : (-wire114)) : (~$signed(wire112))) : $unsigned(wire110[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      for (forvar117 = (1'h0); (forvar117 < (3'h4)); forvar117 = (forvar117 + (1'h1)))
        begin
          reg118 = (((($signed(wire114) >= (wire111 || (8'hb1))) ?
              ($signed(forvar117) ?
                  $unsigned((7'h41)) : {wire112}) : $signed((wire116 | wire111))) ~^ {$unsigned(((8'ha4) ?
                  wire116 : wire111))}) > (^{forvar117[(1'h0):(1'h0)],
              $signed($signed(wire116))}));
          for (forvar119 = (1'h0); (forvar119 < (2'h3)); forvar119 = (forvar119 + (1'h1)))
            begin
              reg120 <= (~|((((wire111 >> wire115) | $signed(wire112)) > $unsigned($unsigned(wire110))) && wire112[(3'h4):(2'h2)]));
              reg121 <= wire110;
              reg122 <= ((~^(forvar119[(3'h6):(3'h6)] ?
                      wire111 : $signed($unsigned(wire116)))) ?
                  reg118 : (+$signed(((reg121 ?
                      reg118 : reg121) ^ $unsigned((8'ha2))))));
            end
          reg123 <= (-wire110[(2'h2):(1'h0)]);
          reg124 <= $signed($unsigned($unsigned($signed(forvar117[(4'h8):(2'h2)]))));
          reg125 <= ((^(^~($signed(reg122) ?
                  (wire110 ? reg122 : reg124) : (!wire114)))) ?
              (8'h9e) : $signed($unsigned($signed($signed(wire113)))));
        end
      reg126 <= (wire113 ?
          (reg124 << $unsigned(wire115)) : (^(((wire111 && reg120) || {wire116}) ?
              ((|reg118) == wire116[(1'h1):(1'h0)]) : wire112[(4'ha):(3'h7)])));
      reg127 = {$signed($unsigned(((reg124 ? reg118 : wire113) <<< (wire112 ?
              reg123 : wire112)))),
          reg123};
      reg128 <= $signed($unsigned($unsigned($unsigned(reg126))));
      reg129 = ({$unsigned($unsigned((reg118 || reg118))),
          ({{reg118, forvar117},
              wire115} & $unsigned($signed(reg124)))} + (8'hac));
    end
  always
    @(posedge clk) begin
      reg130 <= $unsigned((wire114[(3'h6):(1'h1)] ?
          ((reg126 ?
              (forvar119 >> reg128) : reg122[(4'hf):(4'he)]) >= $signed(wire114)) : reg124));
    end
  always
    @(posedge clk) begin
      reg131 = (^~(reg122 >>> $signed($signed($signed(reg127)))));
      reg132 <= reg126;
      reg133 <= ($signed((^reg125)) ?
          ((^~$signed((wire115 ? forvar119 : reg126))) == $signed((^(wire115 ?
              forvar119 : forvar119)))) : $unsigned(($signed((reg128 ~^ reg132)) ?
              $signed((^reg124)) : ($unsigned(wire116) ^ $signed(forvar117)))));
      reg134 <= $signed((^~reg118));
      reg135 <= wire111[(3'h7):(2'h2)];
    end
  module136 modinst505 (.y(wire504), .wire138(reg120), .clk(clk), .wire140(reg132), .wire137(reg118), .wire139(reg130), .wire141(reg124));
  always
    @(posedge clk) begin
      reg506 <= reg132[(4'h9):(3'h5)];
    end
  always
    @(posedge clk) begin
      reg507 <= {$unsigned(($unsigned(wire113[(4'h8):(3'h5)]) ?
              ((reg126 ?
                  reg120 : reg122) ^~ reg118) : $signed((wire115 >= (8'hba)))))};
    end
  always
    @(posedge clk) begin
      reg508 <= reg123;
    end
  assign wire509 = $unsigned((~&(reg125 ?
                       forvar117[(3'h4):(3'h4)] : ((wire112 ?
                           reg125 : reg506) && $signed((8'hb1))))));
  always
    @(posedge clk) begin
      reg510 <= ((8'hbb) - reg508[(3'h6):(2'h3)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module136
#( parameter param503 = {(!(({(8'ha3), (8'ha6)} ? ((8'ha3) >>> (8'hb2)) : ((8'ha8) || (8'hbc))) || (((8'hbb) ? (8'hbd) : (8'haa)) ? ((8'h9d) ? (8'hbb) : (8'hb1)) : {(8'ha2), (8'hb0)}))), (((~(8'ha4)) ? (-((8'ha9) ? (8'hac) : (8'ha4))) : (~(8'ha8))) >>> {{((8'hb3) ^ (7'h43))}, ({(8'hb3)} < (|(8'hb1)))})} )
(y, clk, wire141, wire140, wire139, wire138, wire137);
  output wire [(32'h23a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire141;
  input wire [(4'ha):(1'h0)] wire140;
  input wire signed [(4'he):(1'h0)] wire139;
  input wire [(5'h10):(1'h0)] wire138;
  input wire signed [(5'h13):(1'h0)] wire137;
  reg signed [(2'h3):(1'h0)] reg502 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg501 = (1'h0);
  reg [(3'h5):(1'h0)] reg500 = (1'h0);
  reg [(3'h5):(1'h0)] reg499 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg498 = (1'h0);
  wire [(4'he):(1'h0)] wire497;
  wire [(4'he):(1'h0)] wire496;
  reg signed [(4'hd):(1'h0)] reg495 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg494 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg493 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg492 = (1'h0);
  reg [(5'h10):(1'h0)] reg491 = (1'h0);
  reg [(5'h14):(1'h0)] reg490 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar489 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire488;
  wire [(3'h4):(1'h0)] wire486;
  reg [(3'h5):(1'h0)] reg266 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg265 = (1'h0);
  reg [(4'hb):(1'h0)] reg264 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar262 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg261 = (1'h0);
  reg [(4'hf):(1'h0)] reg260 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire259;
  wire signed [(3'h7):(1'h0)] wire183;
  wire signed [(3'h4):(1'h0)] wire185;
  wire [(4'h9):(1'h0)] wire186;
  wire signed [(3'h7):(1'h0)] wire187;
  reg signed [(4'hf):(1'h0)] reg188 = (1'h0);
  reg [(3'h6):(1'h0)] reg189 = (1'h0);
  reg [(5'h11):(1'h0)] reg190 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg193 = (1'h0);
  reg [(2'h3):(1'h0)] reg194 = (1'h0);
  reg [(4'he):(1'h0)] reg195 = (1'h0);
  reg [(3'h7):(1'h0)] forvar196 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar197 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg198 = (1'h0);
  reg [(4'h9):(1'h0)] reg199 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg200 = (1'h0);
  reg signed [(4'he):(1'h0)] reg201 = (1'h0);
  reg [(5'h10):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg204 = (1'h0);
  reg [(5'h11):(1'h0)] reg205 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg206 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire207;
  reg signed [(4'he):(1'h0)] reg208 = (1'h0);
  wire [(4'hc):(1'h0)] wire209;
  wire signed [(3'h4):(1'h0)] wire257;
  assign y = {reg502,
                 reg501,
                 reg500,
                 reg499,
                 reg498,
                 wire497,
                 wire496,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 reg491,
                 reg490,
                 forvar489,
                 wire488,
                 wire486,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 forvar262,
                 reg261,
                 reg260,
                 wire259,
                 wire183,
                 wire185,
                 wire186,
                 wire187,
                 reg188,
                 reg189,
                 reg190,
                 reg191,
                 reg192,
                 reg193,
                 reg194,
                 reg195,
                 forvar196,
                 forvar197,
                 reg198,
                 reg199,
                 reg200,
                 reg201,
                 reg202,
                 reg203,
                 reg204,
                 reg205,
                 reg206,
                 wire207,
                 reg208,
                 wire209,
                 wire257,
                 (1'h0)};
  module142 modinst184 (.wire147(wire138), .wire143(wire139), .wire146(wire140), .wire144(wire137), .y(wire183), .wire145(wire141), .clk(clk));
  assign wire185 = $signed((-(^~{wire138[(4'hd):(3'h5)]})));
  assign wire186 = $unsigned(((wire185 ?
                       ($signed(wire185) ?
                           (wire138 >= wire140) : wire137) : ((wire141 ?
                               (7'h43) : wire140) ?
                           (wire140 > wire137) : wire185)) < (wire141[(1'h0):(1'h0)] ?
                       $unsigned((wire139 > wire185)) : ((wire141 >> wire183) ?
                           $signed(wire183) : (~wire141)))));
  assign wire187 = (^wire183);
  always
    @(posedge clk) begin
      reg188 <= $signed((wire141 ?
          $signed($signed((~|wire187))) : (((8'ha8) ?
              wire187 : $unsigned(wire141)) != ($unsigned(wire186) && wire141[(3'h7):(3'h7)]))));
      reg189 <= $unsigned(wire137);
    end
  always
    @(posedge clk) begin
      reg190 <= $signed((~^wire140));
      reg191 <= $signed(wire183);
      reg192 <= $unsigned(wire186[(2'h2):(1'h1)]);
      reg193 = (~(8'haa));
    end
  always
    @(posedge clk) begin
      reg194 <= (reg188 >> reg191);
      reg195 <= $unsigned(reg190);
      for (forvar196 = (1'h0); (forvar196 < (3'h4)); forvar196 = (forvar196 + (1'h1)))
        begin
          for (forvar197 = (1'h0); (forvar197 < (1'h0)); forvar197 = (forvar197 + (1'h1)))
            begin
              reg198 <= ($unsigned($unsigned($unsigned(((8'hb1) < (8'hbb))))) ?
                  $unsigned({(~^reg195)}) : reg195);
              reg199 <= (^{(wire137 ?
                      reg198[(3'h5):(1'h1)] : wire141[(1'h0):(1'h0)]),
                  $signed(wire141)});
              reg200 = (forvar197[(1'h1):(1'h0)] ?
                  ($signed(reg191[(4'h9):(1'h1)]) | reg193) : ((&$unsigned($unsigned(reg189))) ?
                      wire138[(4'hf):(4'ha)] : $unsigned(reg193[(2'h3):(2'h3)])));
              reg201 <= (reg192 ? reg193[(2'h3):(2'h2)] : reg191);
            end
          reg202 <= wire137;
          reg203 = (reg202[(1'h1):(1'h1)] ?
              $unsigned((wire183 ?
                  {(^reg189),
                      wire139[(2'h2):(1'h1)]} : $signed({reg189}))) : reg190[(3'h4):(2'h2)]);
        end
      reg204 <= $signed({wire140[(4'h9):(2'h3)],
          $signed((^~(forvar197 ? reg192 : wire137)))});
    end
  always
    @(posedge clk) begin
      reg205 <= (wire137[(4'h9):(1'h0)] ?
          ($signed((reg191[(1'h1):(1'h0)] || (reg194 ?
              wire141 : forvar197))) >> (~(+(reg198 ?
              reg192 : reg203)))) : (($unsigned((reg198 ~^ (8'h9f))) == ((wire183 | (8'hbd)) != (&wire139))) ?
              ((wire183 != forvar197[(1'h0):(1'h0)]) ?
                  forvar196[(3'h6):(1'h0)] : wire186[(3'h4):(2'h2)]) : (~&wire137)));
      reg206 <= ((($signed($unsigned(reg192)) != reg189) * $unsigned(reg198[(2'h3):(2'h2)])) ?
          (reg194[(1'h0):(1'h0)] ?
              {((wire183 << reg198) ? reg199 : $signed(reg189)),
                  reg202} : $unsigned((((8'ha8) >> reg204) >> (wire187 <= wire185)))) : (({$unsigned((8'hac)),
              $unsigned(forvar197)} != reg202) & ($signed((wire138 ?
                  reg199 : forvar197)) ?
              ((~&wire185) || reg194[(1'h1):(1'h1)]) : (reg195[(2'h3):(2'h3)] > (wire185 <= (8'h9e))))));
    end
  assign wire207 = (wire185[(1'h0):(1'h0)] ?
                       $unsigned(reg189[(1'h0):(1'h0)]) : (^~$unsigned(forvar196)));
  always
    @(posedge clk) begin
      reg208 = (+reg194);
    end
  assign wire209 = $unsigned((~$signed({reg203, (wire183 & (8'hab))})));
  module210 modinst258 (.y(wire257), .wire211(wire141), .wire215(reg208), .wire212(forvar197), .wire214(reg200), .clk(clk), .wire213(reg193));
  assign wire259 = (-wire137);
  always
    @(posedge clk) begin
      reg260 <= reg205[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg261 = (-(^({$signed(forvar196)} > $signed((wire183 ^ reg260)))));
      for (forvar262 = (1'h0); (forvar262 < (2'h2)); forvar262 = (forvar262 + (1'h1)))
        begin
          reg263 <= $unsigned($signed($signed({wire141})));
          reg264 = (~({((wire183 ? reg208 : wire138) && (reg192 ?
                  wire209 : reg202))} <= ($unsigned((reg202 | reg201)) | (reg199 ?
              (wire139 ? (7'h41) : reg195) : forvar196))));
          reg265 = reg206;
        end
      reg266 = reg198;
    end
  module267 modinst487 (wire486, clk, reg263, reg205, reg265, wire141);
  assign wire488 = wire141[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      for (forvar489 = (1'h0); (forvar489 < (2'h3)); forvar489 = (forvar489 + (1'h1)))
        begin
          reg490 <= (|$unsigned(((7'h41) ?
              {(forvar196 | (7'h40))} : $signed((8'ha1)))));
          reg491 = ((&((~reg266) ?
              ({reg204, (8'ha0)} ?
                  (reg265 ?
                      (8'ha5) : reg266) : (^wire141)) : forvar262[(1'h0):(1'h0)])) | (~&(-$signed(reg188[(4'ha):(1'h0)]))));
          reg492 <= $signed(($signed(reg192[(1'h1):(1'h0)]) ?
              $unsigned(($unsigned(wire183) ^~ ((8'hba) ?
                  wire139 : wire140))) : (+((forvar196 >>> reg195) >= $signed(reg195)))));
        end
      reg493 = (forvar196 < $unsigned($unsigned(wire140)));
      reg494 = $unsigned($signed(reg192));
      reg495 = ((reg191[(2'h3):(1'h1)] && ($unsigned($unsigned(wire257)) ~^ $unsigned($signed((8'ha5))))) ?
          ((&$signed(forvar197)) ?
              (~^{$unsigned(forvar197)}) : $unsigned(reg494[(4'hb):(3'h7)])) : ($signed(((8'h9d) ?
                  (~^reg190) : (wire259 < reg491))) ?
              $unsigned(wire488[(4'h8):(3'h6)]) : ((+(8'ha2)) ?
                  (~|wire207[(4'h9):(2'h3)]) : wire137[(3'h4):(1'h0)])));
    end
  assign wire496 = ((~|(($unsigned(wire140) <= $unsigned(forvar489)) ?
                       ($signed(reg493) ?
                           (reg205 != reg208) : wire183) : (~|$signed(forvar489)))) - wire139);
  assign wire497 = (~^reg261[(2'h2):(1'h1)]);
  always
    @(posedge clk) begin
      reg498 <= ($signed(($signed($unsigned(wire138)) ?
          wire497[(3'h5):(2'h3)] : $signed((reg203 ?
              (8'hb2) : wire141)))) & ((8'hb2) && (-((wire207 - reg205) | ((8'hac) == wire183)))));
      reg499 <= $signed($signed($signed({forvar262, $unsigned((8'hb7))})));
      reg500 <= $unsigned($unsigned(reg493[(3'h4):(2'h3)]));
      reg501 <= {$unsigned(reg498[(2'h3):(1'h0)])};
      reg502 <= wire488[(5'h13):(3'h7)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module267  (y, clk, wire271, wire270, wire269, wire268);
  output wire [(32'h1dc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire271;
  input wire [(5'h11):(1'h0)] wire270;
  input wire [(5'h12):(1'h0)] wire269;
  input wire signed [(4'hb):(1'h0)] wire268;
  reg [(4'hf):(1'h0)] reg485 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar484 = (1'h0);
  reg [(3'h5):(1'h0)] reg483 = (1'h0);
  reg [(5'h11):(1'h0)] reg482 = (1'h0);
  reg [(4'ha):(1'h0)] reg481 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg480 = (1'h0);
  reg [(5'h10):(1'h0)] forvar479 = (1'h0);
  reg [(4'he):(1'h0)] reg478 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg477 = (1'h0);
  reg [(5'h10):(1'h0)] reg476 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg475 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg474 = (1'h0);
  reg [(5'h10):(1'h0)] forvar473 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg472 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar471 = (1'h0);
  reg [(4'h8):(1'h0)] reg470 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg469 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire468;
  wire [(4'hc):(1'h0)] wire467;
  wire signed [(5'h15):(1'h0)] wire465;
  reg [(5'h11):(1'h0)] reg362 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire361;
  wire [(5'h10):(1'h0)] wire360;
  reg signed [(2'h2):(1'h0)] reg359 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire358;
  reg [(4'he):(1'h0)] reg357 = (1'h0);
  reg [(4'hd):(1'h0)] reg356 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg355 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg354 = (1'h0);
  reg [(4'he):(1'h0)] reg353 = (1'h0);
  reg [(5'h12):(1'h0)] reg352 = (1'h0);
  reg [(5'h14):(1'h0)] reg351 = (1'h0);
  reg [(4'hf):(1'h0)] reg350 = (1'h0);
  wire [(3'h4):(1'h0)] wire349;
  wire signed [(4'hc):(1'h0)] wire348;
  wire [(4'hd):(1'h0)] wire347;
  reg [(4'hf):(1'h0)] reg346 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg345 = (1'h0);
  wire [(3'h7):(1'h0)] wire343;
  wire [(4'hb):(1'h0)] wire273;
  wire signed [(4'hb):(1'h0)] wire272;
  assign y = {reg485,
                 forvar484,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 forvar479,
                 reg478,
                 reg477,
                 reg476,
                 reg475,
                 reg474,
                 forvar473,
                 reg472,
                 forvar471,
                 reg470,
                 reg469,
                 wire468,
                 wire467,
                 wire465,
                 reg362,
                 wire361,
                 wire360,
                 reg359,
                 wire358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 reg350,
                 wire349,
                 wire348,
                 wire347,
                 reg346,
                 reg345,
                 wire343,
                 wire273,
                 wire272,
                 (1'h0)};
  assign wire272 = wire269;
  assign wire273 = $signed(($signed($signed($signed(wire269))) >> wire271));
  module274 modinst344 (.wire275(wire270), .y(wire343), .clk(clk), .wire277(wire273), .wire276(wire268), .wire278(wire269));
  always
    @(posedge clk) begin
      reg345 = $signed({$signed((7'h44)), $unsigned(wire272)});
    end
  always
    @(posedge clk) begin
      reg346 = (&$signed((((wire272 <<< (8'ha6)) ?
              (reg345 ~^ (8'hb8)) : (wire271 <= (8'hbc))) ?
          ((wire272 ?
              wire271 : wire269) && $unsigned((8'h9f))) : $signed((wire271 ?
              (8'hb3) : wire269)))));
    end
  assign wire347 = (~|wire343);
  assign wire348 = $unsigned(((($signed((7'h44)) ?
                       wire343[(1'h1):(1'h0)] : $signed((8'hba))) > (&$signed(reg345))) > (~wire268[(2'h2):(1'h1)])));
  assign wire349 = wire271[(3'h5):(1'h0)];
  always
    @(posedge clk) begin
      reg350 = $signed($unsigned(wire271));
      reg351 <= $signed(wire271[(1'h0):(1'h0)]);
      reg352 <= $unsigned($unsigned(reg351[(4'hb):(3'h5)]));
      reg353 <= reg346;
      reg354 <= ((~^reg353) ?
          wire347[(2'h3):(2'h2)] : (wire268[(1'h1):(1'h1)] ?
              (wire343[(1'h1):(1'h0)] ?
                  ($unsigned(wire268) < $signed(wire270)) : $signed((8'hb6))) : $signed(((^~wire271) << $signed(wire348)))));
    end
  always
    @(posedge clk) begin
      reg355 = reg354[(1'h0):(1'h0)];
      reg356 <= $unsigned((~$signed($signed(wire268[(3'h5):(2'h2)]))));
      reg357 <= wire268[(1'h1):(1'h1)];
    end
  assign wire358 = (^~reg351[(2'h3):(1'h0)]);
  always
    @(posedge clk) begin
      reg359 <= wire349[(1'h1):(1'h1)];
    end
  assign wire360 = $signed(($unsigned(reg352) >>> wire272[(2'h2):(1'h1)]));
  assign wire361 = $signed(reg345[(3'h6):(2'h3)]);
  always
    @(posedge clk) begin
      reg362 <= $unsigned($unsigned($unsigned((reg350[(3'h4):(2'h3)] && $signed(reg345)))));
    end
  module363 modinst466 (wire465, clk, reg351, wire268, reg354, reg356);
  assign wire467 = (wire272 | ($signed($signed(reg362)) == wire348[(3'h6):(2'h3)]));
  assign wire468 = $unsigned((8'haa));
  always
    @(posedge clk) begin
      reg469 = wire358[(4'h8):(3'h4)];
      reg470 <= ($signed(((|wire348) != wire268[(1'h0):(1'h0)])) ^~ ((wire360 ?
              ((~&wire272) ?
                  (reg359 ?
                      (8'hb7) : wire349) : (+wire467)) : (wire348[(2'h3):(2'h3)] ?
                  wire361[(2'h2):(2'h2)] : (|wire273))) ?
          ($unsigned((|wire348)) >> $signed($signed(wire272))) : (^({reg355,
                  wire468} ?
              (reg355 >>> reg355) : (wire272 & wire347)))));
      for (forvar471 = (1'h0); (forvar471 < (1'h0)); forvar471 = (forvar471 + (1'h1)))
        begin
          reg472 <= (~&$signed(wire269));
          for (forvar473 = (1'h0); (forvar473 < (3'h4)); forvar473 = (forvar473 + (1'h1)))
            begin
              reg474 <= $signed(wire273);
              reg475 <= (!((wire343 >> $signed(reg474[(1'h1):(1'h1)])) ?
                  reg470 : {wire467, wire270[(5'h10):(2'h3)]}));
              reg476 <= reg472[(2'h2):(1'h1)];
              reg477 <= ((&$unsigned($unsigned(reg353[(2'h2):(2'h2)]))) <= ((wire349 != ($unsigned(reg353) << $unsigned((8'ha8)))) ^~ $signed($signed({wire468}))));
              reg478 <= $signed(wire465);
            end
          for (forvar479 = (1'h0); (forvar479 < (2'h2)); forvar479 = (forvar479 + (1'h1)))
            begin
              reg480 <= reg478;
              reg481 <= (^(reg356 ?
                  reg346 : ({wire360, $signed(reg345)} ?
                      wire347[(4'hb):(4'h9)] : $signed($unsigned(reg362)))));
              reg482 <= (~|($signed((8'ha9)) ?
                  $signed($unsigned($unsigned(wire358))) : {$signed($unsigned(wire269))}));
              reg483 <= (forvar473[(4'he):(3'h6)] ?
                  (~|$unsigned($unsigned((reg355 ?
                      reg475 : wire271)))) : $unsigned({(~&wire358[(1'h1):(1'h1)])}));
            end
          for (forvar484 = (1'h0); (forvar484 < (2'h3)); forvar484 = (forvar484 + (1'h1)))
            begin
              reg485 <= ($signed((^~forvar471)) <<< ({reg356, wire347} ?
                  reg353 : $signed({reg474[(2'h3):(1'h1)],
                      $signed(forvar473)})));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module210
#( parameter param255 = (({{(!(8'hbd)), ((8'hac) ? (8'haf) : (8'hbc))}, (!(8'ha6))} ? ((((7'h42) >= (8'haf)) ? ((8'hb2) * (8'ha1)) : ((8'hb5) ? (8'hb8) : (8'hba))) ? ((+(8'hb7)) && ((8'ha4) ? (8'hbf) : (8'haa))) : (((8'ha3) ? (7'h40) : (7'h40)) <<< ((8'hb9) < (8'hb6)))) : (~|((+(8'hb7)) ? ((8'hab) + (8'ha9)) : ((8'ha4) * (8'hb1))))) ? (-(8'hbf)) : ((-({(8'had), (8'h9e)} >> (-(8'hbe)))) ~^ (~&((+(8'h9f)) << {(8'hbd), (8'hbd)}))))
, parameter param256 = (({({param255} ? (param255 ? param255 : param255) : (param255 != (8'hab)))} ? ({param255} ^~ (param255 * (param255 ? param255 : param255))) : {param255, (^(param255 ? param255 : param255))}) && {((~^(8'hae)) ? {(~^param255), (param255 ? param255 : param255)} : {param255})}) )
(y, clk, wire215, wire214, wire213, wire212, wire211);
  output wire [(32'h1c3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire215;
  input wire [(4'hb):(1'h0)] wire214;
  input wire [(5'h13):(1'h0)] wire213;
  input wire signed [(3'h6):(1'h0)] wire212;
  input wire signed [(5'h10):(1'h0)] wire211;
  reg signed [(4'hf):(1'h0)] reg254 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg253 = (1'h0);
  reg [(5'h12):(1'h0)] reg252 = (1'h0);
  reg [(5'h13):(1'h0)] reg251 = (1'h0);
  reg [(4'h8):(1'h0)] reg250 = (1'h0);
  reg [(3'h6):(1'h0)] reg249 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar248 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire247;
  wire signed [(3'h5):(1'h0)] wire246;
  reg signed [(4'ha):(1'h0)] reg245 = (1'h0);
  reg [(3'h7):(1'h0)] reg244 = (1'h0);
  reg [(5'h13):(1'h0)] reg243 = (1'h0);
  reg [(3'h7):(1'h0)] reg242 = (1'h0);
  reg [(4'hd):(1'h0)] reg241 = (1'h0);
  reg [(5'h15):(1'h0)] forvar240 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg239 = (1'h0);
  reg [(4'hd):(1'h0)] reg238 = (1'h0);
  wire [(4'ha):(1'h0)] wire237;
  reg signed [(3'h5):(1'h0)] reg236 = (1'h0);
  reg [(4'hb):(1'h0)] reg235 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar234 = (1'h0);
  reg [(3'h4):(1'h0)] reg233 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg232 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire231;
  wire [(4'ha):(1'h0)] wire230;
  wire [(3'h7):(1'h0)] wire229;
  wire [(4'ha):(1'h0)] wire228;
  reg signed [(5'h12):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg226 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg225 = (1'h0);
  reg [(4'ha):(1'h0)] forvar224 = (1'h0);
  reg [(4'h8):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg222 = (1'h0);
  reg [(5'h12):(1'h0)] reg221 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg219 = (1'h0);
  reg [(4'he):(1'h0)] reg218 = (1'h0);
  reg signed [(4'he):(1'h0)] reg217 = (1'h0);
  wire [(5'h12):(1'h0)] wire216;
  assign y = {reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 forvar248,
                 wire247,
                 wire246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 forvar240,
                 reg239,
                 reg238,
                 wire237,
                 reg236,
                 reg235,
                 forvar234,
                 reg233,
                 reg232,
                 wire231,
                 wire230,
                 wire229,
                 wire228,
                 reg227,
                 reg226,
                 reg225,
                 forvar224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 wire216,
                 (1'h0)};
  assign wire216 = (+wire215);
  always
    @(posedge clk) begin
      reg217 <= (wire211 ?
          ((7'h40) ?
              wire212 : ($unsigned(wire214[(1'h1):(1'h0)]) ?
                  $signed((wire214 < wire213)) : $signed((wire212 <= (7'h40))))) : $unsigned(($signed($unsigned(wire211)) || (wire212 > $signed(wire215)))));
      reg218 <= wire214;
      reg219 <= (~&wire216[(4'ha):(3'h5)]);
      reg220 = (|$unsigned((wire211[(3'h4):(1'h1)] << (~wire212[(3'h4):(1'h0)]))));
      reg221 <= (~$signed((7'h40)));
    end
  always
    @(posedge clk) begin
      reg222 <= (wire215[(3'h4):(2'h2)] ?
          $unsigned((({wire211, wire215} >> (8'hbb)) ?
              $signed((&wire213)) : $signed(((8'ha0) & reg220)))) : (wire213[(3'h5):(1'h0)] > (^$unsigned($signed(reg221)))));
      reg223 = reg221[(4'hb):(1'h0)];
      for (forvar224 = (1'h0); (forvar224 < (1'h1)); forvar224 = (forvar224 + (1'h1)))
        begin
          reg225 <= {(~&(^~(reg217 ^~ (+reg219))))};
          reg226 <= reg218[(4'hb):(3'h7)];
          reg227 <= ((~(~|(8'hb4))) & reg219);
        end
    end
  assign wire228 = (7'h40);
  assign wire229 = ($signed(reg222[(3'h4):(1'h0)]) > $signed(reg222[(4'hc):(1'h1)]));
  assign wire230 = reg222;
  assign wire231 = wire214[(4'hb):(3'h7)];
  always
    @(posedge clk) begin
      reg232 <= $signed({$signed(wire230[(2'h2):(1'h1)]), wire229});
      reg233 <= (|$unsigned((+$signed((reg225 & wire211)))));
      for (forvar234 = (1'h0); (forvar234 < (3'h4)); forvar234 = (forvar234 + (1'h1)))
        begin
          reg235 <= $unsigned({$signed((^~$signed(reg219))),
              (wire231[(2'h2):(2'h2)] == $signed($signed(reg219)))});
          reg236 <= (^~(8'h9f));
        end
    end
  assign wire237 = reg219;
  always
    @(posedge clk) begin
      reg238 <= $unsigned($unsigned(($signed((~wire228)) == ((reg235 * wire213) ?
          (reg235 ~^ (8'hbc)) : (|reg225)))));
      reg239 <= {$unsigned($signed(reg221))};
      for (forvar240 = (1'h0); (forvar240 < (2'h3)); forvar240 = (forvar240 + (1'h1)))
        begin
          reg241 <= (($signed((reg217[(3'h6):(2'h3)] ~^ (forvar224 ?
                  reg221 : reg225))) ?
              (~&$signed((~&reg218))) : ({(&reg223)} ?
                  ($signed(wire213) ?
                      $signed((8'hb4)) : reg238[(1'h0):(1'h0)]) : (^(~|reg227)))) - wire215[(1'h1):(1'h0)]);
          reg242 <= wire215[(3'h7):(1'h0)];
          reg243 = (($signed(reg241[(3'h6):(3'h5)]) ?
                  {($signed(reg226) && reg222[(4'h9):(3'h4)]),
                      $unsigned((wire213 | wire230))} : wire229) ?
              {wire237} : wire211);
        end
      reg244 <= $unsigned(wire231[(1'h0):(1'h0)]);
      reg245 <= (-$signed(wire213[(4'he):(1'h0)]));
    end
  assign wire246 = ({(reg217 | ({reg222, reg226} ?
                               (forvar234 & reg239) : $unsigned(reg232)))} ?
                       reg244 : $unsigned(wire229[(2'h2):(1'h1)]));
  assign wire247 = $unsigned({(8'hae)});
  always
    @(posedge clk) begin
      for (forvar248 = (1'h0); (forvar248 < (2'h3)); forvar248 = (forvar248 + (1'h1)))
        begin
          reg249 <= wire211[(3'h7):(2'h2)];
          if ((~($unsigned(reg241) ?
              reg241[(4'h9):(3'h7)] : (((~|wire237) <= (reg220 ?
                  wire247 : reg227)) <= forvar240))))
            begin
              reg250 <= ({{$signed($signed(reg225))},
                  wire246} & $signed((forvar248 ?
                  reg241[(4'hb):(3'h7)] : ((wire246 || reg232) ?
                      $signed(reg225) : (|reg239)))));
            end
          else
            begin
              reg250 <= reg221;
              reg251 <= $unsigned($signed((reg223[(3'h7):(3'h7)] ?
                  $unsigned($unsigned(reg218)) : $signed((-(8'hab))))));
            end
          reg252 <= (7'h43);
        end
      reg253 <= {(($signed((-reg232)) > {reg219}) ?
              $unsigned($unsigned((!reg233))) : $unsigned((~|((8'ha9) ^~ (8'h9c))))),
          (~$signed(reg244[(3'h5):(3'h5)]))};
      reg254 <= wire231;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module142  (y, clk, wire147, wire146, wire145, wire144, wire143);
  output wire [(32'h36):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire147;
  input wire [(4'ha):(1'h0)] wire146;
  input wire signed [(5'h10):(1'h0)] wire145;
  input wire signed [(5'h13):(1'h0)] wire144;
  input wire signed [(3'h6):(1'h0)] wire143;
  wire [(3'h4):(1'h0)] wire182;
  wire [(4'hf):(1'h0)] wire180;
  wire signed [(5'h11):(1'h0)] wire150;
  reg signed [(4'he):(1'h0)] reg149 = (1'h0);
  reg [(2'h3):(1'h0)] reg148 = (1'h0);
  assign y = {wire182, wire180, wire150, reg149, reg148, (1'h0)};
  always
    @(posedge clk) begin
      reg148 <= {$signed({(8'hbe), $unsigned({wire146, (8'hbd)})}),
          ($unsigned(wire147[(3'h7):(1'h0)]) ?
              (8'ha2) : $signed({(wire144 ? wire147 : wire143)}))};
    end
  always
    @(posedge clk) begin
      reg149 <= $signed((+$signed(wire143)));
    end
  assign wire150 = wire145[(4'hb):(1'h0)];
  module151 modinst181 (wire180, clk, wire147, wire145, reg149, wire150);
  assign wire182 = {wire150[(5'h11):(4'he)],
                       ($unsigned((7'h40)) ?
                           $signed(wire143[(2'h3):(1'h1)]) : (~((!reg148) != $unsigned(wire147))))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module151
#( parameter param178 = ((((((8'ha8) ? (8'ha1) : (8'hb1)) ? ((8'haa) >> (8'h9d)) : (^(7'h42))) << ((^~(8'ha9)) ? ((8'hb8) ? (8'ha6) : (8'ha0)) : ((7'h43) ? (8'hbb) : (8'hb5)))) ? (~^(~&{(7'h41)})) : ({((8'h9e) ? (7'h40) : (8'hae)), ((8'hb1) | (8'h9d))} != (((8'hac) - (8'hb1)) ? (8'hb1) : {(8'ha6), (7'h40)}))) ? (^((((8'hab) ^~ (8'hb4)) ? ((8'hb9) ? (8'h9d) : (8'ha6)) : (-(8'ha1))) > (((8'hb4) & (8'ha6)) ? ((8'hbf) >> (8'ha0)) : ((8'ha5) ? (8'haa) : (8'hb8))))) : ((((&(8'hae)) ^ ((8'hb0) & (8'hb9))) * (((8'hb6) * (8'hb1)) ^ ((8'ha1) ? (8'h9c) : (8'hb8)))) ? ((((7'h43) ? (8'hb2) : (8'hba)) > ((8'ha6) < (8'h9f))) ^~ {{(8'ha9)}, ((8'hab) ? (8'ha7) : (8'ha1))}) : (((&(8'ha4)) ? (+(8'hbc)) : (!(7'h42))) ? (~^{(8'haf)}) : (((8'hb4) ? (7'h41) : (8'hb8)) ? ((8'hb9) << (8'ha0)) : ((8'hb7) * (8'hb8))))))
, parameter param179 = (param178 ? ({{(^~param178)}} ^ param178) : (!((!param178) ? ({param178} | param178) : (+{param178})))) )
(y, clk, wire155, wire154, wire153, wire152);
  output wire [(32'hea):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire155;
  input wire signed [(5'h10):(1'h0)] wire154;
  input wire [(3'h6):(1'h0)] wire153;
  input wire [(5'h11):(1'h0)] wire152;
  reg signed [(4'hc):(1'h0)] reg177 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg176 = (1'h0);
  reg [(2'h2):(1'h0)] reg175 = (1'h0);
  reg [(3'h4):(1'h0)] forvar174 = (1'h0);
  reg [(5'h13):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar172 = (1'h0);
  reg [(4'hd):(1'h0)] reg171 = (1'h0);
  reg [(5'h10):(1'h0)] forvar170 = (1'h0);
  wire [(2'h3):(1'h0)] wire169;
  wire signed [(4'hc):(1'h0)] wire168;
  wire [(3'h6):(1'h0)] wire167;
  wire [(4'h9):(1'h0)] wire166;
  reg [(4'he):(1'h0)] reg165 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire164;
  wire [(4'hf):(1'h0)] wire163;
  reg [(4'hb):(1'h0)] reg162 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg161 = (1'h0);
  reg [(5'h13):(1'h0)] reg160 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire159;
  reg [(3'h6):(1'h0)] reg158 = (1'h0);
  wire [(4'hf):(1'h0)] wire157;
  wire signed [(2'h3):(1'h0)] wire156;
  assign y = {reg177,
                 reg176,
                 reg175,
                 forvar174,
                 reg173,
                 forvar172,
                 reg171,
                 forvar170,
                 wire169,
                 wire168,
                 wire167,
                 wire166,
                 reg165,
                 wire164,
                 wire163,
                 reg162,
                 reg161,
                 reg160,
                 wire159,
                 reg158,
                 wire157,
                 wire156,
                 (1'h0)};
  assign wire156 = (($signed({wire155[(2'h3):(1'h0)],
                           ((8'ha5) ?
                               wire155 : wire154)}) & wire152[(4'hd):(4'h9)]) ?
                       $unsigned((wire152[(2'h2):(1'h1)] + ($signed(wire152) == {wire153,
                           wire153}))) : wire153);
  assign wire157 = wire153;
  always
    @(posedge clk) begin
      reg158 <= wire156[(2'h2):(1'h1)];
    end
  assign wire159 = ((($signed($signed((8'hbb))) ?
                           $unsigned(wire152[(4'hc):(3'h5)]) : ((wire157 ?
                                   wire153 : wire152) ?
                               (wire153 <<< wire152) : (reg158 ~^ (8'ha1)))) ~^ wire156[(2'h2):(1'h0)]) ?
                       $unsigned($signed($unsigned($signed(wire157)))) : ((-$signed($unsigned((8'hb9)))) & ($signed((!wire154)) ?
                           {{reg158, wire155},
                               (wire157 ^~ wire156)} : ((^wire153) ?
                               wire152 : $unsigned(wire152)))));
  always
    @(posedge clk) begin
      if ({$signed((wire154[(4'ha):(4'h8)] ?
              $unsigned(wire159[(4'hf):(4'he)]) : ($signed(wire156) ?
                  $unsigned(reg158) : (~^wire152))))})
        begin
          reg160 = wire159[(4'hc):(4'ha)];
          reg161 <= $signed(((8'h9f) ? (~&wire152[(4'hd):(1'h0)]) : (8'hbe)));
          reg162 <= wire159;
        end
      else
        begin
          reg160 <= wire157[(1'h0):(1'h0)];
        end
    end
  assign wire163 = {$signed((-(wire152[(1'h0):(1'h0)] < $signed(reg162))))};
  assign wire164 = ({(~^wire155),
                       (^((&wire155) << $unsigned(reg158)))} && $signed(((^(^wire159)) & reg161)));
  always
    @(posedge clk) begin
      reg165 = $signed($unsigned(($signed($unsigned(wire156)) | wire153[(1'h0):(1'h0)])));
    end
  assign wire166 = wire163;
  assign wire167 = ((wire152 + (^~$unsigned((!(8'hb3))))) ?
                       {$unsigned((wire164 && (wire159 ^ wire157))),
                           wire166[(4'h9):(2'h2)]} : reg160);
  assign wire168 = $unsigned($unsigned($signed(reg160[(4'hf):(3'h4)])));
  assign wire169 = $unsigned((8'ha0));
  always
    @(posedge clk) begin
      for (forvar170 = (1'h0); (forvar170 < (2'h3)); forvar170 = (forvar170 + (1'h1)))
        begin
          reg171 <= reg165[(4'ha):(4'ha)];
        end
      for (forvar172 = (1'h0); (forvar172 < (1'h1)); forvar172 = (forvar172 + (1'h1)))
        begin
          reg173 = reg165[(3'h4):(1'h0)];
        end
      for (forvar174 = (1'h0); (forvar174 < (3'h4)); forvar174 = (forvar174 + (1'h1)))
        begin
          reg175 <= (8'hbf);
          reg176 <= ({($unsigned(wire167[(3'h5):(2'h3)]) ?
                      $signed(reg175[(1'h0):(1'h0)]) : {{reg173}}),
                  (~(wire159[(3'h4):(1'h0)] ?
                      wire156 : wire154[(1'h1):(1'h1)]))} ?
              (reg175[(2'h2):(1'h0)] ?
                  {(((8'ha7) * wire156) ?
                          $unsigned((8'hbe)) : $unsigned((7'h40))),
                      (^~{wire153})} : $unsigned($signed(wire164))) : $unsigned($unsigned(forvar172[(1'h0):(1'h0)])));
          reg177 <= {wire164[(4'hd):(4'ha)]};
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module363
#( parameter param464 = ((((((8'haf) ? (7'h44) : (8'ha8)) - (-(7'h44))) ? {((8'ha9) & (8'h9d))} : (((8'ha6) ? (8'ha4) : (7'h42)) | (8'hb3))) ? (~&(((8'hb1) ? (8'hba) : (7'h44)) >> ((8'ha5) ? (8'h9d) : (8'hbd)))) : (({(8'ha6)} || ((8'haa) ^~ (8'haf))) < (^~{(8'hbe)}))) || (&{(~^((8'hb6) ? (8'ha9) : (7'h44)))})) )
(y, clk, wire367, wire366, wire365, wire364);
  output wire [(32'h464):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire367;
  input wire signed [(4'hb):(1'h0)] wire366;
  input wire signed [(4'hd):(1'h0)] wire365;
  input wire signed [(3'h6):(1'h0)] wire364;
  reg signed [(5'h14):(1'h0)] reg463 = (1'h0);
  reg [(5'h10):(1'h0)] reg462 = (1'h0);
  reg [(5'h15):(1'h0)] reg461 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg460 = (1'h0);
  reg [(3'h7):(1'h0)] reg459 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar458 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar457 = (1'h0);
  reg [(4'ha):(1'h0)] reg456 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire455;
  reg [(4'hb):(1'h0)] reg454 = (1'h0);
  reg [(2'h3):(1'h0)] reg453 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg452 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg451 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg450 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg449 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar448 = (1'h0);
  reg [(4'he):(1'h0)] reg447 = (1'h0);
  reg [(4'h8):(1'h0)] reg446 = (1'h0);
  reg [(3'h4):(1'h0)] forvar445 = (1'h0);
  reg [(4'h8):(1'h0)] reg444 = (1'h0);
  reg [(5'h11):(1'h0)] reg443 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar442 = (1'h0);
  reg [(4'hc):(1'h0)] forvar441 = (1'h0);
  reg [(4'hf):(1'h0)] reg440 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire439;
  reg [(4'hb):(1'h0)] reg438 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg437 = (1'h0);
  reg [(2'h3):(1'h0)] reg436 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg435 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg434 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg433 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg432 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar431 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg430 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg429 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg428 = (1'h0);
  reg [(3'h7):(1'h0)] forvar427 = (1'h0);
  reg [(4'h8):(1'h0)] forvar426 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg425 = (1'h0);
  reg [(3'h5):(1'h0)] reg424 = (1'h0);
  reg [(5'h10):(1'h0)] reg423 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg422 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg421 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg420 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar419 = (1'h0);
  reg [(4'h8):(1'h0)] forvar418 = (1'h0);
  wire [(5'h12):(1'h0)] wire417;
  reg signed [(2'h3):(1'h0)] reg416 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg415 = (1'h0);
  reg [(5'h10):(1'h0)] reg414 = (1'h0);
  reg [(2'h3):(1'h0)] reg413 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire412;
  reg [(4'hd):(1'h0)] reg411 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar410 = (1'h0);
  reg [(4'hf):(1'h0)] reg409 = (1'h0);
  reg [(4'hf):(1'h0)] reg408 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar407 = (1'h0);
  reg [(3'h7):(1'h0)] reg406 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg405 = (1'h0);
  reg [(5'h11):(1'h0)] reg404 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg403 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg402 = (1'h0);
  reg [(4'hd):(1'h0)] reg401 = (1'h0);
  reg [(4'he):(1'h0)] reg400 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg399 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar398 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg397 = (1'h0);
  reg [(4'ha):(1'h0)] reg396 = (1'h0);
  reg [(4'hd):(1'h0)] reg395 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg394 = (1'h0);
  reg [(3'h4):(1'h0)] reg393 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg392 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg391 = (1'h0);
  reg signed [(4'he):(1'h0)] reg390 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar389 = (1'h0);
  reg [(4'h9):(1'h0)] forvar388 = (1'h0);
  reg [(5'h10):(1'h0)] reg387 = (1'h0);
  reg [(4'hd):(1'h0)] reg386 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg385 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg384 = (1'h0);
  reg [(5'h14):(1'h0)] reg383 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar382 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg380 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg379 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg378 = (1'h0);
  reg [(4'ha):(1'h0)] forvar377 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg376 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg375 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire374;
  wire signed [(5'h14):(1'h0)] wire373;
  wire signed [(4'hd):(1'h0)] wire372;
  wire [(3'h5):(1'h0)] wire371;
  reg [(5'h15):(1'h0)] reg370 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg369 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire368;
  assign y = {reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 forvar458,
                 forvar457,
                 reg456,
                 wire455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 forvar448,
                 reg447,
                 reg446,
                 forvar445,
                 reg444,
                 reg443,
                 forvar442,
                 forvar441,
                 reg440,
                 wire439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 forvar431,
                 reg430,
                 reg429,
                 reg428,
                 forvar427,
                 forvar426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 forvar419,
                 forvar418,
                 wire417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 wire412,
                 reg411,
                 forvar410,
                 reg409,
                 reg408,
                 forvar407,
                 reg406,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 forvar398,
                 reg397,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 forvar389,
                 forvar388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 forvar382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 forvar377,
                 reg376,
                 reg375,
                 wire374,
                 wire373,
                 wire372,
                 wire371,
                 reg370,
                 reg369,
                 wire368,
                 (1'h0)};
  assign wire368 = (|(((wire365[(3'h5):(1'h0)] ?
                               (&wire367) : (wire364 ? wire364 : wire366)) ?
                           $unsigned((~wire364)) : $signed((wire366 ?
                               wire365 : wire367))) ?
                       wire365 : ($signed($unsigned(wire364)) + $signed($signed(wire364)))));
  always
    @(posedge clk) begin
      reg369 = wire366;
      reg370 = {wire366};
    end
  assign wire371 = $signed((~^$unsigned($unsigned($signed(wire367)))));
  assign wire372 = wire365[(3'h7):(3'h4)];
  assign wire373 = (wire366[(3'h4):(1'h0)] ?
                       (wire365 ?
                           (^~$unsigned(wire372[(4'hb):(4'ha)])) : (({reg369,
                                   reg370} - {wire367, wire368}) ?
                               (reg369[(3'h6):(1'h0)] ?
                                   $signed(reg370) : {wire371}) : {(wire371 == wire371)})) : $signed(((8'hb2) ?
                           (^(~^wire364)) : ($unsigned(wire372) ?
                               $signed(wire372) : $signed(reg369)))));
  assign wire374 = ($unsigned((reg369 >>> {(reg370 ?
                           (8'hab) : wire367)})) <= $signed($signed(((~wire371) ?
                       (wire364 ? (8'hb4) : wire367) : (-(8'hb1))))));
  always
    @(posedge clk) begin
      reg375 <= (reg369 ?
          $unsigned((8'hb0)) : $unsigned(wire374[(2'h2):(2'h2)]));
      reg376 = (8'hb9);
      for (forvar377 = (1'h0); (forvar377 < (2'h2)); forvar377 = (forvar377 + (1'h1)))
        begin
          reg378 = $signed(wire367[(1'h1):(1'h1)]);
          reg379 <= (forvar377[(3'h5):(2'h3)] ^ reg369);
          reg380 = (((reg375[(4'h9):(2'h3)] ?
                      wire374 : reg379[(5'h12):(4'hd)]) ?
                  {$unsigned(wire368[(4'ha):(1'h1)]),
                      (wire374[(1'h1):(1'h1)] ?
                          (-reg369) : (forvar377 ?
                              (8'ha5) : forvar377))} : $signed((wire364 > (forvar377 ?
                      wire366 : wire373)))) ?
              (wire364 ?
                  wire366[(1'h1):(1'h0)] : wire373) : ($signed((((7'h42) ?
                          reg369 : reg369) ?
                      (+wire374) : (wire371 ? reg376 : reg376))) ?
                  wire373[(5'h11):(4'h9)] : reg369));
          reg381 = $signed(($signed($unsigned(wire372[(1'h1):(1'h1)])) ~^ $signed(({forvar377,
                  wire366} ?
              wire372[(4'hb):(3'h7)] : $unsigned(reg370)))));
          for (forvar382 = (1'h0); (forvar382 < (1'h0)); forvar382 = (forvar382 + (1'h1)))
            begin
              reg383 = reg376;
              reg384 <= $signed(reg370);
              reg385 = $unsigned((reg375 ?
                  ($signed({wire364}) ^~ ((reg380 ? (8'hbd) : wire372) ?
                      ((8'h9e) <<< reg369) : (8'hbf))) : wire365[(4'hd):(4'hc)]));
              reg386 = reg381;
              reg387 <= ($signed($unsigned($signed({reg369}))) ?
                  wire367 : (|reg380[(3'h5):(1'h0)]));
            end
        end
      for (forvar388 = (1'h0); (forvar388 < (2'h2)); forvar388 = (forvar388 + (1'h1)))
        begin
          for (forvar389 = (1'h0); (forvar389 < (2'h2)); forvar389 = (forvar389 + (1'h1)))
            begin
              reg390 <= (+$unsigned(reg380[(2'h2):(2'h2)]));
              reg391 = wire373;
              reg392 <= wire368;
              reg393 <= reg379[(4'hb):(4'hb)];
              reg394 = $signed(reg375);
            end
        end
      reg395 <= reg385;
    end
  always
    @(posedge clk) begin
      reg396 <= ($unsigned($signed(reg392[(1'h0):(1'h0)])) ?
          {{(-(reg385 >>> wire373))}} : reg381[(3'h5):(2'h3)]);
    end
  always
    @(posedge clk) begin
      reg397 = $unsigned(($unsigned($signed((~|wire366))) ~^ (+{reg385,
          (|reg380)})));
      for (forvar398 = (1'h0); (forvar398 < (2'h3)); forvar398 = (forvar398 + (1'h1)))
        begin
          reg399 <= (&(($unsigned($unsigned(reg392)) <<< $unsigned(reg376)) ?
              reg394 : reg395[(3'h4):(2'h2)]));
          reg400 <= ($signed($signed(((forvar389 >>> reg378) ?
                  reg370 : $unsigned(reg394)))) ?
              reg390 : reg395);
          reg401 <= reg390;
          reg402 = (($unsigned(((~(8'hb2)) ?
                      forvar377[(4'ha):(1'h1)] : reg381)) ?
                  $unsigned(reg393) : forvar382[(4'h8):(1'h1)]) ?
              (forvar388 < forvar398) : $signed($signed($unsigned((reg394 ?
                  wire367 : forvar382)))));
          reg403 = ($signed(((~&(reg380 ? reg396 : reg402)) << {(reg397 ?
                  reg391 : reg386),
              $unsigned(wire368)})) <= (^~(reg391[(3'h5):(1'h0)] ^ (reg378 ?
              (|reg397) : (reg401 == wire371)))));
        end
      reg404 <= ($signed(reg386) ?
          $signed($unsigned((^$signed(reg395)))) : $unsigned(forvar388[(2'h2):(1'h1)]));
      reg405 <= (reg376 <<< $signed(((wire366 + (8'hb3)) != ($unsigned(reg400) != forvar388))));
      reg406 = {reg380, reg378};
    end
  always
    @(posedge clk) begin
      for (forvar407 = (1'h0); (forvar407 < (3'h4)); forvar407 = (forvar407 + (1'h1)))
        begin
          reg408 <= reg381[(4'h9):(3'h5)];
          reg409 <= $unsigned(reg392);
        end
      for (forvar410 = (1'h0); (forvar410 < (3'h4)); forvar410 = (forvar410 + (1'h1)))
        begin
          reg411 <= {reg406,
              (|(wire365 ^ ((forvar377 < forvar398) ?
                  $signed(reg405) : wire367)))};
        end
    end
  assign wire412 = wire373[(5'h12):(5'h10)];
  always
    @(posedge clk) begin
      reg413 <= $unsigned((((forvar410[(4'hd):(4'hc)] & (wire365 <= (8'haf))) ~^ ({wire368} ?
              $signed((8'had)) : reg379)) ?
          forvar388 : (8'ha5)));
      reg414 <= (reg397 ?
          wire371 : $unsigned(((reg383[(2'h2):(2'h2)] & reg378[(4'h9):(2'h2)]) ~^ reg391)));
      reg415 <= $signed($unsigned(reg381[(3'h5):(1'h1)]));
      reg416 <= (^~wire365[(1'h0):(1'h0)]);
    end
  assign wire417 = ($unsigned(reg383) ?
                       (&(~|$signed((7'h40)))) : (~^reg409[(2'h2):(1'h1)]));
  always
    @(posedge clk) begin
      for (forvar418 = (1'h0); (forvar418 < (2'h2)); forvar418 = (forvar418 + (1'h1)))
        begin
          for (forvar419 = (1'h0); (forvar419 < (1'h1)); forvar419 = (forvar419 + (1'h1)))
            begin
              reg420 <= reg379;
              reg421 = $signed((~^($signed(reg408[(3'h6):(3'h5)]) ?
                  $unsigned(forvar407) : $unsigned($unsigned(reg369)))));
              reg422 <= {($unsigned(((reg392 ? reg369 : (8'hb1)) ?
                          $unsigned(reg381) : (~forvar377))) ?
                      $unsigned((&$unsigned(reg397))) : (^~({wire417} <= (+reg403)))),
                  reg400[(3'h7):(3'h7)]};
              reg423 <= forvar388;
            end
          reg424 <= wire373;
        end
      reg425 = (|reg383);
      for (forvar426 = (1'h0); (forvar426 < (1'h0)); forvar426 = (forvar426 + (1'h1)))
        begin
          for (forvar427 = (1'h0); (forvar427 < (1'h1)); forvar427 = (forvar427 + (1'h1)))
            begin
              reg428 <= {reg392[(1'h1):(1'h1)],
                  $unsigned($signed(($unsigned((8'ha6)) + ((8'hba) + reg415))))};
              reg429 <= $unsigned($signed($unsigned(forvar419[(4'hd):(2'h2)])));
              reg430 <= (($unsigned({$unsigned(reg391), reg406}) ?
                      {(reg385 ? reg381[(1'h1):(1'h1)] : reg413[(2'h3):(1'h0)]),
                          ($unsigned(reg385) ?
                              $signed(reg400) : reg411)} : $unsigned((reg381 ?
                          $unsigned(wire368) : (-reg401)))) ?
                  (+reg422) : (~|reg403[(1'h0):(1'h0)]));
            end
          for (forvar431 = (1'h0); (forvar431 < (2'h3)); forvar431 = (forvar431 + (1'h1)))
            begin
              reg432 <= (reg391 ^ $unsigned(reg387[(3'h4):(3'h4)]));
            end
          reg433 = (wire368[(1'h0):(1'h0)] ?
              $unsigned({((8'hbd) * {reg399}), (&(8'ha7))}) : reg395);
        end
      reg434 = {reg395};
    end
  always
    @(posedge clk) begin
      reg435 <= ((~^forvar389[(1'h1):(1'h0)]) == $unsigned({($signed(reg370) < $unsigned(forvar388))}));
      reg436 <= forvar419[(4'hf):(3'h7)];
      reg437 <= {reg415};
      reg438 <= reg384[(4'h8):(4'h8)];
    end
  assign wire439 = {((!wire365) ?
                           $unsigned(($signed(reg414) ?
                               reg411[(1'h1):(1'h1)] : (~^wire371))) : ((8'ha3) ?
                               ($unsigned(reg420) ?
                                   $unsigned(reg402) : (forvar418 ?
                                       wire374 : wire372)) : wire374[(2'h3):(1'h1)]))};
  always
    @(posedge clk) begin
      reg440 = $signed({$signed((~(reg379 ^ reg387)))});
    end
  always
    @(posedge clk) begin
      for (forvar441 = (1'h0); (forvar441 < (2'h3)); forvar441 = (forvar441 + (1'h1)))
        begin
          for (forvar442 = (1'h0); (forvar442 < (1'h1)); forvar442 = (forvar442 + (1'h1)))
            begin
              reg443 <= (wire368[(2'h2):(1'h0)] * $signed((reg400 ?
                  forvar389 : $signed(forvar389))));
            end
          reg444 = $unsigned(reg405);
        end
      for (forvar445 = (1'h0); (forvar445 < (2'h2)); forvar445 = (forvar445 + (1'h1)))
        begin
          reg446 <= (~wire412[(4'ha):(1'h1)]);
        end
      reg447 = reg397;
      for (forvar448 = (1'h0); (forvar448 < (2'h3)); forvar448 = (forvar448 + (1'h1)))
        begin
          reg449 <= {((+reg394) << $signed((~&(~^reg396)))),
              $unsigned($signed($unsigned(reg433[(5'h12):(2'h3)])))};
          reg450 <= wire372;
          reg451 <= (wire417 + forvar419[(2'h3):(2'h2)]);
        end
      reg452 <= (~((((reg447 & reg384) ? reg396 : {wire372}) ?
              ((wire412 ?
                  forvar407 : (8'ha8)) & reg446[(3'h4):(2'h2)]) : $signed(reg391[(3'h6):(3'h4)])) ?
          (^(+$signed(reg450))) : (-wire368[(3'h7):(3'h4)])));
    end
  always
    @(posedge clk) begin
      reg453 <= forvar398[(3'h7):(2'h2)];
      reg454 = $signed($signed((+$unsigned(((8'hb2) && reg369)))));
    end
  assign wire455 = reg406;
  always
    @(posedge clk) begin
      reg456 <= ((8'hbb) ? forvar388 : $unsigned((~reg421)));
      for (forvar457 = (1'h0); (forvar457 < (2'h2)); forvar457 = (forvar457 + (1'h1)))
        begin
          for (forvar458 = (1'h0); (forvar458 < (1'h1)); forvar458 = (forvar458 + (1'h1)))
            begin
              reg459 <= reg423;
              reg460 = reg394[(4'h8):(3'h4)];
              reg461 = ((reg381[(3'h6):(3'h6)] ?
                      {(!(-reg370))} : ($unsigned($signed(reg452)) ~^ (~wire364[(2'h2):(2'h2)]))) ?
                  (~{((~^reg375) ? $unsigned(forvar418) : $signed(reg430)),
                      ((reg380 ? reg381 : wire365) ?
                          reg401 : $signed(reg429))}) : (|(~^{(!wire365),
                      reg446[(2'h3):(1'h0)]})));
              reg462 <= reg428[(3'h7):(2'h3)];
            end
          reg463 = reg406[(3'h4):(3'h4)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module274  (y, clk, wire278, wire277, wire276, wire275);
  output wire [(32'h2f5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire278;
  input wire [(2'h3):(1'h0)] wire277;
  input wire [(3'h5):(1'h0)] wire276;
  input wire signed [(4'hf):(1'h0)] wire275;
  reg [(4'he):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg341 = (1'h0);
  reg [(4'h8):(1'h0)] reg340 = (1'h0);
  reg [(4'hb):(1'h0)] reg339 = (1'h0);
  reg [(5'h10):(1'h0)] reg338 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg337 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg336 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg335 = (1'h0);
  reg [(5'h10):(1'h0)] forvar334 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg333 = (1'h0);
  reg [(2'h3):(1'h0)] reg332 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg331 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg329 = (1'h0);
  reg [(4'h9):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar327 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar326 = (1'h0);
  reg [(5'h14):(1'h0)] reg325 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg324 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg322 = (1'h0);
  wire [(5'h11):(1'h0)] wire321;
  reg signed [(3'h6):(1'h0)] reg320 = (1'h0);
  reg [(5'h15):(1'h0)] reg319 = (1'h0);
  reg [(3'h5):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg317 = (1'h0);
  reg [(4'hb):(1'h0)] reg316 = (1'h0);
  reg [(4'he):(1'h0)] reg315 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire314;
  wire signed [(4'h9):(1'h0)] wire313;
  wire [(4'hb):(1'h0)] wire312;
  reg [(5'h11):(1'h0)] reg311 = (1'h0);
  reg [(5'h15):(1'h0)] reg310 = (1'h0);
  reg [(2'h2):(1'h0)] reg309 = (1'h0);
  reg [(5'h11):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg307 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg306 = (1'h0);
  reg [(4'hb):(1'h0)] reg305 = (1'h0);
  reg [(2'h2):(1'h0)] forvar304 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar303 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg302 = (1'h0);
  reg [(4'he):(1'h0)] reg301 = (1'h0);
  reg [(5'h12):(1'h0)] reg300 = (1'h0);
  wire [(2'h2):(1'h0)] wire299;
  reg [(5'h11):(1'h0)] reg298 = (1'h0);
  reg [(4'hb):(1'h0)] reg297 = (1'h0);
  reg [(4'h8):(1'h0)] forvar296 = (1'h0);
  reg [(5'h15):(1'h0)] reg295 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg294 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg293 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg291 = (1'h0);
  reg [(2'h2):(1'h0)] reg290 = (1'h0);
  reg [(2'h3):(1'h0)] reg289 = (1'h0);
  reg [(5'h12):(1'h0)] reg288 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg287 = (1'h0);
  reg [(5'h15):(1'h0)] reg286 = (1'h0);
  reg [(4'h8):(1'h0)] forvar285 = (1'h0);
  reg [(4'he):(1'h0)] reg284 = (1'h0);
  reg [(4'hb):(1'h0)] reg283 = (1'h0);
  reg [(5'h13):(1'h0)] forvar282 = (1'h0);
  reg [(2'h3):(1'h0)] forvar281 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg280 = (1'h0);
  reg [(4'h8):(1'h0)] reg279 = (1'h0);
  assign y = {reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 forvar334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 forvar327,
                 forvar326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 wire321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 wire314,
                 wire313,
                 wire312,
                 reg311,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 forvar304,
                 forvar303,
                 reg302,
                 reg301,
                 reg300,
                 wire299,
                 reg298,
                 reg297,
                 forvar296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 forvar285,
                 reg284,
                 reg283,
                 forvar282,
                 forvar281,
                 reg280,
                 reg279,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg279 = wire277;
      reg280 <= (8'hb0);
      for (forvar281 = (1'h0); (forvar281 < (3'h4)); forvar281 = (forvar281 + (1'h1)))
        begin
          for (forvar282 = (1'h0); (forvar282 < (2'h2)); forvar282 = (forvar282 + (1'h1)))
            begin
              reg283 <= ((~&wire275[(3'h6):(3'h4)]) ?
                  $unsigned($signed($unsigned(reg279))) : (($unsigned((wire278 ?
                      wire275 : wire277)) + wire278) >> forvar281));
              reg284 <= {($signed($signed((wire275 ?
                      forvar281 : wire277))) && reg280)};
            end
          for (forvar285 = (1'h0); (forvar285 < (2'h2)); forvar285 = (forvar285 + (1'h1)))
            begin
              reg286 = $unsigned(((($signed(wire276) ?
                  reg283 : $signed(forvar285)) >> ({(7'h42)} ?
                  ((8'h9d) < wire278) : (wire275 ?
                      forvar282 : reg283))) >>> (~&$signed(reg280))));
              reg287 <= reg286[(5'h12):(4'hd)];
              reg288 <= $signed((wire278[(5'h12):(3'h5)] | $signed((+$unsigned(wire278)))));
              reg289 <= wire276;
            end
          reg290 <= (reg287[(4'hd):(4'hb)] ?
              (~|reg286) : $unsigned((($signed((8'hac)) << reg289[(2'h3):(1'h0)]) & reg279)));
        end
      reg291 <= (($signed(((8'hac) ?
              $unsigned(reg283) : $signed(forvar282))) >>> reg279) ?
          ($signed($unsigned((reg283 - reg283))) ?
              $unsigned(reg289) : forvar282) : $unsigned({reg284[(3'h6):(3'h4)],
              forvar282}));
    end
  always
    @(posedge clk) begin
      reg292 <= $signed(({forvar285[(2'h3):(1'h0)],
          $signed((~forvar285))} && (8'ha5)));
      reg293 <= (~({$unsigned($unsigned((8'ha2))),
              $signed(reg291[(2'h2):(2'h2)])} ?
          {$unsigned((reg289 ? wire278 : reg286))} : reg288));
      reg294 = (({$signed($unsigned(reg292))} & reg289) - ({(~|$signed(reg290))} ?
          {(!(reg280 | (8'h9d)))} : $unsigned($signed((wire277 ?
              wire275 : reg291)))));
      reg295 <= ({$signed(((~(8'hb8)) & $unsigned((8'ha2))))} ?
          (~&forvar282[(4'hc):(1'h0)]) : ($unsigned($unsigned(forvar281)) << (+$signed($unsigned(wire275)))));
      for (forvar296 = (1'h0); (forvar296 < (3'h4)); forvar296 = (forvar296 + (1'h1)))
        begin
          reg297 = ($signed((^~$unsigned((reg291 ? wire275 : (8'hb7))))) ?
              ($unsigned({(-reg280)}) < (8'h9d)) : $unsigned(wire278[(4'ha):(1'h1)]));
          reg298 <= $signed($signed(forvar281[(2'h2):(1'h1)]));
        end
    end
  assign wire299 = (~^(+($unsigned((reg298 ? reg295 : reg287)) ?
                       {(|reg291)} : (reg290 ^~ $signed(reg280)))));
  always
    @(posedge clk) begin
      reg300 <= forvar285[(1'h1):(1'h1)];
      reg301 = $signed(reg300);
      reg302 <= reg301[(1'h0):(1'h0)];
      for (forvar303 = (1'h0); (forvar303 < (1'h0)); forvar303 = (forvar303 + (1'h1)))
        begin
          for (forvar304 = (1'h0); (forvar304 < (1'h1)); forvar304 = (forvar304 + (1'h1)))
            begin
              reg305 <= {$signed(reg280[(2'h2):(2'h2)])};
              reg306 <= $unsigned((&$unsigned(forvar304)));
              reg307 <= $signed(($unsigned(wire276[(3'h4):(1'h0)]) > $unsigned(reg301[(4'hb):(1'h1)])));
              reg308 <= $signed((reg306[(4'h9):(3'h4)] ?
                  {$unsigned((reg283 >= reg291)),
                      reg292[(2'h3):(2'h3)]} : (((7'h43) < (forvar281 ?
                      (8'hba) : reg300)) >>> $signed(reg284[(4'ha):(4'h8)]))));
              reg309 <= reg293[(3'h5):(2'h3)];
            end
          reg310 <= $unsigned(((((reg290 ? forvar281 : (8'ha5)) ?
                      reg309[(1'h0):(1'h0)] : $unsigned(forvar304)) ?
                  ($signed(reg292) ^ reg295) : $signed((reg284 ?
                      reg300 : reg280))) ?
              reg300[(4'hb):(4'h8)] : $unsigned(forvar296)));
          reg311 <= $unsigned(reg298);
        end
    end
  assign wire312 = {(!(^($signed(forvar282) <<< $signed(reg308)))), reg306};
  assign wire313 = forvar296;
  assign wire314 = ($unsigned(($unsigned(((8'ha2) >= reg288)) ?
                           wire276 : reg308[(4'hb):(2'h2)])) ?
                       {($unsigned(reg292) ?
                               forvar296 : (reg295 ?
                                   reg288 : (forvar281 > (8'hbf)))),
                           (~{$signed((8'hab)),
                               $unsigned(forvar281)})} : (^~$unsigned(reg306)));
  always
    @(posedge clk) begin
      reg315 = forvar303;
      reg316 <= $signed($signed((&(^~reg293))));
    end
  always
    @(posedge clk) begin
      reg317 <= (^(^(&($unsigned(reg279) ?
          $unsigned((8'h9f)) : $signed(reg315)))));
      reg318 = reg280[(4'hb):(4'h8)];
      reg319 = $signed((^~($unsigned((reg289 ? reg280 : reg309)) << ((8'hae) ?
          {reg301, reg301} : (forvar296 || reg295)))));
      reg320 = (~$signed((8'hb5)));
    end
  assign wire321 = (~|{wire313, reg319});
  always
    @(posedge clk) begin
      reg322 <= $unsigned(reg319[(1'h1):(1'h0)]);
      reg323 <= reg294;
    end
  always
    @(posedge clk) begin
      reg324 <= forvar282;
      reg325 = $signed((&($signed($unsigned(reg297)) ~^ reg311)));
      for (forvar326 = (1'h0); (forvar326 < (1'h0)); forvar326 = (forvar326 + (1'h1)))
        begin
          for (forvar327 = (1'h0); (forvar327 < (3'h4)); forvar327 = (forvar327 + (1'h1)))
            begin
              reg328 <= reg287;
              reg329 = (({(^{reg328, reg297})} ?
                  (~|((reg305 ?
                      reg320 : (8'hbb)) >> {reg286})) : (($unsigned((8'had)) ?
                      forvar304 : $unsigned(wire276)) >> $signed(reg293))) - $unsigned(reg306[(3'h6):(2'h3)]));
              reg330 <= (reg324 ?
                  $unsigned($unsigned(((^reg279) ?
                      (reg320 ^ reg324) : (~|(7'h43))))) : reg309);
            end
          reg331 <= ($signed((^~reg288[(3'h6):(3'h6)])) >>> reg315[(4'hd):(3'h5)]);
        end
    end
  always
    @(posedge clk) begin
      reg332 = reg301[(3'h6):(3'h5)];
      reg333 <= {forvar326,
          ($unsigned(forvar281[(1'h1):(1'h1)]) - reg332[(2'h3):(1'h0)])};
      for (forvar334 = (1'h0); (forvar334 < (2'h3)); forvar334 = (forvar334 + (1'h1)))
        begin
          reg335 <= $unsigned(reg332);
          reg336 <= $unsigned(reg305[(3'h5):(1'h1)]);
        end
    end
  always
    @(posedge clk) begin
      reg337 <= reg286[(3'h6):(2'h2)];
      reg338 = $signed((wire312[(4'h9):(4'h8)] >> (~({reg328} <<< $signed(wire278)))));
      reg339 <= ((+($unsigned((reg311 != (8'ha4))) ?
          ($signed(wire277) | (|reg301)) : wire276)) & reg286[(5'h11):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg340 <= (forvar334[(4'ha):(1'h0)] * $unsigned((reg323 == {wire277[(1'h1):(1'h1)]})));
      reg341 = ($signed(($unsigned($signed(reg331)) && forvar303[(1'h1):(1'h1)])) ?
          (7'h40) : {$unsigned($unsigned((~reg307))),
              ($signed((&reg310)) + {(+reg286), reg311[(3'h4):(1'h0)]})});
      reg342 <= reg310;
    end
endmodule