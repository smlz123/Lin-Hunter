(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h282):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire0;
  input wire [(5'h13):(1'h0)] wire1;
  input wire [(5'h12):(1'h0)] wire2;
  input wire [(4'hf):(1'h0)] wire3;
  wire [(2'h2):(1'h0)] wire694;
  wire signed [(4'hc):(1'h0)] wire4;
  wire [(4'ha):(1'h0)] wire5;
  wire signed [(5'h10):(1'h0)] wire6;
  reg signed [(5'h13):(1'h0)] reg7 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg8 = (1'h0);
  reg [(4'hc):(1'h0)] reg9 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire10;
  wire signed [(2'h3):(1'h0)] wire11;
  wire [(4'hf):(1'h0)] wire12;
  reg [(3'h7):(1'h0)] reg13 = (1'h0);
  reg [(4'hc):(1'h0)] forvar14 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg15 = (1'h0);
  reg [(5'h10):(1'h0)] reg16 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg17 = (1'h0);
  reg [(5'h11):(1'h0)] forvar18 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg20 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg21 = (1'h0);
  reg [(5'h13):(1'h0)] reg22 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg24 = (1'h0);
  reg [(4'h8):(1'h0)] reg25 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg26 = (1'h0);
  reg [(5'h14):(1'h0)] reg27 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar28 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg29 = (1'h0);
  reg [(5'h14):(1'h0)] reg30 = (1'h0);
  reg [(4'h8):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg33 = (1'h0);
  reg [(4'hc):(1'h0)] forvar34 = (1'h0);
  reg [(3'h5):(1'h0)] forvar35 = (1'h0);
  reg [(5'h13):(1'h0)] reg36 = (1'h0);
  reg [(5'h13):(1'h0)] reg37 = (1'h0);
  reg [(4'he):(1'h0)] reg38 = (1'h0);
  reg [(4'h8):(1'h0)] reg39 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg40 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg41 = (1'h0);
  reg [(5'h14):(1'h0)] reg42 = (1'h0);
  reg [(5'h10):(1'h0)] reg43 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar44 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg45 = (1'h0);
  reg [(5'h15):(1'h0)] reg46 = (1'h0);
  wire signed [(4'he):(1'h0)] wire47;
  wire [(5'h14):(1'h0)] wire48;
  wire signed [(3'h6):(1'h0)] wire49;
  wire [(2'h3):(1'h0)] wire692;
  assign y = {wire694,
                 wire4,
                 wire5,
                 wire6,
                 reg7,
                 reg8,
                 reg9,
                 wire10,
                 wire11,
                 wire12,
                 reg13,
                 forvar14,
                 reg15,
                 reg16,
                 reg17,
                 forvar18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 forvar28,
                 reg29,
                 reg30,
                 reg31,
                 reg32,
                 reg33,
                 forvar34,
                 forvar35,
                 reg36,
                 reg37,
                 reg38,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 forvar44,
                 reg45,
                 reg46,
                 wire47,
                 wire48,
                 wire49,
                 wire692,
                 (1'h0)};
  assign wire4 = (($unsigned(wire2) ?
                     (wire3[(4'hb):(3'h6)] ?
                         (!wire1[(2'h3):(1'h0)]) : (~|(+wire3))) : ((^$unsigned(wire0)) ?
                         (~|((7'h42) ?
                             wire1 : wire2)) : (+$unsigned(wire2)))) == $signed(($unsigned(((8'h9c) ?
                     wire3 : (8'ha6))) || $unsigned((wire2 | wire2)))));
  assign wire5 = $unsigned(((~^wire4) ? wire4[(3'h5):(3'h4)] : (!wire2)));
  assign wire6 = ($signed($signed(wire1)) ?
                     wire5[(1'h1):(1'h1)] : (^~(|($signed(wire4) ?
                         $signed((8'ha2)) : wire2))));
  always
    @(posedge clk) begin
      reg7 <= $unsigned((8'haf));
      reg8 = wire0[(4'hb):(4'ha)];
      reg9 <= (wire3 <= (((-wire0) ^ $unsigned((wire3 * wire5))) >> ((wire6 ?
              (wire2 - wire6) : $unsigned(wire6)) ?
          $signed($unsigned(wire1)) : {(wire0 ~^ wire5), reg7})));
    end
  assign wire10 = (reg8 ? (!wire0[(4'ha):(3'h4)]) : wire0);
  assign wire11 = wire10[(1'h1):(1'h1)];
  assign wire12 = wire11[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg13 <= reg9[(1'h1):(1'h0)];
      for (forvar14 = (1'h0); (forvar14 < (2'h3)); forvar14 = (forvar14 + (1'h1)))
        begin
          reg15 <= ($unsigned({reg8}) * $unsigned((^~(reg13 ?
              (wire12 ? reg7 : wire2) : (~|wire11)))));
          reg16 <= (wire5[(3'h7):(1'h0)] ?
              (reg15 ~^ $signed(wire3[(1'h0):(1'h0)])) : $signed(wire5));
          reg17 <= forvar14;
          for (forvar18 = (1'h0); (forvar18 < (3'h4)); forvar18 = (forvar18 + (1'h1)))
            begin
              reg19 <= (reg17 & wire11);
              reg20 <= $unsigned({($signed($signed(reg7)) >= (((8'hb8) ?
                      reg16 : wire5) ^~ (~&reg19)))});
              reg21 <= wire12;
              reg22 <= reg13[(3'h7):(3'h6)];
              reg23 = (~^$signed($signed(wire3[(4'h9):(4'h8)])));
            end
          reg24 <= (8'ha8);
        end
      if ((|(~|{($unsigned(reg7) & (+reg17)),
          (((8'ha4) ? wire1 : reg19) ? reg19 : ((8'hba) & wire1))})))
        begin
          reg25 = ($unsigned($signed(wire3)) != (~^{(^~(reg17 ?
                  (8'hbe) : (8'hba))),
              $unsigned((forvar18 > reg19))}));
        end
      else
        begin
          reg25 <= reg13;
          reg26 <= (($signed($signed($unsigned(reg25))) ?
                  (|reg8[(4'h9):(3'h6)]) : $unsigned($signed(((8'ha2) ?
                      wire4 : reg24)))) ?
              $signed(reg22) : $signed({(((8'h9f) >>> reg13) ?
                      (reg20 < (8'hbd)) : $unsigned(reg19))}));
          reg27 <= reg23[(4'h9):(2'h2)];
          for (forvar28 = (1'h0); (forvar28 < (2'h3)); forvar28 = (forvar28 + (1'h1)))
            begin
              reg29 = $unsigned(reg8[(5'h10):(4'hf)]);
              reg30 <= $signed(($unsigned(reg7) >> reg26));
              reg31 <= wire1[(1'h0):(1'h0)];
              reg32 <= reg29[(1'h0):(1'h0)];
              reg33 <= reg27;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar34 = (1'h0); (forvar34 < (1'h1)); forvar34 = (forvar34 + (1'h1)))
        begin
          for (forvar35 = (1'h0); (forvar35 < (2'h3)); forvar35 = (forvar35 + (1'h1)))
            begin
              reg36 <= (&$signed({reg20}));
              reg37 <= $signed($unsigned((8'ha7)));
              reg38 <= wire12;
              reg39 = reg15[(3'h5):(3'h4)];
              reg40 = (&forvar14[(2'h3):(1'h0)]);
            end
        end
      reg41 = $unsigned(wire0[(3'h4):(1'h0)]);
      reg42 <= ((~^$signed(reg26[(3'h5):(3'h4)])) ?
          (&(wire6 ?
              (reg40[(3'h4):(1'h0)] ?
                  $unsigned(reg8) : (^forvar35)) : (^(reg27 ?
                  reg13 : reg13)))) : $signed(wire3));
      reg43 <= reg23;
      for (forvar44 = (1'h0); (forvar44 < (1'h1)); forvar44 = (forvar44 + (1'h1)))
        begin
          reg45 = {({reg15, (~|(reg20 <= reg42))} ?
                  $signed(wire12[(4'hb):(3'h7)]) : (~^((forvar44 < forvar28) ?
                      reg37 : (~&reg43))))};
          reg46 = {(~|(^~(reg27 && reg43)))};
        end
    end
  assign wire47 = (reg27 > reg42);
  assign wire48 = reg32[(3'h7):(3'h5)];
  assign wire49 = $unsigned(((+wire3[(4'hb):(3'h7)]) ?
                      wire2[(4'ha):(3'h5)] : reg20[(2'h3):(2'h2)]));
  module50 modinst693 (wire692, clk, reg33, wire48, reg40, reg46, reg21);
  assign wire694 = ($unsigned(($signed($signed(reg16)) ?
                       reg7[(3'h6):(3'h6)] : $unsigned(reg31))) >> $unsigned(((wire692[(2'h2):(1'h1)] ?
                           (reg20 ? reg29 : reg19) : reg7[(5'h10):(4'hf)]) ?
                       (&wire0[(3'h5):(1'h0)]) : (wire10 ?
                           (forvar34 + (8'had)) : ((8'h9e) ? reg20 : reg16)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module50  (y, clk, wire55, wire54, wire53, wire52, wire51);
  output wire [(32'h2aa):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire55;
  input wire signed [(5'h12):(1'h0)] wire54;
  input wire [(5'h13):(1'h0)] wire53;
  input wire [(3'h6):(1'h0)] wire52;
  input wire signed [(4'hb):(1'h0)] wire51;
  wire [(4'hf):(1'h0)] wire691;
  reg signed [(4'hb):(1'h0)] reg690 = (1'h0);
  reg signed [(4'he):(1'h0)] reg689 = (1'h0);
  reg [(4'h9):(1'h0)] reg688 = (1'h0);
  reg [(5'h10):(1'h0)] reg687 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar686 = (1'h0);
  reg [(4'hd):(1'h0)] reg685 = (1'h0);
  reg [(4'hf):(1'h0)] reg684 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire683;
  reg [(4'hf):(1'h0)] reg682 = (1'h0);
  wire [(2'h3):(1'h0)] wire681;
  reg [(5'h13):(1'h0)] reg680 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg679 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg678 = (1'h0);
  reg [(5'h15):(1'h0)] reg677 = (1'h0);
  wire [(5'h14):(1'h0)] wire675;
  wire [(3'h5):(1'h0)] wire92;
  wire [(3'h6):(1'h0)] wire91;
  wire [(5'h12):(1'h0)] wire90;
  reg signed [(4'hd):(1'h0)] reg89 = (1'h0);
  reg [(4'hd):(1'h0)] reg88 = (1'h0);
  reg [(4'hf):(1'h0)] reg87 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg86 = (1'h0);
  reg [(4'ha):(1'h0)] forvar85 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg84 = (1'h0);
  reg [(4'h9):(1'h0)] forvar83 = (1'h0);
  reg [(4'hd):(1'h0)] reg82 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg81 = (1'h0);
  reg [(4'h8):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar78 = (1'h0);
  reg [(4'hd):(1'h0)] reg77 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar76 = (1'h0);
  wire [(5'h11):(1'h0)] wire75;
  wire [(4'hd):(1'h0)] wire74;
  reg [(5'h11):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg72 = (1'h0);
  reg [(4'hd):(1'h0)] reg71 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire70;
  wire signed [(2'h2):(1'h0)] wire69;
  reg [(3'h5):(1'h0)] reg68 = (1'h0);
  reg [(5'h13):(1'h0)] reg67 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg66 = (1'h0);
  reg [(5'h14):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg64 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg63 = (1'h0);
  reg [(5'h13):(1'h0)] forvar62 = (1'h0);
  reg [(3'h7):(1'h0)] forvar61 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg60 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg59 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar57 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg58 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg57 = (1'h0);
  reg [(5'h14):(1'h0)] reg56 = (1'h0);
  assign y = {wire691,
                 reg690,
                 reg689,
                 reg688,
                 reg687,
                 forvar686,
                 reg685,
                 reg684,
                 wire683,
                 reg682,
                 wire681,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 wire675,
                 wire92,
                 wire91,
                 wire90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 forvar85,
                 reg84,
                 forvar83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 forvar78,
                 reg77,
                 forvar76,
                 wire75,
                 wire74,
                 reg73,
                 reg72,
                 reg71,
                 wire70,
                 wire69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 forvar62,
                 forvar61,
                 reg60,
                 reg59,
                 forvar57,
                 reg58,
                 reg57,
                 reg56,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg56 <= wire55[(2'h3):(2'h3)];
      if ((($signed($unsigned(wire51[(4'h9):(3'h4)])) * (+wire52)) >= $signed({wire52,
          ({(8'hbc)} ^~ wire51[(3'h5):(3'h4)])})))
        begin
          reg57 = {(~wire55[(3'h7):(3'h5)])};
          reg58 = ($unsigned(wire54[(4'hd):(3'h7)]) || ($signed(((reg57 ?
              reg57 : wire53) >> (wire53 ?
              wire51 : (8'hb8)))) >> (+(~wire54))));
        end
      else
        begin
          for (forvar57 = (1'h0); (forvar57 < (2'h3)); forvar57 = (forvar57 + (1'h1)))
            begin
              reg58 = (((~^$signed($signed(wire53))) ? reg56 : forvar57) ?
                  (^~$unsigned($signed(wire53[(4'h9):(3'h6)]))) : $unsigned((forvar57[(3'h7):(3'h5)] <<< (8'ha0))));
            end
          reg59 = ($signed(reg58[(1'h0):(1'h0)]) ?
              {$unsigned((^$signed((8'hb6))))} : reg58);
        end
      reg60 = ($signed((|wire55)) ?
          (wire53 ?
              {wire55,
                  reg59[(1'h1):(1'h0)]} : wire55[(1'h0):(1'h0)]) : ($signed(((!reg57) | {wire51,
              wire54})) ~^ (wire51[(1'h1):(1'h0)] ?
              (-(reg56 ? forvar57 : (8'ha0))) : $unsigned((~&wire52)))));
      for (forvar61 = (1'h0); (forvar61 < (2'h2)); forvar61 = (forvar61 + (1'h1)))
        begin
          for (forvar62 = (1'h0); (forvar62 < (2'h3)); forvar62 = (forvar62 + (1'h1)))
            begin
              reg63 <= $unsigned($signed(($signed((reg59 ? reg58 : forvar57)) ?
                  {reg57[(3'h6):(3'h5)]} : ((wire52 > reg60) && (+reg59)))));
              reg64 <= $signed({{(!(wire51 ? wire51 : reg63))},
                  $signed($unsigned((+forvar62)))});
              reg65 <= ($signed(reg63) ?
                  (!reg60[(4'hb):(4'ha)]) : $signed(wire52));
              reg66 = $signed(reg59);
              reg67 = ((($signed($unsigned((8'hb3))) ?
                      reg66[(4'h9):(4'h9)] : {(&wire52),
                          wire51[(4'ha):(2'h2)]}) && reg63) ?
                  (((~|reg64) ?
                          ((8'haa) ?
                              wire53[(4'h8):(3'h7)] : reg65[(1'h1):(1'h0)]) : $unsigned(wire51[(2'h2):(1'h1)])) ?
                      $unsigned(($unsigned(reg59) ?
                          $unsigned(reg63) : $signed(wire51))) : (~|$signed(((8'h9e) || (8'hae))))) : reg63[(4'h8):(2'h2)]);
            end
        end
      reg68 <= (($signed($unsigned(forvar57)) ?
              (^$signed(reg60)) : (~^(^$unsigned((8'ha8))))) ?
          ($signed($unsigned(reg67)) - ((wire52 ?
                  forvar57[(3'h7):(2'h2)] : (reg60 ? reg66 : reg57)) ?
              ({reg65,
                  wire51} - $unsigned((8'hbf))) : $unsigned(reg58))) : wire51[(3'h6):(3'h4)]);
    end
  assign wire69 = $unsigned((reg56[(5'h14):(4'h9)] ?
                      (&{(forvar61 == reg57), reg63}) : reg58));
  assign wire70 = $signed((8'hb0));
  always
    @(posedge clk) begin
      reg71 = forvar62;
      reg72 <= reg65[(5'h13):(2'h3)];
      reg73 <= (-($unsigned({reg58}) ?
          forvar61[(1'h1):(1'h1)] : reg60[(5'h12):(4'hf)]));
    end
  assign wire74 = ((wire52[(3'h4):(1'h0)] | (|((reg60 + forvar62) * (reg59 ?
                      reg71 : wire55)))) <= ($unsigned($signed({reg64})) && $unsigned(wire55[(3'h6):(3'h6)])));
  assign wire75 = {{wire74,
                          (($signed(wire51) ?
                              {forvar57,
                                  wire51} : (wire70 >>> reg71)) >= $signed({reg66,
                              wire55}))},
                      $signed($signed(reg60[(2'h2):(1'h1)]))};
  always
    @(posedge clk) begin
      for (forvar76 = (1'h0); (forvar76 < (3'h4)); forvar76 = (forvar76 + (1'h1)))
        begin
          reg77 <= (forvar62 ? $signed($signed((|wire55))) : reg64);
          for (forvar78 = (1'h0); (forvar78 < (1'h1)); forvar78 = (forvar78 + (1'h1)))
            begin
              reg79 = ($signed($unsigned($unsigned(wire51))) - $signed(((8'h9f) >>> ($signed((8'ha8)) >> wire53[(5'h12):(1'h0)]))));
            end
          reg80 <= wire69[(1'h1):(1'h1)];
          reg81 <= $unsigned($signed($signed($signed({reg58}))));
        end
    end
  always
    @(posedge clk) begin
      reg82 = $unsigned($unsigned($signed(wire53)));
      for (forvar83 = (1'h0); (forvar83 < (3'h4)); forvar83 = (forvar83 + (1'h1)))
        begin
          reg84 = (|reg59[(4'ha):(4'h8)]);
          for (forvar85 = (1'h0); (forvar85 < (1'h1)); forvar85 = (forvar85 + (1'h1)))
            begin
              reg86 <= {$unsigned(reg56[(3'h4):(2'h2)])};
              reg87 <= ({(!$unsigned((reg56 ^ wire74)))} * ((8'hbb) ?
                  ($signed($signed(reg68)) ?
                      (8'hb4) : (^~reg77[(2'h2):(1'h0)])) : $unsigned($unsigned((reg65 <= wire54)))));
              reg88 <= (|(wire69[(1'h1):(1'h0)] ^ $signed($unsigned(reg81[(4'hc):(4'h8)]))));
              reg89 = ($unsigned($signed($signed($signed(reg68)))) ?
                  reg56 : $unsigned($signed(wire53[(4'h9):(3'h7)])));
            end
        end
    end
  assign wire90 = reg72;
  assign wire91 = (wire69[(2'h2):(2'h2)] + reg71[(4'ha):(3'h6)]);
  assign wire92 = wire52[(2'h2):(1'h0)];
  module93 modinst676 (.wire95(reg59), .clk(clk), .wire97(reg67), .wire96(reg72), .y(wire675), .wire94(reg89));
  always
    @(posedge clk) begin
      reg677 <= ({$signed($signed(reg67[(4'he):(3'h6)])),
          reg67} != (reg58[(2'h3):(2'h3)] ?
          (8'ha9) : $unsigned((reg71[(4'hc):(4'h9)] ?
              $signed((7'h41)) : wire70))));
      reg678 = (-$signed({{{reg67}}, reg60[(5'h13):(5'h12)]}));
      reg679 <= reg82[(2'h3):(1'h1)];
      reg680 = ($unsigned($signed(((!wire90) <<< ((8'h9c) ? wire51 : reg57)))) ?
          reg72[(1'h1):(1'h1)] : $signed(forvar61));
    end
  assign wire681 = $unsigned(($unsigned((8'ha9)) > {reg59[(1'h1):(1'h0)]}));
  always
    @(posedge clk) begin
      reg682 <= $unsigned((reg65 ?
          (|reg56) : ($unsigned({(8'ha3), reg88}) ?
              $unsigned((reg79 == (8'h9d))) : (~$unsigned(reg71)))));
    end
  assign wire683 = $signed($signed(wire681));
  always
    @(posedge clk) begin
      reg684 <= ((~($unsigned((~|reg679)) ?
          (reg71 || (|wire91)) : reg680[(3'h4):(1'h1)])) ~^ wire53[(4'h8):(3'h5)]);
    end
  always
    @(posedge clk) begin
      reg685 <= $signed((~&(~$signed((wire75 ? reg82 : wire675)))));
      for (forvar686 = (1'h0); (forvar686 < (2'h3)); forvar686 = (forvar686 + (1'h1)))
        begin
          reg687 <= wire54[(4'he):(2'h2)];
        end
      reg688 = $unsigned(((~{wire70[(2'h2):(2'h2)], {reg685}}) ?
          reg80[(3'h5):(3'h5)] : (reg59[(1'h0):(1'h0)] ?
              {$unsigned(forvar57),
                  (reg685 ?
                      (8'hbd) : (8'hb8))} : ((wire92 & reg86) - {forvar686,
                  reg56}))));
      reg689 = (~&(reg84 ? reg59[(2'h3):(2'h2)] : reg86));
      reg690 <= ($signed((~&(forvar686 << forvar61[(2'h2):(2'h2)]))) & (~&(reg60[(5'h12):(4'he)] & $signed(forvar686))));
    end
  assign wire691 = $unsigned(reg64[(2'h3):(1'h1)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module93
#( parameter param673 = (+(((((8'hbb) ? (8'ha4) : (8'hbf)) ? (|(8'h9d)) : (~(8'hab))) ? (~|(-(8'ha8))) : (((8'hbc) + (8'hbd)) ? ((8'hba) ? (8'hb0) : (8'hb2)) : ((8'hac) ? (8'hbd) : (8'ha2)))) ? (|(!(8'h9f))) : ((8'hbd) ? ({(8'hbe), (8'hb9)} && ((8'h9d) >>> (8'hb2))) : (~((7'h43) && (8'ha0))))))
, parameter param674 = param673 )
(y, clk, wire94, wire95, wire96, wire97);
  output wire [(32'h17d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire94;
  input wire signed [(4'h9):(1'h0)] wire95;
  input wire signed [(4'hf):(1'h0)] wire96;
  input wire [(5'h13):(1'h0)] wire97;
  wire [(3'h4):(1'h0)] wire672;
  reg [(4'h8):(1'h0)] reg671 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar670 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg669 = (1'h0);
  wire [(5'h13):(1'h0)] wire668;
  wire [(2'h3):(1'h0)] wire667;
  wire [(4'h8):(1'h0)] wire666;
  reg signed [(4'hb):(1'h0)] reg665 = (1'h0);
  reg [(3'h7):(1'h0)] reg664 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg663 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire662;
  wire [(5'h14):(1'h0)] wire661;
  wire [(5'h11):(1'h0)] wire660;
  wire signed [(5'h10):(1'h0)] wire659;
  reg [(4'he):(1'h0)] reg658 = (1'h0);
  reg [(5'h14):(1'h0)] reg657 = (1'h0);
  reg [(2'h2):(1'h0)] reg656 = (1'h0);
  reg [(5'h14):(1'h0)] reg655 = (1'h0);
  reg [(4'he):(1'h0)] reg654 = (1'h0);
  reg [(3'h6):(1'h0)] reg653 = (1'h0);
  reg [(4'hb):(1'h0)] reg652 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar651 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg651 = (1'h0);
  reg [(4'hb):(1'h0)] reg650 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg649 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg648 = (1'h0);
  wire [(5'h15):(1'h0)] wire646;
  wire signed [(3'h4):(1'h0)] wire541;
  wire signed [(4'hc):(1'h0)] wire98;
  wire [(5'h11):(1'h0)] wire99;
  wire signed [(5'h10):(1'h0)] wire539;
  assign y = {wire672,
                 reg671,
                 forvar670,
                 reg669,
                 wire668,
                 wire667,
                 wire666,
                 reg665,
                 reg664,
                 reg663,
                 wire662,
                 wire661,
                 wire660,
                 wire659,
                 reg658,
                 reg657,
                 reg656,
                 reg655,
                 reg654,
                 reg653,
                 reg652,
                 forvar651,
                 reg651,
                 reg650,
                 reg649,
                 reg648,
                 wire646,
                 wire541,
                 wire98,
                 wire99,
                 wire539,
                 (1'h0)};
  assign wire98 = {wire94, (wire94 > wire94)};
  assign wire99 = $signed(wire97);
  module100 modinst540 (wire539, clk, wire98, wire99, wire94, wire97, wire96);
  assign wire541 = {$signed(wire539),
                       (~|(wire96 ?
                           (~&{wire96}) : {wire96[(1'h0):(1'h0)],
                               ((8'hb8) >= wire539)}))};
  module542 modinst647 (wire646, clk, wire99, wire94, wire98, wire96);
  always
    @(posedge clk) begin
      reg648 <= (wire541[(1'h0):(1'h0)] ?
          ((^~wire541[(3'h4):(2'h3)]) >= wire541[(2'h2):(2'h2)]) : wire97);
      reg649 <= reg648;
    end
  always
    @(posedge clk) begin
      if ($signed((8'hb3)))
        begin
          reg650 <= $signed(wire541);
          reg651 <= ($signed($signed($unsigned((~wire96)))) ?
              $signed((((8'h9d) - $signed(wire95)) ?
                  reg648[(1'h0):(1'h0)] : ($signed(wire98) * $signed(reg649)))) : ($signed({(^reg648)}) ?
                  $signed((~|{wire646})) : $signed(wire98[(2'h3):(1'h0)])));
        end
      else
        begin
          reg650 = $unsigned($signed(reg650));
          for (forvar651 = (1'h0); (forvar651 < (2'h2)); forvar651 = (forvar651 + (1'h1)))
            begin
              reg652 <= reg649;
              reg653 = ($unsigned((!$signed(reg651))) ^ $signed($signed(((&wire95) ?
                  wire97[(4'hf):(1'h0)] : ((7'h44) <= wire98)))));
              reg654 <= forvar651[(3'h6):(3'h4)];
            end
          reg655 = ((reg649 ?
              $unsigned($signed((reg654 ?
                  reg653 : reg652))) : ((8'haf) ^ reg653[(3'h5):(3'h5)])) - reg649[(2'h3):(2'h3)]);
          reg656 = wire541;
          reg657 = $signed(wire96[(3'h7):(3'h5)]);
        end
      reg658 <= wire98;
    end
  assign wire659 = reg648[(3'h6):(1'h1)];
  assign wire660 = ($signed((!$unsigned((~|reg657)))) ? wire98 : reg658);
  assign wire661 = ((reg655[(2'h3):(1'h0)] ~^ reg648[(1'h1):(1'h1)]) ^ ((~|(8'ha4)) ?
                       (wire98[(1'h1):(1'h0)] <= wire646) : reg654[(4'h8):(2'h3)]));
  assign wire662 = (((&$signed($signed((8'hae)))) ? reg658 : wire94) ?
                       {((forvar651 + $unsigned(reg656)) | $signed(wire97[(4'h9):(2'h3)]))} : reg656);
  always
    @(posedge clk) begin
      reg663 <= (($signed($signed($signed(wire646))) << wire659[(3'h6):(3'h5)]) ?
          (&(reg654[(4'hc):(4'hc)] ?
              reg653 : (reg658[(1'h0):(1'h0)] ?
                  ((8'hae) ~^ wire98) : reg655))) : $signed((($unsigned(reg654) || (-wire661)) >= $unsigned(wire661))));
      reg664 <= (reg651[(1'h0):(1'h0)] ^ $signed((($signed(reg654) ?
              (^~wire94) : (reg655 & reg658)) ?
          {wire97} : reg652)));
      reg665 = reg648[(1'h1):(1'h1)];
    end
  assign wire666 = reg652[(1'h1):(1'h0)];
  assign wire667 = ((^~(({reg648} & wire541) ?
                       $unsigned((~|wire662)) : (wire99[(3'h4):(2'h2)] >= (&reg652)))) >= {wire661[(5'h10):(4'h8)],
                       $signed({reg665[(1'h1):(1'h1)]})});
  assign wire668 = ((~&(wire541 * (((8'hae) ? reg657 : reg652) + (reg651 ?
                           reg652 : (8'ha9))))) ?
                       $unsigned($signed((^wire666[(3'h5):(3'h4)]))) : reg649);
  always
    @(posedge clk) begin
      reg669 <= $signed(wire666[(1'h1):(1'h0)]);
      for (forvar670 = (1'h0); (forvar670 < (2'h2)); forvar670 = (forvar670 + (1'h1)))
        begin
          reg671 = $signed(reg651[(4'h8):(3'h6)]);
        end
    end
  assign wire672 = wire667[(1'h0):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module542
#( parameter param645 = ((-{((8'haf) ? (&(8'hb9)) : ((8'ha3) ? (8'hb2) : (8'ha0)))}) ? (^~((8'hbd) ? (((7'h43) ^ (8'hb9)) ? ((8'hb1) < (8'hac)) : {(8'hba)}) : ({(8'hbb), (8'h9c)} ? {(8'ha1), (7'h43)} : ((8'ha8) ? (8'hb6) : (8'ha7))))) : (((((7'h41) ? (8'hbf) : (7'h43)) ^~ ((8'hb2) && (8'hb7))) ? {(|(8'ha0)), (-(8'ha4))} : ((~|(8'ha4)) ? ((8'hab) && (8'ha5)) : ((8'hb1) ? (8'ha2) : (8'ha5)))) ? ((~((8'h9e) != (8'h9f))) == (~^{(8'ha2), (8'ha2)})) : (|({(8'hbf)} ? (^~(8'hae)) : {(8'h9e), (8'hb8)})))) )
(y, clk, wire546, wire545, wire544, wire543);
  output wire [(32'h45d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire546;
  input wire [(4'hd):(1'h0)] wire545;
  input wire [(4'hc):(1'h0)] wire544;
  input wire [(4'hf):(1'h0)] wire543;
  wire signed [(4'hf):(1'h0)] wire644;
  wire signed [(4'hc):(1'h0)] wire643;
  wire [(5'h12):(1'h0)] wire642;
  reg signed [(5'h15):(1'h0)] reg641 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg640 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg639 = (1'h0);
  reg [(3'h7):(1'h0)] reg638 = (1'h0);
  reg [(5'h11):(1'h0)] forvar637 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg636 = (1'h0);
  reg [(4'hd):(1'h0)] reg635 = (1'h0);
  reg [(3'h7):(1'h0)] reg634 = (1'h0);
  reg [(3'h5):(1'h0)] reg633 = (1'h0);
  reg [(5'h12):(1'h0)] forvar632 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg631 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg630 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg629 = (1'h0);
  reg [(3'h7):(1'h0)] reg628 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg627 = (1'h0);
  reg [(3'h7):(1'h0)] reg626 = (1'h0);
  reg [(5'h13):(1'h0)] reg625 = (1'h0);
  reg [(4'h9):(1'h0)] reg624 = (1'h0);
  reg [(3'h5):(1'h0)] reg623 = (1'h0);
  reg [(4'h9):(1'h0)] forvar622 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar621 = (1'h0);
  wire [(4'hc):(1'h0)] wire620;
  reg signed [(4'hf):(1'h0)] reg619 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg618 = (1'h0);
  reg [(2'h3):(1'h0)] reg617 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg616 = (1'h0);
  reg [(4'h9):(1'h0)] reg615 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg614 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg613 = (1'h0);
  reg [(5'h10):(1'h0)] forvar612 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg611 = (1'h0);
  reg signed [(4'he):(1'h0)] reg610 = (1'h0);
  reg [(3'h7):(1'h0)] reg609 = (1'h0);
  reg [(2'h2):(1'h0)] reg608 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg607 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar606 = (1'h0);
  reg [(5'h15):(1'h0)] reg605 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg604 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg603 = (1'h0);
  reg [(4'hb):(1'h0)] forvar602 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg601 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg600 = (1'h0);
  reg [(4'he):(1'h0)] reg599 = (1'h0);
  reg [(2'h3):(1'h0)] reg598 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar597 = (1'h0);
  reg [(3'h7):(1'h0)] reg596 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg595 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg594 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg593 = (1'h0);
  reg [(5'h13):(1'h0)] reg592 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg591 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar590 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg589 = (1'h0);
  reg [(5'h12):(1'h0)] reg588 = (1'h0);
  reg [(4'hc):(1'h0)] reg587 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg586 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg585 = (1'h0);
  reg [(3'h5):(1'h0)] reg584 = (1'h0);
  reg [(4'h8):(1'h0)] forvar583 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg582 = (1'h0);
  reg [(5'h10):(1'h0)] reg581 = (1'h0);
  reg [(4'hd):(1'h0)] reg580 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg579 = (1'h0);
  reg [(4'hd):(1'h0)] reg578 = (1'h0);
  reg [(3'h7):(1'h0)] reg577 = (1'h0);
  reg [(4'he):(1'h0)] reg576 = (1'h0);
  reg [(5'h13):(1'h0)] forvar575 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar574 = (1'h0);
  reg [(3'h4):(1'h0)] reg573 = (1'h0);
  reg [(4'hb):(1'h0)] reg572 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg571 = (1'h0);
  reg [(4'ha):(1'h0)] forvar570 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg569 = (1'h0);
  reg [(3'h5):(1'h0)] reg568 = (1'h0);
  reg signed [(4'he):(1'h0)] reg567 = (1'h0);
  reg [(3'h7):(1'h0)] reg566 = (1'h0);
  reg [(4'hd):(1'h0)] reg565 = (1'h0);
  reg [(4'hc):(1'h0)] reg564 = (1'h0);
  reg [(4'hd):(1'h0)] reg563 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg562 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire561;
  reg [(2'h3):(1'h0)] reg560 = (1'h0);
  wire [(4'h9):(1'h0)] wire559;
  reg signed [(5'h13):(1'h0)] reg558 = (1'h0);
  reg [(4'hd):(1'h0)] reg557 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg556 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg555 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg554 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg553 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg552 = (1'h0);
  reg signed [(4'he):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar550 = (1'h0);
  reg [(5'h10):(1'h0)] forvar549 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg548 = (1'h0);
  reg [(5'h12):(1'h0)] reg547 = (1'h0);
  assign y = {wire644,
                 wire643,
                 wire642,
                 reg641,
                 reg640,
                 reg639,
                 reg638,
                 forvar637,
                 reg636,
                 reg635,
                 reg634,
                 reg633,
                 forvar632,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 forvar622,
                 forvar621,
                 wire620,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 reg615,
                 reg614,
                 reg613,
                 forvar612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 forvar606,
                 reg605,
                 reg604,
                 reg603,
                 forvar602,
                 reg601,
                 reg600,
                 reg599,
                 reg598,
                 forvar597,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 forvar590,
                 reg589,
                 reg588,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 forvar583,
                 reg582,
                 reg581,
                 reg580,
                 reg579,
                 reg578,
                 reg577,
                 reg576,
                 forvar575,
                 forvar574,
                 reg573,
                 reg572,
                 reg571,
                 forvar570,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 reg565,
                 reg564,
                 reg563,
                 reg562,
                 wire561,
                 reg560,
                 wire559,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 reg551,
                 forvar550,
                 forvar549,
                 reg548,
                 reg547,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg547 <= wire546;
      reg548 <= (^(^(|wire544[(4'hb):(2'h3)])));
      for (forvar549 = (1'h0); (forvar549 < (1'h1)); forvar549 = (forvar549 + (1'h1)))
        begin
          for (forvar550 = (1'h0); (forvar550 < (1'h0)); forvar550 = (forvar550 + (1'h1)))
            begin
              reg551 <= (~|(-((^(forvar549 == forvar549)) ?
                  wire546[(3'h4):(2'h3)] : wire544)));
              reg552 <= $signed(wire544);
              reg553 <= wire543;
              reg554 = {$signed({wire543, reg551})};
              reg555 <= (((~reg548[(1'h1):(1'h1)]) >> (8'hbf)) ^ (~$unsigned((((8'hbd) ~^ reg552) ?
                  (forvar550 ? reg553 : (8'ha9)) : $unsigned((8'hb4))))));
            end
          reg556 <= (reg551 <= reg552);
          reg557 = (8'hb2);
        end
      reg558 = {(~|(|$unsigned($unsigned(reg556))))};
    end
  assign wire559 = ((reg557[(1'h1):(1'h0)] && reg547) ?
                       $signed($signed(wire545)) : ((({reg547} >> (8'h9c)) * $signed(((7'h44) ^~ (8'h9c)))) ?
                           ($signed((wire546 ?
                               forvar550 : wire544)) | $unsigned(reg554[(4'h9):(4'h8)])) : (!((reg555 ?
                                   wire546 : reg548) ?
                               reg547 : $unsigned(reg552)))));
  always
    @(posedge clk) begin
      reg560 = $unsigned((+(reg557[(3'h4):(2'h3)] < $unsigned((!reg547)))));
    end
  assign wire561 = (+((reg555 >>> (reg555[(1'h1):(1'h0)] ?
                       (reg551 ?
                           reg547 : wire543) : reg556)) < $signed((~$signed(wire559)))));
  always
    @(posedge clk) begin
      reg562 <= $unsigned({{reg558[(5'h13):(4'he)], $unsigned((|forvar549))}});
      reg563 = $signed(($unsigned((8'hbf)) ?
          wire545[(2'h2):(1'h0)] : (^$signed($unsigned(wire545)))));
      reg564 <= (({reg552[(2'h2):(2'h2)]} ?
          $signed($signed((reg560 >>> wire543))) : (reg551[(4'hc):(3'h5)] <<< $signed({forvar549}))) || reg552);
      reg565 <= reg553;
      reg566 <= $unsigned(($unsigned(reg565) ? reg548 : reg552[(2'h3):(2'h3)]));
    end
  always
    @(posedge clk) begin
      reg567 <= $unsigned(((wire561[(1'h1):(1'h0)] ?
          (reg552 ^ $signed(wire543)) : reg566) == $signed(reg551)));
      reg568 = (&(~((|(forvar550 ? reg556 : reg562)) == wire561)));
      reg569 <= wire543;
      for (forvar570 = (1'h0); (forvar570 < (1'h1)); forvar570 = (forvar570 + (1'h1)))
        begin
          reg571 = ({(7'h40)} ?
              {(^~$unsigned($unsigned(reg569))),
                  $unsigned(($signed(reg553) ?
                      $unsigned(wire545) : (wire546 < (8'hba))))} : (~^$signed(reg555)));
        end
    end
  always
    @(posedge clk) begin
      reg572 <= (7'h40);
      reg573 <= $signed(reg551);
      for (forvar574 = (1'h0); (forvar574 < (1'h1)); forvar574 = (forvar574 + (1'h1)))
        begin
          for (forvar575 = (1'h0); (forvar575 < (2'h2)); forvar575 = (forvar575 + (1'h1)))
            begin
              reg576 = $signed($signed($unsigned((^(|(8'hb6))))));
              reg577 <= {(^~$signed($unsigned({reg562, reg567}))),
                  (($unsigned(wire543) ?
                      ((!reg560) ?
                          $signed(wire546) : $signed((8'hab))) : (^~(-reg572))) & wire544[(1'h1):(1'h1)])};
              reg578 <= reg571;
              reg579 = {(&(8'hb9))};
              reg580 <= $signed(reg578[(4'h8):(2'h2)]);
            end
        end
      reg581 <= ($signed(reg571) ?
          ($unsigned((8'hb1)) >> reg578) : $unsigned(forvar575[(5'h10):(4'hc)]));
    end
  always
    @(posedge clk) begin
      reg582 = (8'hab);
      for (forvar583 = (1'h0); (forvar583 < (1'h0)); forvar583 = (forvar583 + (1'h1)))
        begin
          reg584 <= {(($signed($signed(reg557)) * (~reg582[(4'h9):(3'h6)])) ~^ $unsigned($signed((~^wire544)))),
              reg581[(4'hc):(3'h5)]};
          reg585 <= (~&(!(reg557[(3'h5):(2'h3)] ~^ $unsigned(reg568))));
          reg586 <= {(reg571 ?
                  $unsigned(reg554[(3'h6):(1'h0)]) : (reg558 && reg567[(4'h9):(2'h2)])),
              reg555};
          reg587 <= (({(8'ha1),
                  (wire559[(4'h8):(3'h6)] ?
                      $signed((8'hb1)) : $signed(reg567))} ^~ (((|reg566) ?
                  (reg564 ?
                      wire559 : reg578) : {reg557}) >= {$signed(wire543)})) ?
              reg566 : ($signed($signed(reg565[(2'h3):(1'h0)])) ?
                  reg552 : $signed(($unsigned(reg566) ?
                      reg571[(1'h0):(1'h0)] : reg562[(4'ha):(3'h4)]))));
        end
      reg588 <= {reg580};
      reg589 = ($unsigned($unsigned((-{reg562, (8'h9d)}))) ?
          $unsigned((~{$unsigned((8'hb3)),
              reg556})) : $signed({{reg585[(3'h7):(2'h2)]},
              {$signed(wire546), (forvar583 * reg581)}}));
    end
  always
    @(posedge clk) begin
      for (forvar590 = (1'h0); (forvar590 < (1'h0)); forvar590 = (forvar590 + (1'h1)))
        begin
          reg591 <= (wire544 ?
              $signed($unsigned($unsigned((~^reg563)))) : $signed($signed(reg567)));
          reg592 = ({(~|reg551[(4'hc):(2'h3)]), $signed((^(^~reg578)))} ?
              $signed($unsigned(wire559)) : (|($unsigned((~forvar575)) ?
                  (reg547 | (&reg567)) : $signed(((8'had) ?
                      (8'ha4) : (8'ha5))))));
          reg593 <= reg591[(4'hc):(3'h6)];
          reg594 <= forvar550;
          reg595 <= ({((reg591[(2'h2):(2'h2)] << reg572) ?
                      ((reg569 >= reg556) < reg589[(1'h0):(1'h0)]) : $signed(wire559[(4'h8):(3'h7)]))} ?
              (reg582 < forvar550[(4'hc):(3'h6)]) : $unsigned(reg587));
        end
      reg596 <= (wire561[(1'h0):(1'h0)] + ($signed(((reg591 >> reg553) ?
              $signed(reg557) : $signed(reg572))) ?
          $signed(reg551[(4'hc):(4'ha)]) : (+(7'h42))));
      for (forvar597 = (1'h0); (forvar597 < (3'h4)); forvar597 = (forvar597 + (1'h1)))
        begin
          reg598 <= forvar550[(4'hb):(2'h2)];
          reg599 <= (~|{($unsigned(reg563[(3'h5):(2'h2)]) ^ $unsigned((8'hb3)))});
          reg600 = $unsigned(reg557);
          reg601 <= {$signed(reg560[(1'h1):(1'h1)]),
              $unsigned($signed(((reg573 ?
                  reg553 : reg578) || (reg547 ^ forvar590))))};
          for (forvar602 = (1'h0); (forvar602 < (3'h4)); forvar602 = (forvar602 + (1'h1)))
            begin
              reg603 <= (wire546 & {reg566,
                  $unsigned(($unsigned(reg573) ^~ {reg598}))});
              reg604 = (reg576 >>> (reg596[(1'h0):(1'h0)] ?
                  (8'hb1) : forvar570));
            end
        end
      reg605 = $unsigned((&(reg548[(2'h2):(1'h0)] ?
          $signed($unsigned(forvar597)) : reg599[(2'h2):(1'h1)])));
      for (forvar606 = (1'h0); (forvar606 < (2'h2)); forvar606 = (forvar606 + (1'h1)))
        begin
          reg607 = ($signed((&$signed((~|forvar575)))) | reg592);
          reg608 <= reg563;
          reg609 <= $signed({$signed((reg571 || $unsigned(reg566)))});
          reg610 <= ((+(reg568 ?
              (reg562 || (7'h42)) : ($signed(reg593) ?
                  forvar602 : $signed((8'haf))))) < {((reg565 ^~ {reg604,
                  (7'h43)}) ^ (~^(reg609 ^ reg573))),
              (|{forvar570[(3'h5):(2'h2)]})});
          reg611 = ((8'ha5) > reg610[(4'hd):(4'hd)]);
        end
    end
  always
    @(posedge clk) begin
      for (forvar612 = (1'h0); (forvar612 < (2'h2)); forvar612 = (forvar612 + (1'h1)))
        begin
          reg613 <= $unsigned((|forvar612[(4'he):(4'ha)]));
          reg614 <= $signed((8'ha6));
          reg615 <= reg607[(3'h5):(1'h0)];
          reg616 <= ($signed($unsigned($unsigned($signed(reg555)))) ?
              (reg593[(1'h0):(1'h0)] ?
                  ($unsigned(reg566) > forvar570) : reg565[(3'h4):(2'h2)]) : ($unsigned($signed(reg579[(4'hb):(1'h1)])) - forvar606[(2'h3):(1'h0)]));
          reg617 <= reg567;
        end
      reg618 <= (reg610[(1'h0):(1'h0)] ?
          (^$unsigned(reg576[(4'ha):(2'h3)])) : (reg609[(1'h1):(1'h0)] >> reg609[(3'h5):(3'h4)]));
    end
  always
    @(posedge clk) begin
      reg619 <= (8'ha7);
    end
  assign wire620 = (reg615[(2'h3):(1'h1)] < (8'hbf));
  always
    @(posedge clk) begin
      for (forvar621 = (1'h0); (forvar621 < (1'h0)); forvar621 = (forvar621 + (1'h1)))
        begin
          for (forvar622 = (1'h0); (forvar622 < (1'h0)); forvar622 = (forvar622 + (1'h1)))
            begin
              reg623 <= $signed(($unsigned({reg578}) | $unsigned($signed($signed(reg618)))));
              reg624 = forvar621[(3'h4):(1'h0)];
              reg625 = {$signed({(|wire561)})};
            end
          if ((reg577[(3'h5):(3'h5)] ?
              {forvar574,
                  $unsigned($signed(((8'ha7) > reg610)))} : (&(|{(wire543 ?
                      reg580 : reg618)}))))
            begin
              reg626 <= reg601[(4'h8):(3'h4)];
              reg627 <= (8'ha1);
              reg628 <= (^({(8'hbb),
                  ($signed(forvar621) ?
                      {forvar570, reg562} : {reg564})} < {($signed(forvar575) ?
                      {wire559, forvar570} : $unsigned(reg552))}));
              reg629 <= ((~&reg562[(1'h1):(1'h0)]) ?
                  $signed(reg568[(3'h5):(2'h3)]) : ((($signed(reg615) << $unsigned(reg593)) ?
                          {((8'ha8) ? (8'ha6) : reg567),
                              $unsigned(reg599)} : (|(reg585 ?
                              reg615 : reg593))) ?
                      $signed($signed((8'haa))) : $signed({(forvar575 ?
                              wire561 : reg596),
                          (reg577 ? reg599 : wire561)})));
              reg630 = (~&(|{((reg610 < reg589) ?
                      (reg557 >> reg593) : $unsigned(reg624)),
                  $signed((forvar597 == reg548))}));
            end
          else
            begin
              reg626 <= {(reg616 ?
                      ((reg608 >>> (reg626 ?
                          reg604 : reg605)) && reg582[(4'h8):(4'h8)]) : reg623[(2'h3):(1'h0)])};
            end
          reg631 <= reg551[(2'h2):(1'h1)];
          for (forvar632 = (1'h0); (forvar632 < (2'h2)); forvar632 = (forvar632 + (1'h1)))
            begin
              reg633 <= reg595[(3'h6):(1'h0)];
              reg634 = forvar612[(3'h4):(1'h0)];
              reg635 <= ($signed(({reg564[(3'h7):(3'h5)]} || reg615)) < {(reg614[(1'h1):(1'h0)] ?
                      $signed(reg625[(5'h12):(3'h4)]) : wire620)});
            end
        end
      reg636 <= (8'ha9);
      for (forvar637 = (1'h0); (forvar637 < (2'h3)); forvar637 = (forvar637 + (1'h1)))
        begin
          reg638 <= $unsigned((&(!$unsigned($unsigned((8'hb6))))));
          reg639 = {($unsigned((-(reg603 && (8'hae)))) ?
                  $unsigned({(reg558 ?
                          forvar602 : reg562)}) : $unsigned($signed((reg627 + reg584))))};
          reg640 <= $signed((((reg569 ?
                  (wire543 ^~ reg580) : (forvar612 || forvar570)) - (!(|(8'ha7)))) ?
              ($signed((8'hbd)) ?
                  ((reg633 <= reg551) ?
                      reg587[(3'h4):(1'h1)] : $unsigned(reg614)) : (8'ha3)) : ((^$signed(reg557)) & $signed((^reg555)))));
        end
      reg641 <= $signed(reg605[(5'h14):(4'hd)]);
    end
  assign wire642 = $signed(reg633);
  assign wire643 = {reg568};
  assign wire644 = $unsigned({reg576[(3'h5):(3'h5)],
                       {((reg560 ^ forvar622) >> (!(8'hb7)))}});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module100  (y, clk, wire105, wire104, wire103, wire102, wire101);
  output wire [(32'h2df):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire105;
  input wire [(5'h11):(1'h0)] wire104;
  input wire [(4'h8):(1'h0)] wire103;
  input wire signed [(5'h13):(1'h0)] wire102;
  input wire signed [(2'h2):(1'h0)] wire101;
  reg signed [(2'h2):(1'h0)] reg538 = (1'h0);
  reg [(5'h15):(1'h0)] reg537 = (1'h0);
  reg [(5'h14):(1'h0)] reg536 = (1'h0);
  reg [(4'hf):(1'h0)] reg535 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire534;
  reg signed [(3'h7):(1'h0)] reg533 = (1'h0);
  reg [(5'h10):(1'h0)] reg532 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg531 = (1'h0);
  reg [(4'he):(1'h0)] reg530 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar529 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire528;
  reg signed [(3'h7):(1'h0)] reg527 = (1'h0);
  reg [(4'hd):(1'h0)] reg526 = (1'h0);
  reg [(2'h2):(1'h0)] forvar525 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg524 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg523 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg522 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar521 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg520 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg519 = (1'h0);
  reg [(3'h5):(1'h0)] forvar518 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg517 = (1'h0);
  reg [(4'h8):(1'h0)] reg516 = (1'h0);
  reg [(5'h10):(1'h0)] reg515 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg514 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg513 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar512 = (1'h0);
  reg [(4'h9):(1'h0)] reg511 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg510 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg509 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg508 = (1'h0);
  wire [(4'h9):(1'h0)] wire507;
  reg [(4'hf):(1'h0)] reg506 = (1'h0);
  reg [(3'h6):(1'h0)] reg505 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg504 = (1'h0);
  reg [(4'hf):(1'h0)] reg503 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg502 = (1'h0);
  wire [(2'h2):(1'h0)] wire382;
  reg signed [(3'h4):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar130 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg129 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg128 = (1'h0);
  reg [(3'h4):(1'h0)] forvar127 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg126 = (1'h0);
  wire [(2'h3):(1'h0)] wire125;
  wire signed [(4'hf):(1'h0)] wire124;
  reg signed [(4'he):(1'h0)] reg123 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg122 = (1'h0);
  reg [(3'h4):(1'h0)] reg121 = (1'h0);
  reg [(4'hb):(1'h0)] reg120 = (1'h0);
  reg [(4'h9):(1'h0)] reg119 = (1'h0);
  reg [(3'h4):(1'h0)] reg118 = (1'h0);
  reg [(4'hd):(1'h0)] reg117 = (1'h0);
  reg [(4'hd):(1'h0)] reg116 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg115 = (1'h0);
  reg [(2'h2):(1'h0)] reg114 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg113 = (1'h0);
  reg [(5'h10):(1'h0)] forvar112 = (1'h0);
  reg [(5'h13):(1'h0)] reg111 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg109 = (1'h0);
  reg [(5'h15):(1'h0)] forvar108 = (1'h0);
  reg [(3'h7):(1'h0)] forvar107 = (1'h0);
  wire [(5'h13):(1'h0)] wire106;
  wire signed [(4'h8):(1'h0)] wire384;
  wire [(5'h13):(1'h0)] wire385;
  wire signed [(3'h4):(1'h0)] wire386;
  wire [(4'hd):(1'h0)] wire500;
  assign y = {reg538,
                 reg537,
                 reg536,
                 reg535,
                 wire534,
                 reg533,
                 reg532,
                 reg531,
                 reg530,
                 forvar529,
                 wire528,
                 reg527,
                 reg526,
                 forvar525,
                 reg524,
                 reg523,
                 reg522,
                 forvar521,
                 reg520,
                 reg519,
                 forvar518,
                 reg517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 forvar512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 wire507,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 wire382,
                 reg131,
                 forvar130,
                 reg129,
                 reg128,
                 forvar127,
                 reg126,
                 wire125,
                 wire124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 forvar112,
                 reg111,
                 reg110,
                 reg109,
                 forvar108,
                 forvar107,
                 wire106,
                 wire384,
                 wire385,
                 wire386,
                 wire500,
                 (1'h0)};
  assign wire106 = $unsigned((~(+((!wire105) ? (+wire104) : (~^wire103)))));
  always
    @(posedge clk) begin
      for (forvar107 = (1'h0); (forvar107 < (1'h0)); forvar107 = (forvar107 + (1'h1)))
        begin
          for (forvar108 = (1'h0); (forvar108 < (2'h2)); forvar108 = (forvar108 + (1'h1)))
            begin
              reg109 <= $unsigned($unsigned($unsigned(wire104)));
              reg110 = (($unsigned((reg109[(4'hd):(3'h5)] ?
                  ((8'ha2) ?
                      wire103 : forvar107) : (wire105 || reg109))) > $unsigned($signed((forvar108 < reg109)))) ^~ {wire102});
              reg111 <= (wire101[(1'h0):(1'h0)] ?
                  (reg109[(1'h0):(1'h0)] ?
                      forvar108[(4'hb):(1'h0)] : (|{((8'hab) & wire102),
                          (wire105 <= wire102)})) : $unsigned($unsigned(((wire101 ?
                          (8'hae) : forvar108) ?
                      (wire101 ? wire105 : (8'had)) : (forvar107 ?
                          wire102 : wire104)))));
            end
          for (forvar112 = (1'h0); (forvar112 < (3'h4)); forvar112 = (forvar112 + (1'h1)))
            begin
              reg113 = ({$unsigned($unsigned($unsigned(wire105)))} ?
                  ((!((-reg109) <= (^forvar108))) >> $signed(((reg110 < wire106) ?
                      (reg111 ?
                          wire103 : forvar108) : $signed(forvar108)))) : $unsigned(wire105[(2'h2):(1'h1)]));
              reg114 <= $signed($signed(((wire101 ?
                      $signed(wire104) : (-reg111)) ?
                  ($unsigned(wire103) ?
                      $unsigned(wire103) : $signed(forvar108)) : $signed({wire101,
                      wire102}))));
              reg115 = (^$unsigned(reg109[(4'ha):(2'h2)]));
              reg116 <= reg109;
              reg117 = wire101;
            end
          reg118 <= $unsigned(wire101);
          reg119 <= (~reg115[(1'h1):(1'h1)]);
        end
      reg120 <= (forvar108 < {(-$signed((|reg110)))});
      reg121 <= ($unsigned($unsigned(($unsigned(wire104) * $signed(reg115)))) ?
          reg117 : reg118);
    end
  always
    @(posedge clk) begin
      reg122 <= ((reg118[(1'h1):(1'h1)] != {(8'hb8), (8'h9d)}) ?
          forvar112 : (+(|{wire105[(1'h1):(1'h0)], {wire101, reg117}})));
      reg123 = (+reg116);
    end
  assign wire124 = wire104[(3'h6):(2'h2)];
  assign wire125 = (reg115[(4'h9):(3'h5)] ?
                       (reg118[(2'h3):(2'h2)] ?
                           (($signed(wire102) == $signed(reg115)) ?
                               reg115 : wire124) : ($unsigned(reg123) ^~ ((reg118 ?
                                   reg117 : forvar107) ?
                               (~(8'h9f)) : (reg123 ?
                                   (8'h9d) : forvar108)))) : ({reg114[(2'h2):(1'h1)],
                               (((8'ha7) ? reg116 : reg111) ?
                                   reg118 : $unsigned(reg113))} ?
                           $signed($unsigned((wire104 & reg123))) : reg111[(2'h2):(2'h2)]));
  always
    @(posedge clk) begin
      reg126 <= $unsigned((|$signed((+$signed(reg109)))));
      for (forvar127 = (1'h0); (forvar127 < (2'h3)); forvar127 = (forvar127 + (1'h1)))
        begin
          reg128 <= {$unsigned($signed(reg122)),
              ($unsigned((|{forvar112, reg114})) != reg110[(3'h4):(2'h2)])};
          reg129 <= $signed((reg114[(1'h0):(1'h0)] ~^ ($signed($signed(reg115)) ?
              (8'hb8) : ((8'hbd) ^ (forvar127 ^ reg115)))));
        end
      for (forvar130 = (1'h0); (forvar130 < (2'h2)); forvar130 = (forvar130 + (1'h1)))
        begin
          reg131 <= reg118[(3'h4):(2'h3)];
        end
    end
  module132 modinst383 (wire382, clk, reg111, forvar130, forvar108, reg128, reg126);
  assign wire384 = (8'ha5);
  assign wire385 = $unsigned(wire106[(1'h1):(1'h1)]);
  assign wire386 = reg111[(4'hb):(3'h6)];
  module387 modinst501 (wire500, clk, forvar112, wire124, reg115, wire384, wire385);
  always
    @(posedge clk) begin
      reg502 <= $signed($unsigned((reg116 ?
          (((8'hb5) ? forvar108 : reg118) ?
              $unsigned(forvar107) : (wire103 ?
                  reg128 : reg117)) : $unsigned(wire125[(2'h2):(1'h0)]))));
      reg503 <= (reg110 <= ($unsigned({$unsigned(wire106)}) != ({(reg121 ?
              forvar130 : wire101),
          reg123[(4'hb):(3'h6)]} ~^ $unsigned(wire500))));
      reg504 <= (^~(reg128 != ($unsigned(reg115) || ((-reg116) ?
          (forvar127 ? reg119 : reg111) : reg128[(1'h1):(1'h1)]))));
      reg505 = ($signed($signed((8'ha8))) + (^forvar107));
      reg506 <= (~^(((7'h41) ?
          $unsigned(wire386[(1'h1):(1'h1)]) : $signed(wire101[(2'h2):(1'h1)])) - {{((8'hb3) ?
                  reg111 : wire125),
              $signed(wire103)}}));
    end
  assign wire507 = wire103[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg508 = (-$signed({(&reg119), $signed({wire103})}));
      reg509 <= (wire125 && (~((+forvar108) ?
          $signed((wire103 | reg508)) : (!{wire105}))));
      if (reg113)
        begin
          reg510 = (8'hac);
          reg511 <= reg503[(3'h4):(3'h4)];
          for (forvar512 = (1'h0); (forvar512 < (2'h2)); forvar512 = (forvar512 + (1'h1)))
            begin
              reg513 <= (&(wire382[(1'h1):(1'h0)] == wire382));
              reg514 = reg121[(1'h0):(1'h0)];
              reg515 <= $signed(($signed(reg116) ?
                  {$unsigned((reg117 <<< reg503)), (-(~reg120))} : (((^reg113) ?
                      reg116 : $signed(forvar127)) >> {$signed(reg118),
                      $unsigned(reg113)})));
              reg516 <= wire125;
              reg517 <= $signed($signed(($unsigned((reg505 & reg117)) ?
                  reg510 : (~&(reg114 ? reg128 : wire106)))));
            end
          for (forvar518 = (1'h0); (forvar518 < (2'h3)); forvar518 = (forvar518 + (1'h1)))
            begin
              reg519 <= reg115;
              reg520 = ((($unsigned($signed(wire382)) ?
                      (-reg109[(5'h12):(4'h9)]) : wire382[(2'h2):(1'h0)]) >>> {wire104,
                      $signed((^(8'hb6)))}) ?
                  (!wire384[(1'h1):(1'h1)]) : $signed($signed((&(reg113 && reg122)))));
            end
          for (forvar521 = (1'h0); (forvar521 < (2'h3)); forvar521 = (forvar521 + (1'h1)))
            begin
              reg522 <= $signed((8'hb9));
              reg523 <= $signed($signed((7'h41)));
            end
        end
      else
        begin
          reg510 <= (8'hab);
        end
      reg524 <= reg520[(1'h0):(1'h0)];
      for (forvar525 = (1'h0); (forvar525 < (2'h2)); forvar525 = (forvar525 + (1'h1)))
        begin
          reg526 <= (|$unsigned(((~reg510[(1'h0):(1'h0)]) ?
              $unsigned({(7'h43), reg113}) : ($signed((8'h9c)) >>> reg506))));
          reg527 <= $signed({((~(reg508 >= forvar127)) ^~ ((!(8'ha3)) | wire101[(2'h2):(2'h2)])),
              ($unsigned((-wire102)) ^ ($signed((8'hbe)) <= reg508[(4'h9):(1'h1)]))});
        end
    end
  assign wire528 = $signed({{{$signed(reg524)}, $signed((~(8'ha3)))}});
  always
    @(posedge clk) begin
      for (forvar529 = (1'h0); (forvar529 < (2'h2)); forvar529 = (forvar529 + (1'h1)))
        begin
          reg530 = reg510[(2'h3):(2'h2)];
        end
      reg531 <= $unsigned($unsigned((({reg116,
              reg516} || (wire384 >>> (8'ha2))) ?
          ($signed((8'ha4)) ^ reg519) : $signed($signed(reg111)))));
      reg532 <= {($unsigned(((~^reg131) ?
              $signed(reg510) : ((8'hbc) & (7'h40)))) != reg510[(1'h1):(1'h0)])};
      reg533 <= $unsigned($unsigned($unsigned(forvar525[(1'h1):(1'h1)])));
    end
  assign wire534 = reg126[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg535 <= ($unsigned((^reg129[(2'h2):(1'h0)])) ?
          $unsigned(($signed({forvar130}) && $signed((~(8'ha1))))) : ($unsigned((~&$unsigned(forvar127))) & {$signed((reg123 > reg129)),
              {reg524[(2'h3):(2'h2)], (wire534 ? wire384 : forvar112)}}));
      reg536 = reg514[(3'h4):(1'h0)];
      reg537 <= (((wire102[(4'ha):(3'h6)] << ({forvar521, wire382} ?
              $signed(wire124) : (~&reg531))) ?
          (8'hab) : $signed(wire507[(3'h7):(3'h6)])) - ($unsigned(($signed(wire386) <<< (8'ha0))) <= $signed($unsigned(reg502[(4'h9):(3'h5)]))));
      reg538 <= reg111;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module387
#( parameter param499 = (~^(^~{(((8'hb9) ^ (8'ha4)) > ((8'hbc) ? (7'h43) : (8'hb7))), ((!(8'h9e)) ? ((7'h44) ? (7'h43) : (8'hb5)) : ((8'ha2) >= (8'hb0)))})) )
(y, clk, wire392, wire391, wire390, wire389, wire388);
  output wire [(32'h264):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire392;
  input wire signed [(4'hf):(1'h0)] wire391;
  input wire [(4'h8):(1'h0)] wire390;
  input wire [(3'h4):(1'h0)] wire389;
  input wire [(4'he):(1'h0)] wire388;
  reg signed [(4'he):(1'h0)] reg498 = (1'h0);
  reg [(5'h14):(1'h0)] reg497 = (1'h0);
  reg [(5'h14):(1'h0)] reg496 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg495 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg494 = (1'h0);
  wire [(4'hf):(1'h0)] wire493;
  reg [(2'h3):(1'h0)] reg492 = (1'h0);
  reg [(5'h11):(1'h0)] reg491 = (1'h0);
  reg [(5'h13):(1'h0)] reg490 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg489 = (1'h0);
  reg [(4'ha):(1'h0)] reg488 = (1'h0);
  reg [(5'h15):(1'h0)] reg487 = (1'h0);
  reg [(5'h10):(1'h0)] reg486 = (1'h0);
  reg [(5'h12):(1'h0)] forvar485 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg484 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg483 = (1'h0);
  reg [(5'h10):(1'h0)] reg482 = (1'h0);
  reg [(3'h5):(1'h0)] reg481 = (1'h0);
  reg [(2'h2):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar479 = (1'h0);
  reg [(5'h11):(1'h0)] reg478 = (1'h0);
  reg [(4'h9):(1'h0)] forvar477 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg476 = (1'h0);
  reg [(2'h2):(1'h0)] reg475 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg474 = (1'h0);
  reg [(4'hb):(1'h0)] reg473 = (1'h0);
  reg [(3'h7):(1'h0)] forvar472 = (1'h0);
  reg [(3'h7):(1'h0)] reg471 = (1'h0);
  reg [(5'h15):(1'h0)] forvar470 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg469 = (1'h0);
  reg [(3'h5):(1'h0)] reg468 = (1'h0);
  reg [(2'h3):(1'h0)] reg467 = (1'h0);
  reg [(5'h10):(1'h0)] reg466 = (1'h0);
  reg [(4'h9):(1'h0)] reg465 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg464 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg463 = (1'h0);
  reg [(5'h15):(1'h0)] reg462 = (1'h0);
  reg [(4'hd):(1'h0)] reg461 = (1'h0);
  reg [(3'h7):(1'h0)] reg460 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire459;
  reg [(5'h13):(1'h0)] reg458 = (1'h0);
  reg [(5'h11):(1'h0)] reg457 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg456 = (1'h0);
  reg [(5'h13):(1'h0)] reg455 = (1'h0);
  reg [(5'h14):(1'h0)] reg454 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire453;
  wire [(3'h4):(1'h0)] wire452;
  wire signed [(4'ha):(1'h0)] wire451;
  wire signed [(4'hd):(1'h0)] wire449;
  wire [(4'h9):(1'h0)] wire393;
  assign y = {reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 wire493,
                 reg492,
                 reg491,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 forvar485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 forvar479,
                 reg478,
                 forvar477,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 forvar472,
                 reg471,
                 forvar470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 wire459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 wire453,
                 wire452,
                 wire451,
                 wire449,
                 wire393,
                 (1'h0)};
  assign wire393 = {wire388[(1'h1):(1'h0)]};
  module394 modinst450 (.wire397(wire392), .wire398(wire393), .wire395(wire388), .wire396(wire391), .clk(clk), .y(wire449));
  assign wire451 = wire393;
  assign wire452 = wire388[(2'h3):(2'h2)];
  assign wire453 = (+wire390[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg454 <= wire391;
      reg455 <= $signed($signed($unsigned((~|$unsigned(reg454)))));
      reg456 <= (($signed((+(+wire449))) != ((&((8'hb6) ? wire390 : wire388)) ?
              {wire452} : (!(&reg454)))) ?
          wire391 : (((8'h9d) | wire453[(1'h1):(1'h1)]) ?
              $signed($unsigned(wire389)) : (~^wire390)));
      reg457 <= (({(&(wire392 ?
              reg454 : (8'ha5)))} << ($signed((~|wire452)) >> $signed($unsigned(wire392)))) + (^wire389[(1'h1):(1'h0)]));
      reg458 = ((|$signed((-wire451[(3'h7):(3'h5)]))) << $signed(($signed((wire453 ?
              wire453 : wire393)) ?
          (reg455 ?
              (wire388 ?
                  (8'ha9) : wire452) : (wire391 <<< (7'h42))) : {(&wire452),
              (reg457 >= reg457)})));
    end
  assign wire459 = wire449;
  always
    @(posedge clk) begin
      reg460 <= reg456[(3'h7):(1'h1)];
      reg461 <= (reg455 ?
          wire392[(4'hd):(2'h3)] : $signed((($unsigned(reg456) << (8'hae)) ^ {(wire393 && reg458)})));
    end
  always
    @(posedge clk) begin
      reg462 <= {{$signed(((~^wire449) < wire389)),
              $unsigned($unsigned(reg461))}};
      reg463 <= reg454;
      reg464 <= (~^$signed(($signed(reg463[(3'h4):(2'h3)]) != $signed((wire451 ?
          reg461 : wire393)))));
      reg465 <= $signed(wire453);
      reg466 <= $unsigned(reg455[(2'h2):(2'h2)]);
    end
  always
    @(posedge clk) begin
      reg467 <= $signed(($signed($signed(reg456[(3'h5):(3'h5)])) ?
          reg460 : (wire451[(3'h5):(3'h5)] + wire449[(1'h0):(1'h0)])));
      reg468 = ({reg467[(1'h0):(1'h0)]} | reg467[(1'h0):(1'h0)]);
      reg469 = (~|{(8'h9e), $signed(wire459)});
      for (forvar470 = (1'h0); (forvar470 < (3'h4)); forvar470 = (forvar470 + (1'h1)))
        begin
          reg471 = reg463;
          for (forvar472 = (1'h0); (forvar472 < (1'h1)); forvar472 = (forvar472 + (1'h1)))
            begin
              reg473 <= (~|$unsigned($unsigned(wire393)));
              reg474 = (($unsigned($signed((~&wire388))) & ($unsigned($signed(reg461)) ?
                      (^$signed(wire451)) : ((~wire391) ?
                          (~|reg464) : $unsigned(wire393)))) ?
                  reg461 : (forvar470 ^ (~(wire452 ?
                      reg468 : (reg456 ~^ wire391)))));
            end
          reg475 <= $signed(((^~$signed((|wire459))) ^ (reg454[(4'h9):(2'h3)] ?
              $unsigned($unsigned(wire392)) : (~{wire391}))));
          reg476 <= ($unsigned((-reg457)) >> wire453);
        end
      for (forvar477 = (1'h0); (forvar477 < (1'h0)); forvar477 = (forvar477 + (1'h1)))
        begin
          reg478 <= ((8'h9c) ?
              reg469[(1'h0):(1'h0)] : (reg467[(2'h3):(1'h1)] ?
                  wire393 : ($unsigned($signed(reg466)) <<< {(wire389 ?
                          forvar472 : reg465)})));
          for (forvar479 = (1'h0); (forvar479 < (1'h1)); forvar479 = (forvar479 + (1'h1)))
            begin
              reg480 <= (^~(~reg468[(3'h4):(2'h2)]));
              reg481 = {$unsigned(reg476[(4'hb):(4'ha)])};
              reg482 <= $unsigned({(!$signed(forvar472))});
              reg483 <= reg478;
            end
          reg484 <= ((reg469 ? reg468[(3'h5):(3'h4)] : reg475[(1'h1):(1'h1)]) ?
              {wire390[(3'h6):(1'h1)],
                  (~^(8'hb5))} : ($signed(reg483[(4'h9):(3'h6)]) >>> {{(&reg462)},
                  $unsigned(wire449)}));
          for (forvar485 = (1'h0); (forvar485 < (1'h0)); forvar485 = (forvar485 + (1'h1)))
            begin
              reg486 <= $signed(reg454);
              reg487 <= $unsigned($signed($signed(wire390[(3'h4):(1'h1)])));
              reg488 <= $unsigned(reg478);
              reg489 <= forvar485[(1'h0):(1'h0)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg490 = $unsigned((reg482 ?
          $unsigned(reg468) : ($unsigned((forvar470 ? forvar470 : (8'ha1))) ?
              $unsigned((wire391 >> wire392)) : $unsigned((wire392 ?
                  forvar485 : reg489)))));
      reg491 = forvar485[(4'h9):(3'h7)];
      reg492 <= $unsigned(reg483);
    end
  assign wire493 = reg490;
  always
    @(posedge clk) begin
      reg494 <= (!{$unsigned(forvar485[(5'h12):(3'h7)])});
      reg495 <= wire451;
      reg496 = $unsigned($signed(reg490[(4'hb):(3'h7)]));
      reg497 <= (~|$signed((~(~(8'haf)))));
      reg498 <= (forvar477[(4'h9):(3'h4)] & ((reg469 <= ({(8'ha5)} * {reg455,
          wire451})) ~^ ((-$signed((8'ha8))) ?
          reg471 : $signed($signed((8'ha6))))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module132
#( parameter param380 = {(((((8'haa) && (8'haf)) ? (~&(7'h41)) : ((8'h9d) | (8'ha0))) >> ((|(8'ha0)) ^~ (|(7'h40)))) != {(((7'h43) ? (8'ha5) : (8'hb4)) ? (&(8'h9c)) : ((8'ha3) ? (8'h9c) : (8'hb5))), {((7'h43) == (8'had)), ((8'ha6) ? (8'hb5) : (8'hb8))}}), (~^{(~&((7'h43) ? (8'hb5) : (8'hb1))), {((8'h9f) ^~ (8'ha6)), {(8'hab), (8'hbb)}}})}
, parameter param381 = param380 )
(y, clk, wire133, wire134, wire135, wire136, wire137);
  output wire [(32'ha1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire133;
  input wire signed [(5'h14):(1'h0)] wire134;
  input wire [(5'h13):(1'h0)] wire135;
  input wire [(4'ha):(1'h0)] wire136;
  input wire [(3'h6):(1'h0)] wire137;
  wire [(2'h2):(1'h0)] wire378;
  wire signed [(2'h3):(1'h0)] wire310;
  reg signed [(5'h15):(1'h0)] reg138 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg139 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire140;
  reg [(4'hb):(1'h0)] reg141 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire142;
  wire signed [(3'h5):(1'h0)] wire200;
  wire signed [(5'h11):(1'h0)] wire246;
  wire signed [(5'h11):(1'h0)] wire248;
  wire signed [(5'h15):(1'h0)] wire249;
  wire signed [(4'hd):(1'h0)] wire308;
  assign y = {wire378,
                 wire310,
                 reg138,
                 reg139,
                 wire140,
                 reg141,
                 wire142,
                 wire200,
                 wire246,
                 wire248,
                 wire249,
                 wire308,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg138 <= (wire135[(3'h5):(2'h3)] ?
          $unsigned((|(~|$signed((8'hb2))))) : (-$unsigned(wire135)));
      reg139 <= wire137;
    end
  assign wire140 = $unsigned($unsigned((((wire133 ? (8'hbf) : wire134) ?
                       (wire134 <<< reg139) : (wire137 * wire135)) + $signed(wire136))));
  always
    @(posedge clk) begin
      reg141 <= ($signed(wire133[(4'h9):(3'h7)]) && wire137);
    end
  assign wire142 = (8'hb9);
  module143 modinst201 (.wire144(wire142), .wire147(reg139), .y(wire200), .wire146(wire133), .wire145(wire134), .clk(clk));
  module202 modinst247 (.clk(clk), .y(wire246), .wire203(wire140), .wire204(wire134), .wire205(wire142), .wire206(wire135));
  assign wire248 = ($unsigned(reg141) ?
                       wire136 : (|$unsigned(($signed(reg139) ?
                           wire142 : (wire137 < wire137)))));
  assign wire249 = wire137;
  module250 modinst309 (wire308, clk, reg139, wire246, wire135, wire248, wire137);
  assign wire310 = ($signed(reg141[(3'h7):(3'h4)]) ?
                       $unsigned($unsigned(wire135)) : $unsigned($unsigned($signed({(8'hb2)}))));
  module311 modinst379 (.wire312(wire308), .wire315(reg138), .wire314(reg139), .y(wire378), .clk(clk), .wire313(wire248));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module311  (y, clk, wire315, wire314, wire313, wire312);
  output wire [(32'h307):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire315;
  input wire signed [(5'h10):(1'h0)] wire314;
  input wire signed [(5'h10):(1'h0)] wire313;
  input wire [(2'h2):(1'h0)] wire312;
  reg [(2'h3):(1'h0)] reg377 = (1'h0);
  reg [(5'h11):(1'h0)] reg376 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg375 = (1'h0);
  reg [(4'hc):(1'h0)] reg374 = (1'h0);
  reg [(2'h2):(1'h0)] reg373 = (1'h0);
  reg [(3'h4):(1'h0)] reg372 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg371 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg370 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg369 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg368 = (1'h0);
  reg [(5'h12):(1'h0)] forvar367 = (1'h0);
  reg [(4'hd):(1'h0)] reg366 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg365 = (1'h0);
  reg signed [(4'he):(1'h0)] reg364 = (1'h0);
  reg [(3'h7):(1'h0)] reg363 = (1'h0);
  reg [(4'ha):(1'h0)] forvar362 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar361 = (1'h0);
  wire [(3'h7):(1'h0)] wire360;
  reg signed [(4'hd):(1'h0)] reg359 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg358 = (1'h0);
  reg [(5'h13):(1'h0)] reg357 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire356;
  reg [(5'h10):(1'h0)] reg355 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg354 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg353 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg352 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg351 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg350 = (1'h0);
  reg signed [(4'he):(1'h0)] reg349 = (1'h0);
  reg [(5'h15):(1'h0)] forvar348 = (1'h0);
  reg [(3'h7):(1'h0)] reg347 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg346 = (1'h0);
  reg [(5'h15):(1'h0)] forvar345 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg344 = (1'h0);
  wire [(5'h13):(1'h0)] wire343;
  reg signed [(3'h7):(1'h0)] reg342 = (1'h0);
  reg [(5'h11):(1'h0)] reg341 = (1'h0);
  reg [(4'he):(1'h0)] reg340 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg339 = (1'h0);
  reg signed [(4'he):(1'h0)] reg338 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire337;
  reg signed [(5'h13):(1'h0)] reg331 = (1'h0);
  reg signed [(4'he):(1'h0)] reg336 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg335 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg333 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg332 = (1'h0);
  reg [(4'hf):(1'h0)] forvar331 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg330 = (1'h0);
  reg [(4'hd):(1'h0)] reg329 = (1'h0);
  reg [(5'h15):(1'h0)] reg328 = (1'h0);
  reg [(5'h11):(1'h0)] reg327 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg326 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg325 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar324 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg323 = (1'h0);
  reg [(4'hb):(1'h0)] reg322 = (1'h0);
  reg [(5'h15):(1'h0)] reg321 = (1'h0);
  reg [(4'hf):(1'h0)] forvar320 = (1'h0);
  reg [(4'hd):(1'h0)] reg319 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire318;
  wire signed [(5'h11):(1'h0)] wire317;
  wire signed [(5'h10):(1'h0)] wire316;
  assign y = {reg377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 forvar367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 forvar362,
                 forvar361,
                 wire360,
                 reg359,
                 reg358,
                 reg357,
                 wire356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 reg350,
                 reg349,
                 forvar348,
                 reg347,
                 reg346,
                 forvar345,
                 reg344,
                 wire343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 wire337,
                 reg331,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 forvar331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 forvar324,
                 reg323,
                 reg322,
                 reg321,
                 forvar320,
                 reg319,
                 wire318,
                 wire317,
                 wire316,
                 (1'h0)};
  assign wire316 = $signed($unsigned((((wire312 || wire314) ?
                           $unsigned(wire313) : wire314) ?
                       (^((8'hab) ?
                           wire313 : wire314)) : wire312[(2'h2):(1'h1)])));
  assign wire317 = (wire315[(4'h9):(4'h8)] <= $signed(wire315));
  assign wire318 = wire312;
  always
    @(posedge clk) begin
      reg319 <= wire313[(2'h3):(2'h2)];
      for (forvar320 = (1'h0); (forvar320 < (1'h0)); forvar320 = (forvar320 + (1'h1)))
        begin
          reg321 <= wire315;
          reg322 <= $signed(($signed((!(^wire317))) && wire312));
          reg323 <= $unsigned(((8'hb4) >>> reg319[(4'ha):(3'h4)]));
          for (forvar324 = (1'h0); (forvar324 < (2'h2)); forvar324 = (forvar324 + (1'h1)))
            begin
              reg325 <= reg319[(4'hc):(2'h3)];
              reg326 <= wire316[(2'h2):(2'h2)];
              reg327 = ((~&$signed((((8'hb8) >> reg323) >> (^~wire317)))) - $signed(wire318[(4'h8):(1'h1)]));
              reg328 <= reg327;
            end
          reg329 <= $unsigned((~|reg322));
        end
      reg330 <= $unsigned((8'hbc));
      if (reg326[(3'h4):(3'h4)])
        begin
          for (forvar331 = (1'h0); (forvar331 < (2'h2)); forvar331 = (forvar331 + (1'h1)))
            begin
              reg332 = reg323[(2'h3):(2'h2)];
              reg333 <= $unsigned((8'hb1));
              reg334 <= reg327;
              reg335 = ({reg327[(4'hf):(4'hd)]} != (reg322 != ((^~$unsigned((7'h41))) ?
                  $unsigned((reg334 >>> reg334)) : ($unsigned(wire317) ^ $signed(wire316)))));
              reg336 <= (&(({(+reg333)} << reg329[(4'h9):(3'h7)]) || $signed({(reg322 >>> reg334),
                  $signed(reg325)})));
            end
        end
      else
        begin
          reg331 <= (reg328 ?
              ((-$signed(forvar320)) ?
                  forvar324 : (~|(^{wire316,
                      forvar331}))) : ($unsigned(wire313) && (^((wire318 && (8'h9f)) | (reg321 ?
                  (7'h44) : (8'haa))))));
          reg332 <= ({(((^reg321) ? reg329[(4'hb):(3'h4)] : $signed(reg327)) ?
                      $signed((reg336 ^ forvar331)) : (&$signed(wire317))),
                  (((reg333 ? forvar331 : reg326) >> (reg328 ?
                          reg332 : reg319)) ?
                      (&{wire317, reg319}) : $unsigned((~|reg327)))} ?
              (($unsigned($unsigned((8'hb5))) ?
                  $signed(((7'h41) ?
                      reg329 : wire312)) : {(|(8'had))}) ^~ ($signed((~&forvar331)) ^ ($signed(reg329) ?
                  $unsigned((8'hb9)) : $signed(wire316)))) : ((8'haa) << $signed(wire312[(1'h1):(1'h0)])));
          reg333 <= ((~^(((reg325 ? reg334 : wire312) && ((7'h44) ?
              wire313 : wire316)) < $signed($signed(reg335)))) >> ($signed(($unsigned(reg327) << $signed(reg323))) >= $signed(wire312[(1'h1):(1'h1)])));
          reg334 = $signed(wire317);
          reg335 <= (((|$unsigned((wire313 ?
                  forvar320 : wire317))) >>> $signed((^~$unsigned(reg326)))) ?
              $signed(reg325[(3'h4):(2'h3)]) : (8'ha3));
        end
    end
  assign wire337 = (+($unsigned(((wire315 ? reg334 : reg331) <= (&reg322))) ?
                       (reg326[(3'h6):(2'h3)] <= {wire317[(3'h7):(2'h2)],
                           (wire317 ? forvar331 : reg335)}) : (8'hae)));
  always
    @(posedge clk) begin
      reg338 = (|((~(~(+wire337))) ?
          (!$signed((&(8'hbb)))) : (~&((|reg336) * $signed((8'hbe))))));
      reg339 <= ($unsigned({(wire313 ? reg325 : wire313)}) ?
          reg334[(3'h7):(3'h6)] : wire313);
      reg340 = $signed(($unsigned((~|reg326)) ~^ $unsigned(((reg334 ?
              reg327 : reg336) ?
          (wire314 - reg328) : reg338[(2'h2):(1'h1)]))));
      reg341 <= reg326;
      reg342 <= reg326[(1'h1):(1'h1)];
    end
  assign wire343 = ($unsigned((~&reg338)) ^~ {({{(7'h40)}} ?
                           (+$signed(wire318)) : (wire316[(2'h2):(1'h0)] ?
                               $unsigned(forvar320) : (reg331 | (8'hbf)))),
                       $signed((+reg321))});
  always
    @(posedge clk) begin
      reg344 <= ((+(((8'ha8) << $unsigned(reg338)) ?
              ((reg339 ? wire313 : reg325) ?
                  wire317[(3'h5):(3'h4)] : {reg334,
                      reg331}) : (-reg332[(2'h3):(1'h1)]))) ?
          {(-$signed((-forvar331)))} : forvar324);
      for (forvar345 = (1'h0); (forvar345 < (1'h1)); forvar345 = (forvar345 + (1'h1)))
        begin
          reg346 <= (wire315 != $signed(wire316));
          reg347 <= ($signed(reg338[(4'he):(3'h4)]) ^ $unsigned((($signed((8'ha9)) ?
                  {reg322, reg340} : {reg344}) ?
              $unsigned($signed(reg335)) : (wire312[(1'h1):(1'h1)] <<< reg332))));
          for (forvar348 = (1'h0); (forvar348 < (2'h2)); forvar348 = (forvar348 + (1'h1)))
            begin
              reg349 = $unsigned(($signed({$unsigned(reg336)}) ^~ $unsigned((&(!reg342)))));
              reg350 = $signed((((~&reg342[(2'h3):(1'h1)]) - reg323) ^ ({$unsigned(forvar324)} ?
                  (~|(^reg347)) : (reg349[(4'h8):(3'h6)] ~^ wire314))));
              reg351 <= $signed(reg347);
              reg352 = reg323;
              reg353 <= (({(reg338 ? wire312[(1'h1):(1'h0)] : reg352),
                  (-(wire313 & reg333))} << (~&reg331[(3'h5):(2'h3)])) || ($unsigned(wire314) ?
                  (wire315[(4'h8):(3'h6)] ?
                      reg350 : ({reg321} ?
                          {reg321, (8'hba)} : $signed(reg325))) : reg327));
            end
          reg354 <= wire343[(2'h2):(1'h1)];
          reg355 = (!reg344);
        end
    end
  assign wire356 = ({(((&wire337) & (&forvar345)) <= ($unsigned(reg347) != (reg342 ?
                               wire343 : reg341))),
                           ({(reg321 ? wire313 : reg353)} >>> wire312)} ?
                       $signed((wire314 ? reg349 : $signed(reg339))) : reg347);
  always
    @(posedge clk) begin
      reg357 <= forvar348[(1'h0):(1'h0)];
      reg358 <= $signed($signed(wire315[(1'h0):(1'h0)]));
      reg359 <= {wire315};
    end
  assign wire360 = reg354;
  always
    @(posedge clk) begin
      for (forvar361 = (1'h0); (forvar361 < (3'h4)); forvar361 = (forvar361 + (1'h1)))
        begin
          for (forvar362 = (1'h0); (forvar362 < (2'h3)); forvar362 = (forvar362 + (1'h1)))
            begin
              reg363 <= (((~(forvar361 ?
                  $unsigned((8'hbd)) : wire315)) & (($unsigned(reg332) ?
                  (reg332 >> reg340) : (wire316 < reg352)) ^ ($unsigned(reg335) ?
                  (~&reg336) : $signed(forvar324)))) + reg328[(5'h12):(4'hc)]);
              reg364 <= (wire313[(3'h4):(2'h2)] ?
                  (-{wire360}) : $signed($signed((&(reg332 ?
                      reg341 : wire312)))));
            end
          reg365 <= {$unsigned((reg334[(3'h6):(2'h3)] != ({reg325,
                  reg364} >> (forvar320 ? reg331 : wire314)))),
              {$unsigned((^$signed(wire313)))}};
          reg366 <= (~(~&$unsigned((~&reg331[(1'h0):(1'h0)]))));
        end
      for (forvar367 = (1'h0); (forvar367 < (2'h3)); forvar367 = (forvar367 + (1'h1)))
        begin
          reg368 <= (({(8'ha1)} != $unsigned(((forvar324 ?
              wire312 : (8'ha3)) - (^reg319)))) < reg331[(5'h11):(4'h9)]);
          reg369 <= forvar348[(4'hd):(2'h3)];
          reg370 <= ((~|{forvar361,
              (reg342 * {reg349,
                  wire343})}) - ($signed((reg364 != (~|reg327))) << reg351));
        end
    end
  always
    @(posedge clk) begin
      reg371 <= $unsigned(reg365);
      reg372 <= $signed((~^forvar324[(1'h1):(1'h0)]));
      reg373 = $signed(({$unsigned((reg327 ? forvar361 : forvar324))} ?
          reg331[(3'h6):(1'h0)] : reg340[(2'h3):(2'h2)]));
      reg374 <= $signed($unsigned((reg340[(3'h6):(2'h3)] ~^ (8'hba))));
      reg375 = reg373;
    end
  always
    @(posedge clk) begin
      reg376 <= reg340;
      reg377 <= (~|{(reg363[(2'h3):(1'h1)] || (~&(reg344 ? reg325 : reg338))),
          (8'had)});
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module250
#( parameter param307 = ({(((^(8'had)) ? ((8'ha9) < (7'h41)) : ((7'h40) & (7'h43))) <= (-((8'hb1) <= (8'ha8))))} >>> ((8'ha1) >> {(((8'ha0) ? (8'hb2) : (8'hb4)) ? {(8'hb8)} : ((8'ha3) > (8'hb2)))})) )
(y, clk, wire255, wire254, wire253, wire252, wire251);
  output wire [(32'h27b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire255;
  input wire [(4'he):(1'h0)] wire254;
  input wire signed [(5'h13):(1'h0)] wire253;
  input wire signed [(5'h11):(1'h0)] wire252;
  input wire signed [(2'h2):(1'h0)] wire251;
  wire signed [(5'h14):(1'h0)] wire306;
  reg [(5'h12):(1'h0)] reg305 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg304 = (1'h0);
  reg [(4'hd):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg302 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg301 = (1'h0);
  reg [(4'he):(1'h0)] reg300 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire299;
  wire [(2'h3):(1'h0)] wire298;
  wire [(4'he):(1'h0)] wire297;
  reg signed [(4'hd):(1'h0)] reg296 = (1'h0);
  reg [(4'he):(1'h0)] reg295 = (1'h0);
  reg [(4'hd):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg293 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg292 = (1'h0);
  reg [(3'h4):(1'h0)] reg291 = (1'h0);
  reg [(4'h9):(1'h0)] reg290 = (1'h0);
  reg [(5'h11):(1'h0)] reg289 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg288 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg287 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg286 = (1'h0);
  reg [(5'h15):(1'h0)] reg285 = (1'h0);
  reg [(3'h6):(1'h0)] reg284 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar283 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar282 = (1'h0);
  reg [(5'h13):(1'h0)] reg281 = (1'h0);
  wire [(5'h11):(1'h0)] wire280;
  reg signed [(4'hb):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg278 = (1'h0);
  reg [(4'hf):(1'h0)] reg277 = (1'h0);
  reg [(3'h6):(1'h0)] forvar276 = (1'h0);
  reg [(3'h4):(1'h0)] reg275 = (1'h0);
  reg [(4'hd):(1'h0)] reg274 = (1'h0);
  reg [(2'h2):(1'h0)] reg273 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar272 = (1'h0);
  reg [(4'h9):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg270 = (1'h0);
  reg [(3'h5):(1'h0)] reg269 = (1'h0);
  reg [(4'hf):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar267 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg266 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg265 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg264 = (1'h0);
  reg [(4'h9):(1'h0)] forvar263 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg262 = (1'h0);
  wire [(4'hb):(1'h0)] wire261;
  wire signed [(5'h11):(1'h0)] wire260;
  wire [(3'h6):(1'h0)] wire259;
  reg [(4'h9):(1'h0)] reg258 = (1'h0);
  reg [(4'hb):(1'h0)] reg257 = (1'h0);
  reg [(5'h11):(1'h0)] reg256 = (1'h0);
  assign y = {wire306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 wire299,
                 wire298,
                 wire297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 forvar283,
                 forvar282,
                 reg281,
                 wire280,
                 reg279,
                 reg278,
                 reg277,
                 forvar276,
                 reg275,
                 reg274,
                 reg273,
                 forvar272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 forvar267,
                 reg266,
                 reg265,
                 reg264,
                 forvar263,
                 reg262,
                 wire261,
                 wire260,
                 wire259,
                 reg258,
                 reg257,
                 reg256,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg256 = (wire252[(4'hf):(4'hf)] << $signed(({$signed(wire252), wire251} ?
          {((7'h44) ? wire255 : wire252),
              wire253[(2'h3):(1'h0)]} : (~&wire253[(5'h11):(5'h11)]))));
      reg257 <= ((8'hb0) ? (^wire254) : $signed((|wire251[(1'h1):(1'h0)])));
      reg258 <= wire251;
    end
  assign wire259 = (&$unsigned(wire254[(1'h1):(1'h1)]));
  assign wire260 = {wire259, reg256};
  assign wire261 = reg256[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg262 <= wire251[(2'h2):(2'h2)];
      for (forvar263 = (1'h0); (forvar263 < (1'h1)); forvar263 = (forvar263 + (1'h1)))
        begin
          reg264 = forvar263;
        end
      reg265 <= reg257[(2'h2):(1'h1)];
      reg266 <= wire253[(5'h11):(4'ha)];
      for (forvar267 = (1'h0); (forvar267 < (2'h2)); forvar267 = (forvar267 + (1'h1)))
        begin
          reg268 <= ((((+(!wire254)) ?
                  reg265[(3'h4):(2'h2)] : $signed((^forvar267))) == (forvar267[(5'h10):(4'h8)] || ((wire261 != wire254) | (-(8'hb1))))) ?
              (~|(8'h9f)) : reg257[(4'h8):(3'h7)]);
          reg269 <= ((7'h43) ? (8'hb8) : $unsigned($unsigned(forvar267)));
          reg270 <= forvar267;
        end
    end
  always
    @(posedge clk) begin
      reg271 <= $signed(reg266[(3'h5):(1'h0)]);
      for (forvar272 = (1'h0); (forvar272 < (2'h2)); forvar272 = (forvar272 + (1'h1)))
        begin
          reg273 <= (!wire255);
          reg274 <= $signed(wire261[(2'h2):(1'h0)]);
          reg275 <= wire253;
          for (forvar276 = (1'h0); (forvar276 < (2'h3)); forvar276 = (forvar276 + (1'h1)))
            begin
              reg277 = (~|((8'ha7) ?
                  {({reg273} <= (forvar267 & (8'h9e))),
                      reg264[(4'h8):(3'h5)]} : reg264));
              reg278 <= $unsigned((~^{$signed((wire261 ? wire260 : reg270)),
                  (8'hb2)}));
              reg279 = reg264;
            end
        end
    end
  assign wire280 = ($signed($signed((~|(8'hb5)))) == ((&($signed(wire252) != (^reg262))) >= wire255));
  always
    @(posedge clk) begin
      reg281 <= (~&((!((wire255 ? (8'hbb) : reg278) * (wire280 ?
              reg271 : reg269))) ?
          (((!(7'h43)) ? $unsigned(wire255) : $signed(reg279)) ?
              reg257[(3'h7):(2'h3)] : (reg258 ?
                  {forvar272} : $unsigned(reg277))) : (({reg257} - $signed(wire254)) & $signed((reg266 ?
              reg266 : reg269)))));
      for (forvar282 = (1'h0); (forvar282 < (3'h4)); forvar282 = (forvar282 + (1'h1)))
        begin
          for (forvar283 = (1'h0); (forvar283 < (2'h2)); forvar283 = (forvar283 + (1'h1)))
            begin
              reg284 <= {wire254[(3'h4):(3'h4)]};
              reg285 = $unsigned(((-wire261[(2'h2):(1'h0)]) < (~|((^wire261) > forvar272[(3'h6):(2'h2)]))));
              reg286 = reg269[(3'h4):(1'h1)];
              reg287 <= $signed({reg264, $unsigned((!$signed(reg278)))});
            end
          reg288 = {$unsigned((~^reg268[(3'h4):(2'h3)])), reg279};
          reg289 <= {($signed($signed(wire261[(1'h0):(1'h0)])) ?
                  (8'ha7) : {{reg288[(3'h5):(1'h1)]}}),
              {((^$signed(forvar263)) | reg278[(3'h4):(2'h2)]),
                  $unsigned(($unsigned(reg262) <= $signed(reg257)))}};
        end
      reg290 <= $unsigned(reg274[(1'h1):(1'h0)]);
      reg291 <= forvar276[(2'h2):(1'h1)];
      reg292 <= $signed(reg286);
    end
  always
    @(posedge clk) begin
      reg293 <= (reg287 ? $unsigned(reg287) : forvar263[(4'h8):(2'h3)]);
      reg294 <= ((((~|(reg274 * (8'hab))) != reg258) ? (&reg269) : {wire254}) ?
          reg265[(3'h6):(3'h6)] : (~$unsigned(reg281)));
      reg295 <= reg265;
      reg296 = $unsigned((wire260 ^~ (~|$unsigned(((8'h9f) ?
          reg278 : reg294)))));
    end
  assign wire297 = (8'hbb);
  assign wire298 = reg268[(2'h3):(2'h2)];
  assign wire299 = $signed($unsigned(((|$unsigned(reg258)) ?
                       (!wire253[(3'h4):(1'h0)]) : ($signed(reg281) ?
                           {(8'hbd), reg287} : (reg258 ^~ reg264)))));
  always
    @(posedge clk) begin
      reg300 <= $unsigned(($unsigned(reg291) ? wire261 : $unsigned((8'ha0))));
      reg301 <= (~&wire255[(1'h1):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg302 <= (wire260 | ($signed(($unsigned(reg285) * reg300[(4'hd):(4'hc)])) ?
          $signed(((^~wire252) < reg295[(4'hb):(3'h4)])) : (wire259[(2'h3):(2'h3)] <= ($signed(wire255) >>> reg292[(4'hc):(4'hc)]))));
      reg303 <= ((~&reg301) ? reg290[(2'h2):(2'h2)] : reg269);
      reg304 <= $signed(({$signed($unsigned(wire298)),
          ($signed(wire299) ?
              wire259 : ((8'hb9) ?
                  reg273 : forvar267))} >> (^~$unsigned($signed(reg268)))));
      reg305 = $unsigned((~(reg266 ?
          $unsigned(wire252) : $unsigned((forvar263 ? wire259 : reg300)))));
    end
  assign wire306 = (reg290[(4'h9):(2'h2)] < $unsigned(reg294[(2'h2):(2'h2)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module202
#( parameter param244 = (((-((|(8'had)) ? (~^(8'ha6)) : ((8'hb7) - (8'hb0)))) ? {(^((8'h9e) | (8'ha8))), {(^(8'ha2))}} : (&(((8'hbc) ? (8'hac) : (8'hb6)) > ((8'ha5) ? (8'hac) : (8'had))))) | (~((((8'ha3) << (8'hb8)) ^ ((8'hae) ? (8'hb0) : (8'ha8))) <= (((8'hbc) << (8'hb0)) ^~ ((8'ha6) ? (8'hbe) : (7'h44))))))
, parameter param245 = param244 )
(y, clk, wire206, wire205, wire204, wire203);
  output wire [(32'h1ef):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire206;
  input wire [(4'he):(1'h0)] wire205;
  input wire [(5'h12):(1'h0)] wire204;
  input wire [(4'hd):(1'h0)] wire203;
  reg [(5'h14):(1'h0)] reg243 = (1'h0);
  reg [(3'h7):(1'h0)] reg242 = (1'h0);
  reg [(5'h15):(1'h0)] forvar238 = (1'h0);
  reg [(4'hd):(1'h0)] reg241 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg240 = (1'h0);
  reg [(5'h12):(1'h0)] reg239 = (1'h0);
  reg [(5'h14):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg237 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg236 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire235;
  reg [(4'hd):(1'h0)] reg234 = (1'h0);
  reg [(4'he):(1'h0)] reg233 = (1'h0);
  reg [(4'he):(1'h0)] reg232 = (1'h0);
  reg [(4'h9):(1'h0)] reg231 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg230 = (1'h0);
  wire [(3'h5):(1'h0)] wire229;
  wire [(4'ha):(1'h0)] wire228;
  reg signed [(4'hd):(1'h0)] reg227 = (1'h0);
  reg [(4'he):(1'h0)] reg226 = (1'h0);
  reg [(3'h4):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar224 = (1'h0);
  reg [(5'h11):(1'h0)] reg223 = (1'h0);
  reg [(5'h14):(1'h0)] reg222 = (1'h0);
  wire [(4'h9):(1'h0)] wire221;
  wire [(3'h4):(1'h0)] wire220;
  wire [(4'hb):(1'h0)] wire219;
  wire [(4'h8):(1'h0)] wire218;
  reg signed [(4'hb):(1'h0)] reg217 = (1'h0);
  reg [(4'he):(1'h0)] reg216 = (1'h0);
  reg [(5'h13):(1'h0)] reg215 = (1'h0);
  reg [(3'h6):(1'h0)] reg214 = (1'h0);
  reg [(5'h13):(1'h0)] reg213 = (1'h0);
  reg [(5'h14):(1'h0)] reg212 = (1'h0);
  reg [(3'h7):(1'h0)] forvar211 = (1'h0);
  reg [(4'ha):(1'h0)] reg211 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg209 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg207 = (1'h0);
  assign y = {reg243,
                 reg242,
                 forvar238,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 wire235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 wire229,
                 wire228,
                 reg227,
                 reg226,
                 reg225,
                 forvar224,
                 reg223,
                 reg222,
                 wire221,
                 wire220,
                 wire219,
                 wire218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 forvar211,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg207 <= ((^(!(!(wire204 ? wire204 : wire204)))) + (8'hb8));
      reg208 <= {wire205};
      if (wire204)
        begin
          reg209 = $unsigned(wire204[(1'h0):(1'h0)]);
          reg210 <= ({reg207[(5'h11):(4'ha)]} ?
              ($unsigned(wire204) << (^~$unsigned((wire205 ?
                  (7'h41) : reg208)))) : (~&wire204[(5'h10):(4'h9)]));
          reg211 <= {$unsigned(reg210)};
        end
      else
        begin
          reg209 <= (|{(((wire206 >>> reg211) ?
                  $signed(reg211) : (reg208 ?
                      wire204 : reg210)) & ($unsigned(wire206) || (reg207 ?
                  wire204 : (8'hae))))});
          reg210 = ((wire206 <<< $unsigned(reg207)) ?
              reg211[(1'h0):(1'h0)] : ($signed(reg211[(1'h1):(1'h0)]) ?
                  reg209 : wire203));
          for (forvar211 = (1'h0); (forvar211 < (2'h2)); forvar211 = (forvar211 + (1'h1)))
            begin
              reg212 <= $unsigned((wire203 ?
                  {(~&(!wire205))} : (^wire204[(1'h1):(1'h0)])));
              reg213 <= reg210[(3'h4):(2'h3)];
              reg214 <= (reg213[(5'h11):(1'h0)] ?
                  (+$signed((~&reg212))) : (-(~&(-$unsigned(wire204)))));
            end
          reg215 <= ((((&(reg208 & (8'h9c))) < wire206[(4'h8):(4'h8)]) & wire203[(2'h2):(2'h2)]) != (((&((8'hba) ^ reg213)) ~^ ($unsigned((7'h43)) ?
              $unsigned(reg213) : $unsigned(wire205))) < $unsigned((~&reg211))));
        end
      reg216 <= {wire205};
      reg217 <= (reg215[(4'he):(4'hb)] ? reg212 : reg214[(2'h3):(1'h0)]);
    end
  assign wire218 = reg216[(4'h8):(1'h1)];
  assign wire219 = $signed((~((~wire204) - wire204)));
  assign wire220 = reg208;
  assign wire221 = wire219[(4'h9):(2'h2)];
  always
    @(posedge clk) begin
      reg222 <= wire218;
      reg223 <= $signed(reg208[(1'h0):(1'h0)]);
      for (forvar224 = (1'h0); (forvar224 < (2'h3)); forvar224 = (forvar224 + (1'h1)))
        begin
          reg225 <= ((reg217[(4'ha):(3'h4)] != ($unsigned((reg211 ?
                  forvar211 : (8'hbe))) ?
              $signed((wire206 ?
                  forvar224 : reg223)) : (~$unsigned(reg207)))) > reg215[(2'h3):(2'h3)]);
          reg226 <= (reg210[(3'h5):(2'h2)] ^~ reg211[(4'h8):(3'h7)]);
          reg227 <= $unsigned(wire206[(4'h8):(2'h2)]);
        end
    end
  assign wire228 = $signed($signed((wire218 | reg227)));
  assign wire229 = wire203[(3'h6):(1'h1)];
  always
    @(posedge clk) begin
      reg230 = wire206;
      reg231 <= (~$signed({{{(8'hb1)}},
          ((reg210 & reg222) * ((8'ha4) != wire204))}));
      reg232 = (8'hac);
      reg233 <= {reg208[(1'h1):(1'h1)]};
      reg234 <= reg207;
    end
  assign wire235 = {wire206[(1'h1):(1'h0)]};
  always
    @(posedge clk) begin
      reg236 <= ((reg225 ~^ $signed($unsigned($signed(forvar211)))) ~^ (~(+(wire228[(3'h7):(3'h7)] ?
          $unsigned(wire228) : {(8'hb8), reg217}))));
      if ((((((8'ha6) == (reg234 ? reg234 : (8'h9f))) ?
          ((^~reg210) - (wire235 ? reg231 : reg215)) : ($unsigned(wire204) ?
              (reg215 ?
                  reg215 : (8'hbf)) : (|wire220))) <= ((reg223 >> {reg225}) ?
          $unsigned((~forvar224)) : reg214)) + $signed($signed({wire235}))))
        begin
          reg237 = (^(reg208[(1'h1):(1'h1)] ?
              $unsigned((|$signed(wire228))) : ((8'hbd) ?
                  $signed(reg216[(4'he):(4'h8)]) : ((reg222 * (8'ha4)) ?
                      {reg212, reg232} : reg222))));
          reg238 <= wire203[(4'hd):(4'h8)];
          reg239 <= reg232;
          reg240 <= $unsigned({$signed((+wire219)), reg207[(4'h8):(3'h5)]});
          reg241 <= ((($signed((reg237 >>> (8'h9c))) ?
              reg238 : ((&forvar211) ?
                  (reg232 ^~ reg217) : $signed(reg239))) ^~ reg231[(2'h2):(1'h1)]) ~^ (~&($unsigned((^reg207)) && {wire206,
              $unsigned(reg238)})));
        end
      else
        begin
          reg237 = (!reg212[(5'h13):(2'h3)]);
          for (forvar238 = (1'h0); (forvar238 < (1'h1)); forvar238 = (forvar238 + (1'h1)))
            begin
              reg239 = (+$unsigned($signed({(~|(8'hac)),
                  (reg238 ? (8'hb6) : reg213)})));
              reg240 <= (reg227[(4'hc):(4'hc)] ?
                  $unsigned((-((forvar224 ^ reg217) >= (~(8'hbc))))) : (~|(8'hb4)));
            end
          reg241 = wire206[(3'h4):(1'h1)];
        end
      reg242 = $unsigned((~$unsigned($signed($unsigned(forvar224)))));
      reg243 <= (&reg217[(3'h4):(1'h0)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module143  (y, clk, wire147, wire146, wire145, wire144);
  output wire [(32'h269):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire147;
  input wire [(5'h13):(1'h0)] wire146;
  input wire signed [(4'ha):(1'h0)] wire145;
  input wire signed [(5'h15):(1'h0)] wire144;
  reg [(5'h12):(1'h0)] reg199 = (1'h0);
  reg [(2'h3):(1'h0)] reg198 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire197;
  wire signed [(5'h12):(1'h0)] wire196;
  reg signed [(4'hd):(1'h0)] reg195 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg194 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg193 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg192 = (1'h0);
  wire signed [(4'he):(1'h0)] wire191;
  reg signed [(3'h5):(1'h0)] reg190 = (1'h0);
  reg [(2'h2):(1'h0)] reg189 = (1'h0);
  reg [(2'h2):(1'h0)] reg188 = (1'h0);
  reg [(3'h5):(1'h0)] reg187 = (1'h0);
  reg [(3'h5):(1'h0)] reg186 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire185;
  wire signed [(5'h12):(1'h0)] wire184;
  wire signed [(5'h11):(1'h0)] wire183;
  reg [(5'h14):(1'h0)] reg182 = (1'h0);
  reg [(4'ha):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg180 = (1'h0);
  reg [(4'h8):(1'h0)] reg179 = (1'h0);
  reg [(4'ha):(1'h0)] reg178 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg177 = (1'h0);
  reg [(3'h6):(1'h0)] forvar176 = (1'h0);
  reg [(5'h14):(1'h0)] reg175 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg173 = (1'h0);
  reg [(4'he):(1'h0)] reg172 = (1'h0);
  reg [(3'h6):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg170 = (1'h0);
  reg [(5'h13):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar168 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg167 = (1'h0);
  reg [(3'h6):(1'h0)] reg166 = (1'h0);
  reg signed [(4'he):(1'h0)] reg165 = (1'h0);
  wire [(5'h12):(1'h0)] wire164;
  wire signed [(4'hc):(1'h0)] wire163;
  reg signed [(5'h15):(1'h0)] reg162 = (1'h0);
  reg [(4'h8):(1'h0)] reg161 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg160 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg159 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg158 = (1'h0);
  reg [(4'hc):(1'h0)] reg157 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg156 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg155 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg154 = (1'h0);
  reg [(4'hb):(1'h0)] reg153 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg152 = (1'h0);
  reg [(2'h2):(1'h0)] forvar151 = (1'h0);
  wire [(4'ha):(1'h0)] wire150;
  wire [(4'h9):(1'h0)] wire149;
  reg [(5'h13):(1'h0)] reg148 = (1'h0);
  assign y = {reg199,
                 reg198,
                 wire197,
                 wire196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 wire191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 wire185,
                 wire184,
                 wire183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 forvar176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 forvar168,
                 reg167,
                 reg166,
                 reg165,
                 wire164,
                 wire163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 forvar151,
                 wire150,
                 wire149,
                 reg148,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg148 <= (~&$signed((8'h9e)));
    end
  assign wire149 = wire144[(4'h8):(3'h7)];
  assign wire150 = $signed((!wire149));
  always
    @(posedge clk) begin
      for (forvar151 = (1'h0); (forvar151 < (3'h4)); forvar151 = (forvar151 + (1'h1)))
        begin
          reg152 <= wire150;
          reg153 = (~$unsigned(wire149));
        end
    end
  always
    @(posedge clk) begin
      reg154 = {{($signed($signed((8'hab))) * $signed((wire144 ?
                  wire145 : forvar151)))},
          (8'ha9)};
      reg155 = ((wire144 + wire146[(3'h7):(2'h3)]) ?
          wire144[(5'h11):(5'h11)] : $unsigned($signed($signed((~wire149)))));
      reg156 <= reg148[(4'h9):(3'h6)];
      reg157 = $signed({$signed({{reg153, (8'h9e)}, wire150[(4'ha):(3'h4)]}),
          {wire147, (~^wire147)}});
      reg158 <= (wire149[(2'h2):(2'h2)] || $unsigned($unsigned($unsigned(reg152))));
    end
  always
    @(posedge clk) begin
      reg159 <= {$unsigned(($unsigned((reg155 & reg153)) * reg153[(4'ha):(2'h3)]))};
      reg160 = ((($signed($unsigned(wire144)) ?
              $signed((wire146 <<< (8'hac))) : (~&$unsigned(wire149))) << (~^wire146)) ?
          reg153[(4'ha):(4'ha)] : wire144[(4'hc):(4'ha)]);
      reg161 <= $signed((((~&$signed(wire147)) ^~ (wire147 ?
              ((7'h40) ^ reg157) : $signed(wire149))) ?
          {(forvar151[(1'h0):(1'h0)] ?
                  (reg155 ?
                      reg153 : (8'haf)) : wire146)} : {wire150[(3'h6):(2'h2)]}));
      reg162 = reg160[(4'hb):(3'h5)];
    end
  assign wire163 = $signed((({$unsigned(forvar151), reg158[(2'h3):(1'h1)]} ?
                           (wire150[(4'h8):(1'h0)] >>> (8'hbb)) : reg154[(2'h2):(1'h1)]) ?
                       $signed(((reg148 ? wire147 : reg155) ?
                           reg162[(4'h9):(1'h0)] : (reg161 ?
                               (8'hbc) : reg156))) : $unsigned(reg162[(1'h1):(1'h1)])));
  assign wire164 = (~|$unsigned((+$signed($unsigned(wire145)))));
  always
    @(posedge clk) begin
      reg165 <= $unsigned(((reg156 ?
              (reg161 ?
                  (reg152 >> reg155) : (wire163 * reg162)) : ({(8'hb7)} << {(8'hb6)})) ?
          $signed((^~wire150[(1'h0):(1'h0)])) : reg160[(2'h2):(1'h1)]));
      reg166 <= $signed((7'h42));
      reg167 = {(^{((wire164 + reg152) ^~ ((8'ha9) + (8'hae)))})};
      for (forvar168 = (1'h0); (forvar168 < (1'h0)); forvar168 = (forvar168 + (1'h1)))
        begin
          reg169 <= $unsigned((reg162 << ($unsigned($unsigned(wire146)) ?
              reg148[(4'h9):(3'h6)] : (reg159[(2'h3):(1'h1)] & wire145[(3'h7):(3'h6)]))));
          reg170 <= ((($signed(reg165) ?
              ((wire164 ? (8'hba) : wire145) >>> {wire164,
                  forvar151}) : $unsigned(reg166)) & reg155[(1'h0):(1'h0)]) <<< (wire150[(1'h1):(1'h1)] ?
              reg155[(1'h1):(1'h0)] : $signed((~&$unsigned(reg154)))));
          reg171 <= reg148;
          reg172 <= $unsigned(reg170);
        end
      if ((+reg155))
        begin
          reg173 = wire150;
          reg174 <= reg172;
        end
      else
        begin
          if ((~|(~&forvar151[(2'h2):(2'h2)])))
            begin
              reg173 <= $signed($unsigned(((((8'ha1) ? reg160 : (8'ha2)) ?
                      {wire164, wire164} : {reg160, (8'h9f)}) ?
                  wire164[(3'h7):(2'h3)] : $signed(((8'ha3) ?
                      reg167 : forvar168)))));
              reg174 <= (reg156[(1'h0):(1'h0)] <= reg160);
              reg175 <= reg162[(3'h4):(2'h2)];
            end
          else
            begin
              reg173 <= (!$unsigned($unsigned($unsigned(forvar151))));
              reg174 <= wire163[(4'h9):(3'h6)];
            end
          for (forvar176 = (1'h0); (forvar176 < (3'h4)); forvar176 = (forvar176 + (1'h1)))
            begin
              reg177 <= (8'hbb);
              reg178 <= $unsigned(wire147);
              reg179 <= $signed($signed(($signed((^~reg156)) ^ reg153)));
              reg180 <= reg169[(3'h4):(2'h2)];
              reg181 <= (reg152[(2'h3):(2'h2)] > $unsigned($unsigned(($signed(reg177) & (+reg162)))));
            end
          reg182 <= (((-{reg178,
              reg166[(3'h5):(1'h1)]}) * reg174) - $signed(($signed(wire164) - reg162)));
        end
    end
  assign wire183 = ((&reg171) ?
                       $signed((reg155 ?
                           ($signed(reg161) ?
                               (reg161 ? (8'h9d) : reg177) : {reg159,
                                   (8'hb4)}) : ((reg182 ? reg177 : wire144) ?
                               reg157 : (reg171 <= reg159)))) : ((reg158 ?
                           (+(wire147 ? reg173 : wire164)) : ((reg180 ?
                               forvar151 : (7'h44)) | reg177)) ^~ (~|(~&(wire150 < reg177)))));
  assign wire184 = reg160;
  assign wire185 = {(|reg162[(3'h6):(3'h5)])};
  always
    @(posedge clk) begin
      reg186 <= $unsigned(wire183[(3'h6):(1'h1)]);
      reg187 <= reg174;
      reg188 = wire149[(3'h7):(3'h7)];
      reg189 = ($unsigned($unsigned(reg173)) <<< ($unsigned(((wire185 <= reg171) ?
          (reg188 - reg167) : $unsigned((8'ha8)))) != (8'ha6)));
      reg190 <= reg160;
    end
  assign wire191 = $signed((8'hb8));
  always
    @(posedge clk) begin
      reg192 = ((+$unsigned(reg167)) <= (^({(-reg175),
          $signed((8'haa))} & $signed($unsigned(reg172)))));
      reg193 <= $signed(reg188[(2'h2):(1'h0)]);
      reg194 = {reg173[(3'h6):(1'h0)],
          {$unsigned($unsigned((reg173 >= wire147))),
              $signed($signed(reg159))}};
      reg195 = (^((reg172[(4'hb):(1'h0)] <<< $unsigned((reg188 & reg162))) ^~ $signed(reg179[(1'h1):(1'h0)])));
    end
  assign wire196 = $unsigned(($unsigned({(|wire149)}) ?
                       ({((8'ha3) & reg154)} ?
                           ($unsigned(reg180) ?
                               (wire183 ?
                                   reg173 : wire163) : (^reg193)) : reg178[(3'h4):(1'h1)]) : reg193));
  assign wire197 = $unsigned(wire144);
  always
    @(posedge clk) begin
      reg198 <= $signed(wire145[(4'ha):(1'h0)]);
      reg199 <= reg193[(5'h10):(3'h7)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module394
#( parameter param447 = ((^({((8'ha8) ? (8'h9c) : (7'h40))} > ((8'hbe) < ((8'hbf) <<< (8'h9c))))) ? (~|{(8'hb4)}) : (&(~&(((8'h9f) ? (8'h9c) : (8'ha9)) ? (~(8'ha2)) : ((8'hb7) - (8'hae))))))
, parameter param448 = ((8'h9c) == ({param447, ((param447 ? (8'ha8) : param447) ? param447 : ((8'ha4) >= param447))} ? {(8'had)} : (((param447 ? (8'hbc) : param447) >= param447) ? ({param447, param447} ? (~^param447) : (&param447)) : (~&((8'hb3) ? param447 : param447))))) )
(y, clk, wire398, wire397, wire396, wire395);
  output wire [(32'h209):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire398;
  input wire signed [(5'h10):(1'h0)] wire397;
  input wire [(4'hf):(1'h0)] wire396;
  input wire signed [(2'h2):(1'h0)] wire395;
  wire signed [(4'hc):(1'h0)] wire446;
  wire signed [(4'h9):(1'h0)] wire445;
  reg signed [(4'he):(1'h0)] reg444 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg443 = (1'h0);
  reg [(5'h10):(1'h0)] reg442 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg428 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg440 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar439 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg438 = (1'h0);
  reg [(3'h7):(1'h0)] reg437 = (1'h0);
  reg [(3'h7):(1'h0)] reg436 = (1'h0);
  reg [(4'hc):(1'h0)] reg435 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg434 = (1'h0);
  reg [(3'h6):(1'h0)] reg433 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar432 = (1'h0);
  reg [(2'h3):(1'h0)] reg431 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg430 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg429 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar428 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg427 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire426;
  wire [(4'hb):(1'h0)] wire425;
  wire signed [(3'h4):(1'h0)] wire424;
  reg signed [(5'h12):(1'h0)] reg423 = (1'h0);
  reg [(2'h3):(1'h0)] reg422 = (1'h0);
  reg [(3'h6):(1'h0)] forvar421 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg420 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg419 = (1'h0);
  reg [(5'h13):(1'h0)] reg418 = (1'h0);
  wire [(4'ha):(1'h0)] wire417;
  reg signed [(2'h2):(1'h0)] reg416 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg415 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg413 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg412 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg411 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire410;
  reg [(4'ha):(1'h0)] reg409 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg408 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg407 = (1'h0);
  reg [(4'hc):(1'h0)] reg406 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire405;
  reg [(5'h14):(1'h0)] reg404 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg403 = (1'h0);
  reg [(3'h4):(1'h0)] reg402 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar401 = (1'h0);
  reg [(3'h7):(1'h0)] reg400 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire399;
  assign y = {wire446,
                 wire445,
                 reg444,
                 reg443,
                 reg442,
                 reg428,
                 reg441,
                 reg440,
                 forvar439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 forvar432,
                 reg431,
                 reg430,
                 reg429,
                 forvar428,
                 reg427,
                 wire426,
                 wire425,
                 wire424,
                 reg423,
                 reg422,
                 forvar421,
                 reg420,
                 reg419,
                 reg418,
                 wire417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 wire410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 wire405,
                 reg404,
                 reg403,
                 reg402,
                 forvar401,
                 reg400,
                 wire399,
                 (1'h0)};
  assign wire399 = (^~$signed((wire395[(1'h1):(1'h0)] ?
                       $unsigned((wire398 ? wire395 : wire396)) : wire395)));
  always
    @(posedge clk) begin
      reg400 <= ((7'h40) ?
          (~&(wire399 || (-(&wire397)))) : (wire397 | ($signed(wire396[(3'h5):(3'h4)]) < ($signed(wire397) ?
              (~|wire396) : (wire395 & (8'ha2))))));
      for (forvar401 = (1'h0); (forvar401 < (2'h3)); forvar401 = (forvar401 + (1'h1)))
        begin
          reg402 <= {wire398,
              ($signed(wire395[(1'h1):(1'h0)]) && ($signed({forvar401}) >> (~^$unsigned((8'ha9)))))};
          reg403 <= (({$unsigned((~|(8'hab))),
                  $unsigned((wire396 ?
                      wire396 : wire398))} > $signed($signed({(8'ha9)}))) ?
              ((reg402[(2'h3):(2'h2)] ?
                      ((wire397 ?
                          wire398 : (8'hb8)) < $signed(wire399)) : ($signed((8'h9c)) << (^wire395))) ?
                  wire396[(4'h9):(2'h2)] : $unsigned(((reg400 ?
                          wire398 : wire398) ?
                      (^wire396) : ((8'hb1) < reg402)))) : reg402);
        end
      reg404 <= $unsigned(wire395);
    end
  assign wire405 = ((reg402 >= wire398[(3'h7):(1'h0)]) ?
                       ($signed(({wire398} ~^ (^~wire398))) && {(wire397[(1'h0):(1'h0)] ?
                               reg402[(1'h0):(1'h0)] : (wire396 ?
                                   wire398 : wire399)),
                           (8'ha1)}) : {{wire398[(3'h4):(2'h3)],
                               wire397[(4'h9):(4'h8)]},
                           (-$signed($signed((8'hb7))))});
  always
    @(posedge clk) begin
      reg406 = (($unsigned(wire398[(4'h8):(1'h1)]) && $unsigned(((8'hb0) ^~ (reg403 ?
              wire399 : reg400)))) ?
          ((wire405 >> (reg403 ?
              wire398[(3'h5):(3'h5)] : (wire398 ?
                  reg402 : wire397))) * ($unsigned(((8'had) ?
                  reg404 : forvar401)) ?
              ((8'ha9) <<< $signed(wire405)) : forvar401)) : $signed((7'h41)));
      reg407 <= (|(wire397[(3'h7):(1'h1)] ^ {($signed(wire397) ?
              wire399 : (reg402 ? wire395 : (8'hb9)))}));
      reg408 <= $signed((($signed(forvar401[(2'h2):(2'h2)]) <= wire397) ?
          $unsigned((+(wire405 >>> wire397))) : $signed($signed((wire405 ?
              wire399 : forvar401)))));
      reg409 <= wire397[(2'h2):(2'h2)];
    end
  assign wire410 = $unsigned(((wire396[(4'ha):(3'h7)] * ((~|reg402) << wire396)) ?
                       reg400 : $unsigned((reg400[(3'h4):(1'h0)] >> {(8'hb8),
                           reg407}))));
  always
    @(posedge clk) begin
      reg411 = {(+($signed((reg406 > wire410)) ?
              $unsigned($signed(wire396)) : ($signed(reg400) ?
                  ((8'ha4) << wire399) : (wire397 >= reg408))))};
      reg412 = $unsigned(((8'h9e) ?
          ($unsigned(wire399) >>> reg406) : $signed(reg400[(3'h6):(3'h4)])));
      reg413 <= (-(($unsigned(wire397) ? reg408 : (wire396 >>> (~forvar401))) ?
          wire397 : ($signed((&wire399)) == (wire398 ?
              $signed(reg403) : {reg406}))));
      reg414 = (reg400[(2'h2):(2'h2)] ?
          (~$unsigned($unsigned($unsigned(reg404)))) : (wire399 ?
              wire395[(2'h2):(1'h1)] : $signed($unsigned({reg400}))));
    end
  always
    @(posedge clk) begin
      reg415 = ((~|(~&(~|(reg414 ?
          wire410 : (8'ha8))))) * ($unsigned((~(~^reg409))) || $signed((!reg409[(3'h7):(2'h2)]))));
    end
  always
    @(posedge clk) begin
      reg416 <= (((((forvar401 ? reg409 : forvar401) ^ ((8'hab) ?
              reg402 : reg415)) < wire405[(1'h1):(1'h1)]) ?
          ((~^(~&reg411)) || reg404[(4'h9):(3'h4)]) : $unsigned((wire396 ~^ $unsigned(wire398)))) >> forvar401);
    end
  assign wire417 = (reg409[(4'ha):(3'h7)] ^ $unsigned($signed($signed(reg414[(4'hd):(3'h4)]))));
  always
    @(posedge clk) begin
      reg418 <= $signed((((+(reg400 && wire410)) ?
          {(^~reg402)} : ((reg402 >> reg409) > (!wire417))) >= reg403));
      reg419 <= $signed((-($signed((wire398 ?
          forvar401 : reg402)) || reg402[(2'h3):(1'h0)])));
      reg420 <= (reg402[(2'h3):(1'h1)] ~^ (8'hbc));
    end
  always
    @(posedge clk) begin
      for (forvar421 = (1'h0); (forvar421 < (2'h2)); forvar421 = (forvar421 + (1'h1)))
        begin
          reg422 = reg408;
        end
      reg423 <= $signed((-$unsigned((~|$signed(reg420)))));
    end
  assign wire424 = (~reg407);
  assign wire425 = $unsigned($unsigned(($unsigned({reg422, reg408}) ?
                       $signed((!reg412)) : (~|((8'ha1) <<< wire395)))));
  assign wire426 = $unsigned((^reg414));
  always
    @(posedge clk) begin
      reg427 <= (&(reg415[(1'h1):(1'h1)] ?
          (($unsigned(wire405) ~^ (reg409 ? forvar401 : reg411)) ?
              ($signed(forvar401) & {reg404, (8'ha9)}) : $signed(((8'hba) ?
                  reg411 : (7'h44)))) : reg418[(4'hd):(4'ha)]));
      if ($signed($unsigned(wire410)))
        begin
          for (forvar428 = (1'h0); (forvar428 < (2'h3)); forvar428 = (forvar428 + (1'h1)))
            begin
              reg429 <= wire425;
              reg430 <= ($signed((~((-reg423) | reg423[(4'h9):(2'h3)]))) ?
                  forvar428[(2'h2):(1'h0)] : {($unsigned({(8'hbc),
                          (8'hb1)}) & (wire426[(4'hc):(3'h7)] - (~|reg423))),
                      {wire395, (!$signed(reg412))}});
              reg431 <= {$unsigned(wire410[(4'hf):(4'ha)]),
                  (wire397[(4'he):(3'h4)] >> (8'haf))};
            end
          for (forvar432 = (1'h0); (forvar432 < (2'h3)); forvar432 = (forvar432 + (1'h1)))
            begin
              reg433 <= reg431;
              reg434 = $unsigned((reg431 ?
                  (reg403 ?
                      reg420 : ($unsigned((8'hb2)) || forvar428[(3'h4):(1'h0)])) : wire417));
              reg435 = $signed((reg413[(4'hf):(2'h3)] ?
                  (^(~&((8'haa) ?
                      wire405 : forvar421))) : (((7'h40) <= {reg408}) ?
                      $unsigned($unsigned(reg431)) : (|(reg422 ?
                          forvar421 : (8'hbc))))));
              reg436 <= reg400[(2'h3):(2'h3)];
              reg437 = $unsigned(reg419[(4'he):(3'h7)]);
            end
          reg438 <= reg416[(1'h1):(1'h1)];
          for (forvar439 = (1'h0); (forvar439 < (2'h3)); forvar439 = (forvar439 + (1'h1)))
            begin
              reg440 <= $unsigned(({reg427} ?
                  $signed($signed(reg407[(1'h1):(1'h1)])) : $signed($signed((reg408 ?
                      wire425 : (8'hb5))))));
              reg441 <= reg430;
            end
        end
      else
        begin
          reg428 <= {(~&$unsigned(($unsigned((8'h9c)) < reg438[(1'h1):(1'h0)]))),
              {((wire405[(2'h3):(1'h1)] ?
                          ((7'h41) ? reg422 : reg400) : (reg406 ?
                              (7'h40) : reg402)) ?
                      (reg416[(1'h0):(1'h0)] ?
                          wire417[(4'h9):(3'h5)] : $unsigned(forvar421)) : {reg434[(1'h1):(1'h1)]}),
                  (($unsigned(reg441) <= (reg407 ? wire424 : wire399)) ?
                      reg400[(2'h2):(1'h0)] : $unsigned((forvar428 - (8'hb4))))}};
        end
      reg442 = ((&$unsigned((~&$signed(reg419)))) ?
          ((^~(^~(+reg409))) ?
              $unsigned((+wire397)) : $signed(reg441)) : wire426[(3'h7):(3'h6)]);
      reg443 = {reg431[(2'h3):(1'h0)], {{wire424[(2'h2):(1'h0)]}}};
      reg444 <= reg411[(3'h5):(2'h3)];
    end
  assign wire445 = $unsigned(((+reg402) ?
                       (($unsigned((8'hac)) >>> $unsigned(wire426)) ?
                           (reg443 ?
                               $signed(reg400) : (~reg423)) : forvar401[(2'h2):(1'h0)]) : (reg413[(4'h9):(4'h8)] ^ {wire405[(1'h1):(1'h0)]})));
  assign wire446 = (-(8'hb4));
endmodule