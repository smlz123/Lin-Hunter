(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h8c9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire0;
  input wire [(3'h7):(1'h0)] wire1;
  input wire signed [(4'hb):(1'h0)] wire2;
  input wire [(5'h10):(1'h0)] wire3;
  reg [(4'hc):(1'h0)] reg3327 = (1'h0);
  reg [(4'he):(1'h0)] reg3326 = (1'h0);
  reg [(4'h8):(1'h0)] reg3325 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3324 = (1'h0);
  reg [(4'hb):(1'h0)] reg3323 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3322 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3321 = (1'h0);
  reg [(4'hb):(1'h0)] reg3320 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3319 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3318 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3317 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3316 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar3315 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3314 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3313 = (1'h0);
  reg [(5'h16):(1'h0)] reg3312 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3311 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar3310 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3309 = (1'h0);
  reg [(4'h9):(1'h0)] reg3308 = (1'h0);
  reg [(4'he):(1'h0)] reg3307 = (1'h0);
  reg [(5'h13):(1'h0)] reg3306 = (1'h0);
  reg [(5'h15):(1'h0)] reg3305 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3304 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3303 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3302 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3301 = (1'h0);
  reg [(3'h6):(1'h0)] reg3300 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3299 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3298 = (1'h0);
  reg [(5'h13):(1'h0)] reg3297 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3296 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3295 = (1'h0);
  wire signed [(5'h19):(1'h0)] wire3294;
  reg [(4'ha):(1'h0)] reg3293 = (1'h0);
  reg [(3'h5):(1'h0)] reg3292 = (1'h0);
  reg [(5'h11):(1'h0)] forvar3291 = (1'h0);
  reg [(3'h6):(1'h0)] reg3290 = (1'h0);
  reg [(4'he):(1'h0)] reg3289 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3279 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3278 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3288 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3287 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3286 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3285 = (1'h0);
  reg [(5'h15):(1'h0)] reg3284 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3283 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3282 = (1'h0);
  reg [(3'h6):(1'h0)] reg3281 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3280 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3279 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3278 = (1'h0);
  reg [(5'h11):(1'h0)] reg3277 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3276 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3275 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire3221;
  wire signed [(4'hf):(1'h0)] wire3219;
  wire [(5'h15):(1'h0)] wire3217;
  wire [(5'h18):(1'h0)] wire3216;
  reg [(4'hf):(1'h0)] reg3215 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3214 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3213 = (1'h0);
  wire [(5'h15):(1'h0)] wire3212;
  reg [(5'h19):(1'h0)] forvar4 = (1'h0);
  reg [(5'h1a):(1'h0)] reg5 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg6 = (1'h0);
  reg [(5'h16):(1'h0)] reg7 = (1'h0);
  reg [(5'h19):(1'h0)] forvar8 = (1'h0);
  reg [(5'h12):(1'h0)] reg9 = (1'h0);
  reg [(5'h14):(1'h0)] reg10 = (1'h0);
  reg [(5'h1a):(1'h0)] reg11 = (1'h0);
  reg [(4'hb):(1'h0)] reg12 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg13 = (1'h0);
  reg [(4'hb):(1'h0)] reg14 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg15 = (1'h0);
  reg [(5'h13):(1'h0)] reg16 = (1'h0);
  reg [(4'ha):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar13 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar17 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg20 = (1'h0);
  reg [(4'he):(1'h0)] reg21 = (1'h0);
  reg [(5'h18):(1'h0)] reg22 = (1'h0);
  reg [(5'h1a):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar24 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg28 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg29 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar30 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg31 = (1'h0);
  reg [(5'h19):(1'h0)] reg32 = (1'h0);
  reg [(5'h11):(1'h0)] reg33 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire3210;
  wire [(5'h19):(1'h0)] wire3223;
  wire signed [(5'h18):(1'h0)] wire3225;
  wire [(5'h11):(1'h0)] wire3227;
  wire [(5'h19):(1'h0)] wire3229;
  reg signed [(5'h16):(1'h0)] forvar3230 = (1'h0);
  reg [(5'h19):(1'h0)] reg3231 = (1'h0);
  reg [(2'h2):(1'h0)] reg3232 = (1'h0);
  reg [(5'h10):(1'h0)] reg3233 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3234 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3235 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3236 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3237 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3238 = (1'h0);
  reg [(4'hc):(1'h0)] reg3239 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3240 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3241 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3242 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3243 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3244 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3245 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3246 = (1'h0);
  reg [(2'h3):(1'h0)] reg3247 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3248 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg3249 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3242 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3250 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3251 = (1'h0);
  wire [(2'h3):(1'h0)] wire3252;
  wire signed [(5'h18):(1'h0)] wire3254;
  reg signed [(5'h14):(1'h0)] forvar3255 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3256 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3257 = (1'h0);
  reg [(5'h11):(1'h0)] reg3258 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3259 = (1'h0);
  reg [(5'h12):(1'h0)] reg3260 = (1'h0);
  reg [(2'h3):(1'h0)] reg3261 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3262 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3263 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3264 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3265 = (1'h0);
  reg [(5'h12):(1'h0)] reg3266 = (1'h0);
  reg [(3'h5):(1'h0)] reg3267 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3268 = (1'h0);
  reg [(5'h10):(1'h0)] reg3269 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire3270;
  wire signed [(5'h10):(1'h0)] wire3271;
  wire [(4'ha):(1'h0)] wire3272;
  wire [(4'h9):(1'h0)] wire3273;
  assign y = {reg3327,
                 reg3326,
                 reg3325,
                 reg3324,
                 reg3323,
                 reg3322,
                 reg3321,
                 reg3320,
                 reg3319,
                 reg3318,
                 reg3317,
                 reg3316,
                 forvar3315,
                 reg3314,
                 reg3313,
                 reg3312,
                 reg3311,
                 forvar3310,
                 forvar3309,
                 reg3308,
                 reg3307,
                 reg3306,
                 reg3305,
                 reg3304,
                 reg3303,
                 forvar3302,
                 forvar3301,
                 reg3300,
                 reg3299,
                 reg3298,
                 reg3297,
                 forvar3296,
                 forvar3295,
                 wire3294,
                 reg3293,
                 reg3292,
                 forvar3291,
                 reg3290,
                 reg3289,
                 reg3279,
                 forvar3278,
                 reg3288,
                 reg3287,
                 reg3286,
                 reg3285,
                 reg3284,
                 reg3283,
                 reg3282,
                 reg3281,
                 reg3280,
                 forvar3279,
                 reg3278,
                 reg3277,
                 forvar3276,
                 reg3275,
                 wire3221,
                 wire3219,
                 wire3217,
                 wire3216,
                 reg3215,
                 reg3214,
                 reg3213,
                 wire3212,
                 forvar4,
                 reg5,
                 reg6,
                 reg7,
                 forvar8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 forvar13,
                 forvar17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 forvar24,
                 reg25,
                 reg26,
                 reg27,
                 reg28,
                 reg29,
                 forvar30,
                 reg31,
                 reg32,
                 reg33,
                 wire3210,
                 wire3223,
                 wire3225,
                 wire3227,
                 wire3229,
                 forvar3230,
                 reg3231,
                 reg3232,
                 reg3233,
                 reg3234,
                 forvar3235,
                 reg3236,
                 reg3237,
                 reg3238,
                 reg3239,
                 reg3240,
                 reg3241,
                 forvar3242,
                 reg3243,
                 reg3244,
                 reg3245,
                 reg3246,
                 reg3247,
                 reg3248,
                 reg3249,
                 reg3242,
                 reg3250,
                 reg3251,
                 wire3252,
                 wire3254,
                 forvar3255,
                 reg3256,
                 forvar3257,
                 reg3258,
                 reg3259,
                 reg3260,
                 reg3261,
                 reg3262,
                 reg3263,
                 reg3264,
                 reg3265,
                 reg3266,
                 reg3267,
                 reg3268,
                 reg3269,
                 wire3270,
                 wire3271,
                 wire3272,
                 wire3273,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar4 = (1'h0); (forvar4 < (2'h2)); forvar4 = (forvar4 + (1'h1)))
        begin
          reg5 <= wire3[(1'h1):(1'h1)];
          reg6 <= wire2;
          reg7 <= $unsigned((forvar4[(3'h4):(1'h1)] ?
              ({(wire3 <= wire1)} ?
                  "vJS4Ztf01IkX32sW" : {(wire1 | (7'h47))}) : wire3));
          for (forvar8 = (1'h0); (forvar8 < (2'h3)); forvar8 = (forvar8 + (1'h1)))
            begin
              reg9 <= ($signed(wire3[(2'h2):(2'h2)]) ?
                  {$signed(({forvar4, (8'hbc)} ?
                          (~^(7'h4c)) : "wsQspv85A9xahZhXrAm7"))} : $signed({wire2,
                      $unsigned($unsigned(wire1))}));
              reg10 <= wire2;
              reg11 <= wire0;
            end
          if (($unsigned("7pJ0XbdIFe1K8") ?
              $signed(wire1[(3'h6):(2'h2)]) : "NMgYgaFVcqSwlIpRgVN"))
            begin
              reg12 <= (+"LP");
              reg13 = "vwxH3WbkNluLG9rEm9ZwSBIv";
              reg14 <= $signed($signed(wire0[(3'h6):(1'h0)]));
              reg15 <= ((|reg14[(3'h4):(2'h2)]) ?
                  ((8'hb6) ?
                      reg10 : ($unsigned((reg12 * reg7)) | $unsigned((reg14 ?
                          reg14 : wire0)))) : (~"3LUVzPdTs"));
              reg16 <= wire1[(2'h3):(2'h3)];
              reg17 = (+("dmsNCgg" ?
                  forvar4 : ((reg13[(1'h0):(1'h0)] - "ofpktKtyteBE5a7c9oZWZKCK") ?
                      "FWVLidpJkWnOfymdd" : $signed(reg13))));
            end
          else
            begin
              reg12 <= forvar8[(3'h7):(3'h7)];
              for (forvar13 = (1'h0); (forvar13 < (3'h4)); forvar13 = (forvar13 + (1'h1)))
                begin
                  reg14 <= $signed($unsigned((8'hab)));
                  reg15 <= $unsigned((~&((8'hb0) * ($signed(reg14) ?
                      {(8'ha0)} : $signed(reg5)))));
                end
              reg16 <= wire2[(3'h6):(3'h5)];
              for (forvar17 = (1'h0); (forvar17 < (3'h5)); forvar17 = (forvar17 + (1'h1)))
                begin
                  reg18 <= (8'hbf);
                  reg19 = $signed((^(("e" != ((8'ha6) ?
                      (8'had) : reg9)) + wire2)));
                  reg20 <= wire1;
                  reg21 <= $signed(forvar17[(2'h2):(2'h2)]);
                  reg22 <= ($signed($unsigned($signed($signed(forvar4)))) & $signed((^reg12)));
                  reg23 = reg14;
                end
              for (forvar24 = (1'h0); (forvar24 < (1'h1)); forvar24 = (forvar24 + (1'h1)))
                begin
                  reg25 <= ("Mh4s" ^ $signed(forvar13));
                  reg26 = reg25[(1'h0):(1'h0)];
                  reg27 <= reg23[(4'h9):(3'h7)];
                end
              reg28 <= "gZhTc3WyGJQqBJIHZwrb6JYl";
            end
        end
      reg29 <= $signed("8ZxonOPMtuA");
      for (forvar30 = (1'h0); (forvar30 < (1'h1)); forvar30 = (forvar30 + (1'h1)))
        begin
          reg31 <= (!reg29[(1'h0):(1'h0)]);
          reg32 <= (forvar13 ^~ "i1oKOi6euiuEJW9q");
          reg33 <= $signed($unsigned(wire2));
        end
    end
  module34 modinst3211 (wire3210, clk, reg25, wire3, reg28, reg11, forvar4);
  assign wire3212 = wire2[(4'h8):(3'h4)];
  always
    @(posedge clk) begin
      reg3213 <= ($unsigned(($unsigned((reg14 <= reg5)) <= reg13[(3'h4):(2'h2)])) >= "WP");
      reg3214 = $unsigned((~"5P9G21GQD8I5VpAZlwkSRv"));
      reg3215 <= ("cEZ2wrEunU" ?
          {($unsigned("8I") ?
                  $signed("bToY4FCMP9NcrJy4") : $signed(wire3[(5'h10):(4'h8)]))} : $unsigned(wire3212[(3'h5):(2'h3)]));
    end
  assign wire3216 = ($unsigned("c") ?
                        ({$unsigned((forvar24 ?
                                reg26 : wire0))} || (((|forvar4) || {reg28}) ?
                            {reg32} : wire3210[(1'h1):(1'h1)])) : forvar17);
  module48 modinst3218 (wire3217, clk, reg28, reg23, reg19, forvar30);
  module1753 modinst3220 (wire3219, clk, reg18, forvar4, reg23, reg31);
  module1953 modinst3222 (.y(wire3221), .wire1955(wire3217), .wire1958(reg28), .clk(clk), .wire1957(reg31), .wire1956(reg7), .wire1954(reg3213));
  module2298 modinst3224 (wire3223, clk, reg3215, reg9, reg6, reg19);
  module1753 modinst3226 (wire3225, clk, wire3216, reg32, reg3213, reg3215);
  module2349 modinst3228 (.wire2351(reg32), .y(wire3227), .wire2350(reg31), .wire2352(forvar8), .clk(clk), .wire2353(reg6));
  assign wire3229 = ({({(reg32 < wire3221)} ~^ "s"),
                            ($signed(reg23) >= wire3223)} ?
                        "pHDtl1" : reg20);
  always
    @(posedge clk) begin
      for (forvar3230 = (1'h0); (forvar3230 < (3'h4)); forvar3230 = (forvar3230 + (1'h1)))
        begin
          reg3231 = $signed((wire0[(4'h8):(3'h5)] ~^ wire3221));
        end
      reg3232 <= wire3225[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg3233 <= ("3XvBlJdSyvoN5TcPrDYv0" ?
          ({$signed((forvar3230 ? (7'h49) : wire3221)),
              (reg32 ?
                  $unsigned(reg6) : "A")} == (!wire0[(2'h2):(1'h1)])) : (reg29[(1'h0):(1'h0)] ?
              reg3231 : "zdV3t0wpcAxUi"));
      reg3234 <= "gvhalIu0";
      for (forvar3235 = (1'h0); (forvar3235 < (3'h4)); forvar3235 = (forvar3235 + (1'h1)))
        begin
          reg3236 <= $unsigned((~^{wire3212, (~^"4ITrxdgkCC3qCqx390npg")}));
          reg3237 <= "zOmMRRtU8DV9fc";
          reg3238 <= reg5;
        end
    end
  always
    @(posedge clk) begin
      reg3239 <= (forvar30[(3'h4):(1'h0)] ? reg9[(5'h10):(3'h6)] : (+wire3229));
      reg3240 = $unsigned(forvar17[(4'ha):(4'h9)]);
      reg3241 <= reg3214;
      if (reg27)
        begin
          for (forvar3242 = (1'h0); (forvar3242 < (2'h3)); forvar3242 = (forvar3242 + (1'h1)))
            begin
              reg3243 = $signed((reg14 ?
                  {"e4CmMoOi3Nw9QssH8"} : (|{$signed(wire3223)})));
              reg3244 <= (((-{(wire3217 && (8'ha5)),
                      reg12[(4'hb):(1'h1)]}) < (~^$signed((reg32 * reg33)))) ?
                  (((8'hb8) != "KAQolgMm5Mnze") ?
                      {"yvlwoFw",
                          (wire3227 + (reg23 ?
                              forvar24 : wire3219))} : (8'hb8)) : (((reg20 > (forvar30 ?
                              reg3231 : reg12)) ?
                          reg3232 : ((reg7 < reg12) < (reg6 + reg12))) ?
                      $signed($signed((reg6 - reg3237))) : ({reg21} & $unsigned(forvar4))));
            end
          reg3245 = (+($signed(((^forvar3230) ^ "vGiQttSLYRwXN9XEWX")) ~^ (reg3214[(2'h2):(1'h0)] ?
              $signed((!wire3221)) : ((^wire3229) ~^ forvar3242[(3'h5):(1'h0)]))));
          reg3246 = $signed($signed(forvar4));
          reg3247 <= $unsigned("hGCBw34UoZwx7BPxbV");
          reg3248 <= $signed(reg3236[(4'h8):(2'h3)]);
          reg3249 <= wire3216[(4'hb):(3'h6)];
        end
      else
        begin
          reg3242 <= "0e6qSd";
          reg3243 <= {(~&reg3236)};
          reg3244 <= (~&forvar13[(1'h0):(1'h0)]);
        end
      reg3250 <= ($signed(reg33[(4'hd):(1'h0)]) >> reg23[(2'h3):(2'h2)]);
      reg3251 = (^~forvar8[(4'h9):(4'h8)]);
    end
  module2028 modinst3253 (.wire2030(wire3212), .wire2031(wire3219), .clk(clk), .y(wire3252), .wire2029(reg3245), .wire2032(reg3241));
  assign wire3254 = (^{$unsigned($unsigned((^~reg28)))});
  always
    @(posedge clk) begin
      for (forvar3255 = (1'h0); (forvar3255 < (1'h1)); forvar3255 = (forvar3255 + (1'h1)))
        begin
          reg3256 <= ($signed((((8'hbb) || $unsigned(forvar24)) && reg27)) ?
              ((+reg3249[(4'hc):(3'h6)]) ?
                  $signed(wire3219[(1'h1):(1'h0)]) : $signed(((reg5 ?
                          reg3242 : (8'h9e)) ?
                      "XMz5or4rvPFMBd9Y3oZ" : $signed((8'hb0))))) : reg3241);
          for (forvar3257 = (1'h0); (forvar3257 < (3'h5)); forvar3257 = (forvar3257 + (1'h1)))
            begin
              reg3258 <= forvar17;
              reg3259 <= ($unsigned(forvar3230[(3'h5):(3'h5)]) - forvar3235);
              reg3260 <= (forvar3255[(5'h14):(1'h0)] ?
                  "NPX" : (&($unsigned("AXS1CGxFtBhXo23WOGu") >= (&reg3242[(3'h5):(2'h3)]))));
              reg3261 <= (!"BMvoZXqsMow3fGZ6");
              reg3262 <= $unsigned({(((8'hb3) != "Wwrofxw6CzfHfl") ?
                      reg3242[(2'h3):(2'h3)] : {(~&(7'h4a))}),
                  reg6[(4'hd):(3'h5)]});
              reg3263 <= (8'ha3);
            end
          reg3264 <= "7kUyLnlUfMC";
          reg3265 <= ((("Sm9fZ8DCxOA57G2ii7iaf0" <= $signed(reg7[(4'ha):(2'h3)])) ?
                  $unsigned((^~(wire3221 ?
                      reg29 : forvar30))) : $unsigned($unsigned((|forvar3230)))) ?
              ($unsigned((reg3232[(2'h2):(1'h0)] | reg3238[(1'h0):(1'h0)])) + reg3250[(4'hc):(4'h9)]) : ("xNFIeVOV4DBUN140zq3F4" < (~|$signed(reg3232))));
          reg3266 <= (&$signed((8'hae)));
          reg3267 <= reg9[(4'h8):(2'h3)];
        end
      reg3268 = "1Je6";
      reg3269 <= (reg31[(4'h9):(3'h6)] != (($signed(((8'hb0) ?
              forvar17 : reg18)) ?
          ((reg23 ? reg9 : wire0) ?
              (reg3263 ~^ reg5) : $signed(wire3219)) : (!(~|wire3216))) ^~ "KWWkSN84QPJrOyQwc"));
    end
  assign wire3270 = (((^$signed((7'h47))) == (~$signed((reg33 ?
                            reg11 : reg11)))) ?
                        $signed($signed(("" ?
                            reg22[(1'h0):(1'h0)] : {forvar30,
                                reg26}))) : $unsigned($unsigned("sw4CkRb7eWOs0DLMNkTNNgR")));
  assign wire3271 = (((~^reg3243) ?
                        wire3217[(4'hf):(4'hc)] : reg3232) ~^ forvar13[(1'h0):(1'h0)]);
  assign wire3272 = wire3223[(1'h1):(1'h1)];
  module662 modinst3274 (.wire663(forvar13), .y(wire3273), .wire665(reg20), .clk(clk), .wire667(reg10), .wire664(forvar8), .wire666(reg3249));
  always
    @(posedge clk) begin
      reg3275 <= (wire3254[(5'h11):(3'h5)] ?
          {{(~|((8'h9d) ? reg3258 : reg14))},
              $unsigned((reg3234 ?
                  $signed(reg3237) : (~&reg3237)))} : reg11[(3'h5):(2'h3)]);
      for (forvar3276 = (1'h0); (forvar3276 < (1'h1)); forvar3276 = (forvar3276 + (1'h1)))
        begin
          reg3277 <= (^$signed(reg3239[(4'h8):(3'h4)]));
          if (("Vk8Jw46BqK" ?
              "a4A8i1ECw1HGuaCv2gcH" : $unsigned(wire3223[(5'h16):(5'h15)])))
            begin
              reg3278 = (8'ha8);
              for (forvar3279 = (1'h0); (forvar3279 < (1'h1)); forvar3279 = (forvar3279 + (1'h1)))
                begin
                  reg3280 <= ((&($unsigned("uABigyDqDytTAyT") != "")) ?
                      (reg3247[(2'h3):(2'h3)] ?
                          "qqqZMHXcJyW2K1QyR3z" : (reg26 ?
                              $unsigned((~|reg3246)) : "")) : (wire3225 ?
                          $unsigned(((8'hb8) && (wire3210 - (8'hae)))) : {((wire3225 > wire3221) ~^ $unsigned(reg3233))}));
                  reg3281 = forvar3276[(3'h6):(2'h2)];
                  reg3282 <= (($unsigned("slFKQwzAoayl5NfAv2BDH") >>> ($unsigned("nOY") + {reg3238,
                      $signed(reg3237)})) >= $signed(wire3229[(5'h15):(3'h6)]));
                  reg3283 <= ((((8'hb5) ?
                          "DmoPaWbSunW4lOaxpOp" : (~&reg18)) && "6bQiMS") ?
                      wire2[(4'ha):(3'h4)] : "Z89hFpylns9");
                  reg3284 <= reg3282;
                  reg3285 = reg27;
                end
              reg3286 <= reg3249[(4'h9):(3'h6)];
              reg3287 <= ("iED8lHCL8sJpxi9IPKX" && $unsigned(reg3214));
              reg3288 <= (reg9 ? reg3251 : $unsigned(forvar8));
            end
          else
            begin
              for (forvar3278 = (1'h0); (forvar3278 < (3'h5)); forvar3278 = (forvar3278 + (1'h1)))
                begin
                  reg3279 <= "5Fo4GiP7SQ0o";
                  reg3280 <= reg3286;
                  reg3281 <= $signed($unsigned((~&$signed((wire1 ?
                      forvar3257 : reg28)))));
                  reg3282 <= "nZ2Hr7qoYhDO9x31lGJl";
                  reg3283 <= reg3248;
                  reg3284 <= ({(~(reg7 ?
                              $unsigned(reg3269) : (reg23 ?
                                  reg3287 : reg22)))} ?
                      {"SlolF920ZPGnGLe",
                          "UUIVIvuS2zU8"} : "4Qy6NMbVqTK77ELxAfwq");
                end
              reg3285 <= (reg3249 ?
                  reg25 : ("shv6GJfoL9n8nJIIKgc" == (reg3240[(3'h6):(3'h4)] - "")));
            end
          reg3289 <= $unsigned(forvar30[(5'h14):(4'h8)]);
          reg3290 <= (reg3244 ^ reg3243[(2'h2):(1'h0)]);
          for (forvar3291 = (1'h0); (forvar3291 < (2'h2)); forvar3291 = (forvar3291 + (1'h1)))
            begin
              reg3292 <= $unsigned((^~reg3268[(3'h4):(2'h3)]));
            end
          reg3293 = {"s7xfZHN0g7lDI77DztXIH8OT", "Gv57qNqDAui0Swm"};
        end
    end
  assign wire3294 = ((reg32[(4'hf):(3'h7)] ?
                            forvar30 : $signed($signed(wire3210))) ?
                        forvar3257 : $signed("oYdxGhrC9v3IqCSexim0"));
  always
    @(posedge clk) begin
      for (forvar3295 = (1'h0); (forvar3295 < (2'h2)); forvar3295 = (forvar3295 + (1'h1)))
        begin
          for (forvar3296 = (1'h0); (forvar3296 < (1'h0)); forvar3296 = (forvar3296 + (1'h1)))
            begin
              reg3297 <= $unsigned({{reg3279[(2'h3):(2'h3)]}});
              reg3298 <= ($unsigned((reg3231 - $signed($unsigned(reg3285)))) < forvar3257[(1'h0):(1'h0)]);
              reg3299 <= wire0;
              reg3300 <= ($signed($unsigned((~&(reg3283 ?
                  (8'h9f) : (7'h48))))) & reg12[(4'ha):(1'h0)]);
            end
          for (forvar3301 = (1'h0); (forvar3301 < (3'h5)); forvar3301 = (forvar3301 + (1'h1)))
            begin
              for (forvar3302 = (1'h0); (forvar3302 < (3'h4)); forvar3302 = (forvar3302 + (1'h1)))
                begin
                  reg3303 <= $signed((forvar3302 | $unsigned(("Rv7Rq56Xv1GwDR5G7DD6mfu4O" >= ((8'hb0) <<< reg20)))));
                  reg3304 <= reg20[(5'h12):(4'hd)];
                  reg3305 <= ($signed(((~^reg3290) <= (+$signed((8'ha6))))) < "k1koDOiVPx8lHBvTNn");
                  reg3306 <= $signed("JKmOnqaXd9");
                end
            end
          reg3307 <= $unsigned($unsigned("xcPMK8tD9pA3iTtGU"));
          reg3308 <= ({(^($unsigned(reg3306) | $unsigned(reg3262))),
              "YwkvgPq30LZFIXk6"} << $signed($signed(reg21)));
          for (forvar3309 = (1'h0); (forvar3309 < (2'h2)); forvar3309 = (forvar3309 + (1'h1)))
            begin
              for (forvar3310 = (1'h0); (forvar3310 < (1'h0)); forvar3310 = (forvar3310 + (1'h1)))
                begin
                  reg3311 <= $unsigned($signed(wire3272[(3'h6):(2'h2)]));
                  reg3312 <= reg3298[(4'hc):(3'h5)];
                  reg3313 <= wire1[(3'h4):(1'h0)];
                end
              reg3314 <= reg3298[(4'ha):(4'ha)];
              for (forvar3315 = (1'h0); (forvar3315 < (3'h4)); forvar3315 = (forvar3315 + (1'h1)))
                begin
                  reg3316 <= ({(((reg3261 ? forvar3257 : reg3247) ?
                              wire3219 : reg3287[(3'h4):(2'h3)]) ?
                          (8'h9c) : (8'ha4)),
                      reg9} < forvar3301);
                  reg3317 <= reg3238[(2'h2):(1'h1)];
                  reg3318 <= reg31[(4'hc):(3'h4)];
                  reg3319 <= $unsigned(wire3216[(2'h3):(1'h0)]);
                end
              reg3320 <= {((-reg3285[(3'h4):(1'h1)]) << {(wire3 * {reg3316,
                          reg3307})})};
            end
          reg3321 <= $signed(reg3260);
        end
      reg3322 <= "BtexY7bUS3YfwxpgVuF5iXKRf";
      reg3323 <= wire3216;
      reg3324 <= $unsigned((reg3239 ?
          reg3307 : $unsigned(reg3236[(1'h0):(1'h0)])));
      reg3325 <= $unsigned((^~(^~((~&reg33) ?
          (~|(8'hae)) : (reg3268 != wire2)))));
      reg3326 = {{(|reg3289[(4'ha):(3'h6)]),
              (reg17 ? reg26 : $unsigned($unsigned(reg3319)))}};
    end
  always
    @(posedge clk) begin
      reg3327 <= reg3260;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module34
#( parameter param3208 = {({(~^((8'hbc) < (8'ha8))), ((~(8'ha4)) - ((8'hbf) || (7'h40)))} & (+(((8'hba) ? (8'hae) : (7'h4b)) ? ((8'hbe) >= (8'ha0)) : ((7'h4d) == (8'hba))))), ((((-(8'hb9)) ? (~^(7'h44)) : ((8'hbc) ? (8'hb4) : (7'h41))) ? (8'hbc) : {((8'ha6) | (7'h48))}) ^ ((((7'h40) >>> (8'hbe)) > (8'hbf)) != (((7'h4a) >= (8'ha5)) | ((7'h49) ^ (8'h9f)))))}
, parameter param3209 = (((({param3208} > {param3208, param3208}) ? (~^param3208) : param3208) ? (param3208 ? (8'hb8) : ((param3208 ? param3208 : (8'hae)) | (param3208 | param3208))) : (~^(&(param3208 ? param3208 : param3208)))) && {{param3208}, (~|(((7'h4b) ? param3208 : param3208) ? ((8'h9f) ? param3208 : param3208) : (~^param3208)))}) )
(y, clk, wire39, wire38, wire37, wire36, wire35);
  output wire [(32'h60f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h17):(1'h0)] wire39;
  input wire [(5'h10):(1'h0)] wire38;
  input wire signed [(5'h17):(1'h0)] wire37;
  input wire [(5'h1a):(1'h0)] wire36;
  input wire signed [(5'h19):(1'h0)] wire35;
  reg signed [(5'h10):(1'h0)] reg3207 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3206 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3205 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3204 = (1'h0);
  reg [(4'h8):(1'h0)] reg3203 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3202 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3201 = (1'h0);
  reg [(4'he):(1'h0)] forvar3200 = (1'h0);
  reg [(4'hf):(1'h0)] reg3199 = (1'h0);
  reg [(5'h17):(1'h0)] reg3198 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3197 = (1'h0);
  reg [(5'h12):(1'h0)] reg3196 = (1'h0);
  reg [(5'h11):(1'h0)] reg3195 = (1'h0);
  reg [(4'hc):(1'h0)] reg3194 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3193 = (1'h0);
  reg [(5'h15):(1'h0)] reg3192 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar3191 = (1'h0);
  reg [(5'h13):(1'h0)] reg3190 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3189 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3188 = (1'h0);
  wire [(5'h15):(1'h0)] wire3176;
  wire signed [(5'h15):(1'h0)] wire3172;
  wire [(5'h15):(1'h0)] wire3171;
  wire [(5'h13):(1'h0)] wire3163;
  wire [(5'h14):(1'h0)] wire3162;
  wire [(5'h10):(1'h0)] wire3160;
  wire signed [(5'h17):(1'h0)] wire3102;
  wire [(5'h19):(1'h0)] wire40;
  wire [(5'h17):(1'h0)] wire3104;
  reg [(4'hd):(1'h0)] forvar3106 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3107 = (1'h0);
  reg [(4'hf):(1'h0)] reg3108 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3109 = (1'h0);
  reg [(5'h19):(1'h0)] reg3110 = (1'h0);
  reg [(3'h4):(1'h0)] reg3111 = (1'h0);
  reg [(5'h14):(1'h0)] reg3112 = (1'h0);
  reg [(4'hc):(1'h0)] reg3113 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3114 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3115 = (1'h0);
  reg [(5'h17):(1'h0)] reg3116 = (1'h0);
  reg [(4'hc):(1'h0)] reg3117 = (1'h0);
  reg [(5'h16):(1'h0)] reg3118 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3119 = (1'h0);
  reg [(4'hc):(1'h0)] reg3120 = (1'h0);
  reg [(2'h3):(1'h0)] reg3121 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar3122 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3123 = (1'h0);
  reg [(5'h1a):(1'h0)] reg3124 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3125 = (1'h0);
  reg [(5'h19):(1'h0)] reg3126 = (1'h0);
  reg [(5'h13):(1'h0)] reg3127 = (1'h0);
  reg [(4'he):(1'h0)] reg3128 = (1'h0);
  reg [(4'hb):(1'h0)] reg3129 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3130 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3131 = (1'h0);
  reg [(5'h18):(1'h0)] reg3132 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3133 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3134 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3135 = (1'h0);
  reg [(4'hd):(1'h0)] reg3136 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3137 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3138 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar3139 = (1'h0);
  reg [(5'h17):(1'h0)] forvar3140 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3141 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3142 = (1'h0);
  reg [(5'h17):(1'h0)] reg3143 = (1'h0);
  reg [(5'h19):(1'h0)] reg3144 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar3145 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3146 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3147 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3148 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3149 = (1'h0);
  reg [(5'h17):(1'h0)] reg3150 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar3151 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3152 = (1'h0);
  reg [(5'h14):(1'h0)] reg3153 = (1'h0);
  reg [(2'h2):(1'h0)] reg3154 = (1'h0);
  reg [(5'h12):(1'h0)] reg3155 = (1'h0);
  reg [(5'h15):(1'h0)] reg3156 = (1'h0);
  reg [(4'hb):(1'h0)] reg3157 = (1'h0);
  wire [(3'h4):(1'h0)] wire3158;
  reg [(4'h8):(1'h0)] reg3165 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3166 = (1'h0);
  reg [(5'h11):(1'h0)] reg3167 = (1'h0);
  reg [(3'h4):(1'h0)] reg3168 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire3169;
  wire signed [(5'h12):(1'h0)] wire3174;
  wire [(5'h15):(1'h0)] wire3178;
  wire signed [(3'h4):(1'h0)] wire3180;
  wire [(4'ha):(1'h0)] wire3182;
  wire signed [(5'h19):(1'h0)] wire3184;
  wire signed [(2'h2):(1'h0)] wire3186;
  assign y = {reg3207,
                 reg3206,
                 reg3205,
                 reg3204,
                 reg3203,
                 forvar3202,
                 reg3201,
                 forvar3200,
                 reg3199,
                 reg3198,
                 reg3197,
                 reg3196,
                 reg3195,
                 reg3194,
                 forvar3193,
                 reg3192,
                 forvar3191,
                 reg3190,
                 forvar3189,
                 reg3188,
                 wire3176,
                 wire3172,
                 wire3171,
                 wire3163,
                 wire3162,
                 wire3160,
                 wire3102,
                 wire40,
                 wire3104,
                 forvar3106,
                 forvar3107,
                 reg3108,
                 forvar3109,
                 reg3110,
                 reg3111,
                 reg3112,
                 reg3113,
                 forvar3114,
                 reg3115,
                 reg3116,
                 reg3117,
                 reg3118,
                 forvar3119,
                 reg3120,
                 reg3121,
                 forvar3122,
                 reg3123,
                 reg3124,
                 reg3125,
                 reg3126,
                 reg3127,
                 reg3128,
                 reg3129,
                 reg3130,
                 reg3131,
                 reg3132,
                 reg3133,
                 reg3134,
                 forvar3135,
                 reg3136,
                 reg3137,
                 reg3138,
                 forvar3139,
                 forvar3140,
                 reg3141,
                 reg3142,
                 reg3143,
                 reg3144,
                 forvar3145,
                 reg3146,
                 reg3147,
                 reg3148,
                 reg3149,
                 reg3150,
                 forvar3151,
                 reg3152,
                 reg3153,
                 reg3154,
                 reg3155,
                 reg3156,
                 reg3157,
                 wire3158,
                 reg3165,
                 reg3166,
                 reg3167,
                 reg3168,
                 wire3169,
                 wire3174,
                 wire3178,
                 wire3180,
                 wire3182,
                 wire3184,
                 wire3186,
                 (1'h0)};
  assign wire40 = (((({(8'ha7)} ? wire37 : wire38[(3'h4):(3'h4)]) ?
                              (wire36[(4'hb):(2'h3)] <<< (wire35 > wire38)) : "nV71") ?
                          wire36[(1'h1):(1'h0)] : (wire38[(1'h0):(1'h0)] ?
                              (-(wire39 != wire39)) : $unsigned($signed(wire36)))) ?
                      ({$signed(wire39[(5'h14):(4'hd)]), "IwNRl5IDgzkgXo"} ?
                          "kdpt" : $signed({(wire36 ? wire37 : (8'ha9)),
                              (~wire35)})) : (~&wire39));
  module41 modinst3103 (wire3102, clk, wire36, wire39, wire40, wire37, wire35);
  module48 modinst3105 (wire3104, clk, wire35, wire36, wire40, wire38);
  always
    @(posedge clk) begin
      for (forvar3106 = (1'h0); (forvar3106 < (2'h3)); forvar3106 = (forvar3106 + (1'h1)))
        begin
          for (forvar3107 = (1'h0); (forvar3107 < (2'h3)); forvar3107 = (forvar3107 + (1'h1)))
            begin
              reg3108 <= ((wire39[(4'ha):(2'h2)] ?
                      "2BaNFKtPr8nVfnDpIv" : (~"bDFO19CvMxrkOor")) ?
                  "Gkfmx" : (^"XkD3AVCoo1gRLaMqy4RpZ6i"));
              for (forvar3109 = (1'h0); (forvar3109 < (3'h5)); forvar3109 = (forvar3109 + (1'h1)))
                begin
                  reg3110 <= $signed($signed(($unsigned($unsigned(wire3104)) ?
                      (~&((8'hbc) ^~ (8'hb6))) : wire37)));
                end
              reg3111 <= (~|(($unsigned({reg3108, (8'hbf)}) ?
                      (~^(^~forvar3106)) : $unsigned($unsigned(forvar3106))) ?
                  "wqfqO6fKcfZovSkuefQqTdm" : ((^(wire3102 & wire3104)) ?
                      (|{wire35,
                          wire35}) : ($unsigned((8'hb3)) ~^ $signed(wire40)))));
              reg3112 <= $signed((({(wire37 ? wire39 : forvar3107)} >> wire38) ?
                  $signed($unsigned(wire36)) : wire35));
              reg3113 <= "vEkK";
              for (forvar3114 = (1'h0); (forvar3114 < (3'h5)); forvar3114 = (forvar3114 + (1'h1)))
                begin
                  reg3115 <= forvar3114;
                end
            end
        end
      reg3116 <= reg3112[(5'h10):(4'hc)];
      reg3117 <= ("zvosDrOm6nGVJL07Lz31MT" ?
          (-$signed((|(~|reg3115)))) : {forvar3109[(4'h9):(3'h5)],
              (wire35[(1'h1):(1'h1)] ?
                  {(~forvar3107),
                      ((8'haf) ?
                          wire37 : (8'hbf))} : ($unsigned((8'h9e)) ^ forvar3109))});
      reg3118 = $unsigned((reg3108[(4'h9):(2'h3)] > forvar3106[(4'hc):(3'h7)]));
      for (forvar3119 = (1'h0); (forvar3119 < (3'h5)); forvar3119 = (forvar3119 + (1'h1)))
        begin
          reg3120 <= reg3117;
          reg3121 <= $unsigned(forvar3114);
          for (forvar3122 = (1'h0); (forvar3122 < (1'h1)); forvar3122 = (forvar3122 + (1'h1)))
            begin
              reg3123 <= $signed($unsigned((8'haa)));
              reg3124 <= reg3116;
              reg3125 = "IMEOX7W9FKKFb1VAAw6yN";
              reg3126 <= $signed(reg3113);
              reg3127 = wire35[(4'h9):(3'h7)];
              reg3128 <= $signed($unsigned($signed((reg3108 ?
                  (&reg3124) : (~wire3104)))));
            end
          reg3129 = wire35[(4'hf):(1'h0)];
          reg3130 <= "Ga";
        end
      reg3131 <= (($signed($signed((reg3126 ? reg3115 : reg3115))) ?
              ("tS8ic5o2DAtsn" ?
                  reg3127 : {"CWP91LMybivAnXwFbc7ERxTc"}) : "FUPEBqi") ?
          $unsigned(($unsigned({(8'hb3),
              reg3124}) + "AyuBuAnnMa")) : (&$unsigned($unsigned(forvar3122[(1'h1):(1'h1)]))));
    end
  always
    @(posedge clk) begin
      reg3132 <= ("ahZ6UP4oc9Thk7909T" ? "1RLXuNOEl977YN" : "bNkxxU");
      reg3133 <= ((8'hbe) ?
          {((^wire38) ~^ ($signed(reg3115) ?
                  (!reg3131) : ((8'hba) ~^ wire37)))} : {(~^(reg3131 ?
                  reg3125 : $unsigned(reg3110)))});
      reg3134 = "dW4iVume4NKx1zaUshwoNVL9e";
      for (forvar3135 = (1'h0); (forvar3135 < (2'h2)); forvar3135 = (forvar3135 + (1'h1)))
        begin
          reg3136 <= ((~|"RGG7VbpQK3XNwk0OdD72sJn6Q") && (~^reg3130));
          reg3137 <= reg3118;
          reg3138 <= ($signed({$signed($signed(reg3113)), reg3116}) ?
              reg3134[(5'h12):(5'h10)] : {"D3"});
          for (forvar3139 = (1'h0); (forvar3139 < (3'h4)); forvar3139 = (forvar3139 + (1'h1)))
            begin
              for (forvar3140 = (1'h0); (forvar3140 < (3'h4)); forvar3140 = (forvar3140 + (1'h1)))
                begin
                  reg3141 <= wire39;
                  reg3142 <= (|reg3133[(3'h6):(2'h2)]);
                  reg3143 <= $unsigned(forvar3114[(1'h1):(1'h1)]);
                end
              reg3144 <= wire35[(5'h19):(1'h0)];
              for (forvar3145 = (1'h0); (forvar3145 < (1'h1)); forvar3145 = (forvar3145 + (1'h1)))
                begin
                  reg3146 <= reg3138[(4'ha):(2'h3)];
                  reg3147 = $unsigned($unsigned(forvar3122));
                  reg3148 <= "NlaDRv3rG21xUT2I3xPtR";
                  reg3149 <= ("KiIG" ^ ((reg3124 >= forvar3122[(1'h0):(1'h0)]) != (~|((reg3133 ?
                          reg3120 : forvar3140) ?
                      reg3147[(5'h14):(3'h6)] : reg3128[(1'h1):(1'h0)]))));
                  reg3150 = (reg3115 ? (7'h4a) : "iQQJ7keWsWf0ymHs0DUMIt8S");
                end
              for (forvar3151 = (1'h0); (forvar3151 < (3'h5)); forvar3151 = (forvar3151 + (1'h1)))
                begin
                  reg3152 <= $unsigned(wire39);
                  reg3153 <= {"VDmtNiGgt9bdL144M"};
                end
              reg3154 <= forvar3151[(2'h3):(2'h2)];
              reg3155 <= "yZyaw1RoAeDvKH1Bw";
            end
        end
      reg3156 = ($signed(($signed("dMzUYvsdPh85") ?
              (+(reg3131 ?
                  reg3137 : reg3150)) : ($unsigned(reg3149) >= (&reg3134)))) ?
          $signed((("8JTL" ?
              forvar3151 : $unsigned(forvar3119)) ^~ "22961YVbwYJGOdLiD1K4yfW77")) : reg3116[(4'he):(3'h7)]);
    end
  always
    @(posedge clk) begin
      reg3157 <= $signed((-({$signed(reg3143)} <<< (^"OYbR"))));
    end
  module1953 modinst3159 (.wire1958(reg3141), .clk(clk), .wire1957(wire38), .wire1955(reg3156), .wire1956(reg3115), .y(wire3158), .wire1954(forvar3140));
  module1383 modinst3161 (.wire1386(reg3124), .clk(clk), .wire1384(wire36), .y(wire3160), .wire1387(reg3127), .wire1385(wire3102));
  assign wire3162 = wire3160[(1'h0):(1'h0)];
  module76 modinst3164 (.wire80(reg3124), .wire78(wire36), .y(wire3163), .wire79(reg3153), .clk(clk), .wire77(reg3115), .wire81(reg3155));
  always
    @(posedge clk) begin
      reg3165 <= ({(({reg3125} <<< (reg3116 ?
              reg3115 : (8'hb0))) == wire3102[(5'h17):(5'h17)]),
          ($unsigned("1LyfJ") <<< (^((7'h41) || wire38)))} || "dhEKL6vMc4");
      reg3166 <= (~&($unsigned((wire3160 ?
              (forvar3106 ? reg3134 : (8'ha4)) : (reg3143 ?
                  wire3102 : forvar3139))) ?
          wire38 : $unsigned(reg3136[(4'h9):(2'h2)])));
      reg3167 <= (&"aZWzxpmSBDObbuKRLqfKo");
      reg3168 <= wire39[(5'h17):(4'h8)];
    end
  module957 modinst3170 (wire3169, clk, wire39, forvar3151, wire3162, reg3155, reg3123);
  assign wire3171 = $unsigned((^~reg3148[(5'h10):(2'h3)]));
  module2707 modinst3173 (.wire2711(reg3150), .y(wire3172), .wire2712(wire3102), .clk(clk), .wire2710(reg3142), .wire2708(forvar3122), .wire2709(reg3124));
  module217 modinst3175 (.wire219(forvar3109), .wire220(wire35), .y(wire3174), .wire221(reg3153), .wire222(reg3123), .clk(clk), .wire218(reg3117));
  module957 modinst3177 (wire3176, clk, reg3129, reg3131, reg3153, reg3127, reg3142);
  module690 modinst3179 (.wire691(forvar3145), .wire694(reg3118), .y(wire3178), .wire693(reg3112), .clk(clk), .wire692(reg3132));
  module1383 modinst3181 (.wire1385(wire35), .wire1386(reg3129), .clk(clk), .y(wire3180), .wire1384(wire39), .wire1387(reg3137));
  module492 modinst3183 (wire3182, clk, wire3163, wire3174, wire3160, reg3138);
  module2592 modinst3185 (.y(wire3184), .wire2593(wire3171), .clk(clk), .wire2594(wire36), .wire2596(wire3176), .wire2595(reg3167));
  module54 modinst3187 (wire3186, clk, reg3146, forvar3145, forvar3140, reg3130, reg3149);
  always
    @(posedge clk) begin
      reg3188 = $unsigned(({((reg3125 ^ reg3156) ?
                  reg3128[(2'h3):(2'h2)] : reg3136)} ?
          $signed(($signed(reg3142) ?
              "2Kn0U0sW" : (reg3129 ?
                  wire3186 : reg3121))) : $signed($signed((+reg3118)))));
      for (forvar3189 = (1'h0); (forvar3189 < (3'h5)); forvar3189 = (forvar3189 + (1'h1)))
        begin
          reg3190 <= reg3118;
          for (forvar3191 = (1'h0); (forvar3191 < (2'h2)); forvar3191 = (forvar3191 + (1'h1)))
            begin
              reg3192 <= $signed(forvar3145);
            end
        end
      for (forvar3193 = (1'h0); (forvar3193 < (3'h5)); forvar3193 = (forvar3193 + (1'h1)))
        begin
          reg3194 = (~wire3176[(4'h9):(2'h2)]);
          reg3195 = (^{$unsigned(("RZ3ITxUuUeC" ?
                  ((8'hb7) >>> wire3184) : reg3165[(3'h6):(3'h5)])),
              "7ver2le7Nxa5asB"});
          reg3196 <= reg3132;
          reg3197 = "nkt3z0l2PzQC7bL18EtxPgAvV";
        end
      reg3198 = (^($signed((-wire3172[(5'h15):(4'he)])) ?
          "qHHyRIfKBeJK4Cu46oiTMH" : ((^~$unsigned(forvar3107)) ?
              ($unsigned(wire3180) ?
                  $signed(reg3167) : $unsigned(wire3162)) : $signed((reg3113 * wire40)))));
    end
  always
    @(posedge clk) begin
      reg3199 <= (wire3171[(3'h5):(2'h3)] ? reg3194 : "PMzCL84f5lmIW");
      for (forvar3200 = (1'h0); (forvar3200 < (1'h0)); forvar3200 = (forvar3200 + (1'h1)))
        begin
          reg3201 <= $signed(forvar3107);
          for (forvar3202 = (1'h0); (forvar3202 < (3'h5)); forvar3202 = (forvar3202 + (1'h1)))
            begin
              reg3203 <= $unsigned("4gTLTD2xC64s");
              reg3204 <= $unsigned((+(~$unsigned((forvar3202 >= reg3143)))));
              reg3205 = (({((forvar3109 ? reg3110 : reg3127) >= (7'h46))} ?
                      $signed((8'h9d)) : {forvar3109[(3'h6):(2'h2)],
                          wire3102}) ?
                  ((reg3144[(4'h8):(1'h1)] >> wire3102[(3'h4):(1'h0)]) ?
                      "MZF" : $signed($unsigned(forvar3107))) : "Bulvtkms");
            end
          reg3206 <= "NhHfNxnE";
        end
      reg3207 <= reg3198;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module41
#( parameter param3100 = (~(((((8'hb5) ? (8'hb3) : (8'ha7)) ? ((8'haa) >>> (7'h46)) : (!(8'h9f))) ? (!((8'h9e) ? (8'ha4) : (8'h9d))) : (((8'hb0) ? (8'ha5) : (7'h46)) + ((8'hb2) ~^ (8'ha1)))) | (8'hb2)))
, parameter param3101 = (-(!(((param3100 ? param3100 : param3100) << ((8'haf) ? param3100 : param3100)) ? (~&{param3100, param3100}) : (7'h4d)))) )
(y, clk, wire42, wire43, wire44, wire45, wire46);
  output wire [(32'h446):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire42;
  input wire signed [(5'h17):(1'h0)] wire43;
  input wire [(5'h19):(1'h0)] wire44;
  input wire [(5'h17):(1'h0)] wire45;
  input wire [(5'h19):(1'h0)] wire46;
  reg signed [(5'h10):(1'h0)] reg3099 = (1'h0);
  wire [(3'h7):(1'h0)] wire3095;
  wire [(5'h14):(1'h0)] wire3094;
  reg signed [(2'h2):(1'h0)] reg3093 = (1'h0);
  reg [(5'h12):(1'h0)] reg3092 = (1'h0);
  reg [(5'h14):(1'h0)] reg3091 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3090 = (1'h0);
  wire [(5'h11):(1'h0)] wire3076;
  wire signed [(3'h6):(1'h0)] wire3075;
  reg [(5'h19):(1'h0)] reg3074 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3073 = (1'h0);
  reg [(5'h15):(1'h0)] reg3072 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar3071 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3063 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar3060 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3057 = (1'h0);
  reg [(5'h11):(1'h0)] reg3070 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3069 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg3068 = (1'h0);
  reg [(5'h11):(1'h0)] reg3067 = (1'h0);
  reg [(5'h19):(1'h0)] reg3066 = (1'h0);
  reg [(5'h19):(1'h0)] reg3065 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3064 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar3063 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3062 = (1'h0);
  reg [(5'h13):(1'h0)] reg3061 = (1'h0);
  reg [(5'h11):(1'h0)] reg3060 = (1'h0);
  reg [(5'h18):(1'h0)] reg3059 = (1'h0);
  reg [(4'hf):(1'h0)] reg3058 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3057 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3056 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3055 = (1'h0);
  reg [(5'h16):(1'h0)] reg3054 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg3053 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3052 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg3051 = (1'h0);
  reg [(5'h11):(1'h0)] reg3050 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar3049 = (1'h0);
  reg [(5'h15):(1'h0)] reg3048 = (1'h0);
  reg [(2'h3):(1'h0)] reg3047 = (1'h0);
  reg [(5'h17):(1'h0)] forvar3046 = (1'h0);
  reg [(4'h8):(1'h0)] reg3045 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3044 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3043 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3042 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3041 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3040 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg3039 = (1'h0);
  reg [(4'ha):(1'h0)] reg3038 = (1'h0);
  reg [(5'h13):(1'h0)] reg3037 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3036 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg3035 = (1'h0);
  wire [(5'h1a):(1'h0)] wire47;
  wire [(4'hc):(1'h0)] wire3031;
  wire [(5'h17):(1'h0)] wire3033;
  wire signed [(5'h19):(1'h0)] wire3078;
  wire signed [(5'h14):(1'h0)] wire3080;
  wire signed [(5'h19):(1'h0)] wire3082;
  reg [(4'h9):(1'h0)] reg3084 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire3085;
  wire [(5'h1a):(1'h0)] wire3087;
  wire signed [(2'h3):(1'h0)] wire3088;
  wire [(5'h14):(1'h0)] wire3097;
  assign y = {reg3099,
                 wire3095,
                 wire3094,
                 reg3093,
                 reg3092,
                 reg3091,
                 reg3090,
                 wire3076,
                 wire3075,
                 reg3074,
                 reg3073,
                 reg3072,
                 forvar3071,
                 reg3063,
                 forvar3060,
                 reg3057,
                 reg3070,
                 reg3069,
                 reg3068,
                 reg3067,
                 reg3066,
                 reg3065,
                 reg3064,
                 forvar3063,
                 reg3062,
                 reg3061,
                 reg3060,
                 reg3059,
                 reg3058,
                 forvar3057,
                 reg3056,
                 forvar3055,
                 reg3054,
                 reg3053,
                 reg3052,
                 reg3051,
                 reg3050,
                 forvar3049,
                 reg3048,
                 reg3047,
                 forvar3046,
                 reg3045,
                 reg3044,
                 reg3043,
                 reg3042,
                 reg3041,
                 forvar3040,
                 reg3039,
                 reg3038,
                 reg3037,
                 reg3036,
                 reg3035,
                 wire47,
                 wire3031,
                 wire3033,
                 wire3078,
                 wire3080,
                 wire3082,
                 reg3084,
                 wire3085,
                 wire3087,
                 wire3088,
                 wire3097,
                 (1'h0)};
  assign wire47 = wire44;
  module48 modinst3032 (.wire50(wire43), .wire52(wire44), .y(wire3031), .clk(clk), .wire49(wire46), .wire51(wire47));
  module2538 modinst3034 (wire3033, clk, wire45, wire47, wire3031, wire43, wire46);
  always
    @(posedge clk) begin
      reg3035 = "R5rnzEB3niatRd";
      reg3036 <= $signed($signed({wire47[(4'h9):(1'h1)]}));
      reg3037 = wire45;
      reg3038 <= (8'h9c);
      reg3039 <= wire3033;
    end
  always
    @(posedge clk) begin
      for (forvar3040 = (1'h0); (forvar3040 < (2'h2)); forvar3040 = (forvar3040 + (1'h1)))
        begin
          reg3041 <= $unsigned((&(($unsigned(wire43) && reg3035) == ("UlrSbNVyAviwsONW" * "4RVbbL1fk5T"))));
          reg3042 <= (~|reg3036[(3'h5):(3'h4)]);
          reg3043 <= $signed({$unsigned($signed($unsigned(reg3039))),
              "IeOCuRDwB2eE"});
          reg3044 <= reg3035;
        end
      reg3045 = (8'hb5);
      for (forvar3046 = (1'h0); (forvar3046 < (1'h0)); forvar3046 = (forvar3046 + (1'h1)))
        begin
          reg3047 <= reg3038;
          reg3048 <= ($signed(wire42) * wire47[(2'h3):(2'h3)]);
          for (forvar3049 = (1'h0); (forvar3049 < (2'h3)); forvar3049 = (forvar3049 + (1'h1)))
            begin
              reg3050 = (8'hb6);
              reg3051 <= (-$unsigned("8UIdPId8k39"));
              reg3052 = (($signed(reg3044) < wire47) >>> forvar3046[(1'h0):(1'h0)]);
              reg3053 <= (+(forvar3049[(1'h1):(1'h1)] ? reg3048 : (8'hb3)));
              reg3054 <= "YCqT4OANAeoWNuztkwQBzWtm";
            end
          for (forvar3055 = (1'h0); (forvar3055 < (3'h4)); forvar3055 = (forvar3055 + (1'h1)))
            begin
              reg3056 <= $unsigned($unsigned($signed("IEL3")));
            end
          if ("tJUERQwzeAXBmNmsZb51cLJ")
            begin
              for (forvar3057 = (1'h0); (forvar3057 < (3'h5)); forvar3057 = (forvar3057 + (1'h1)))
                begin
                  reg3058 <= (-"MM6AAsmhY9OcF1ILeI4");
                  reg3059 = $signed("JfC8ZfEz6r6mLfJtBb");
                  reg3060 <= reg3047[(1'h0):(1'h0)];
                  reg3061 <= reg3056[(5'h12):(4'h9)];
                  reg3062 <= {wire42, "dTpoZuoRG0OFv5vQGO1gW5uA"};
                end
              for (forvar3063 = (1'h0); (forvar3063 < (2'h3)); forvar3063 = (forvar3063 + (1'h1)))
                begin
                  reg3064 <= (-"PWXn0YK4AnV");
                  reg3065 = reg3047[(1'h1):(1'h1)];
                  reg3066 <= (reg3050[(4'h8):(3'h6)] >= (8'hac));
                  reg3067 <= ((+{(^~wire46)}) ?
                      $signed((~|("3xuL9SkS97kpbcegbC" || (reg3062 ?
                          (8'h9d) : reg3035)))) : (~&reg3054[(2'h2):(1'h1)]));
                  reg3068 = $signed($signed((~(wire3031[(4'ha):(4'h9)] ?
                      {reg3065} : reg3047[(1'h1):(1'h1)]))));
                  reg3069 <= $signed((~&($unsigned($unsigned(forvar3049)) - reg3047)));
                end
              reg3070 = $unsigned((^~$unsigned($unsigned((reg3042 <<< reg3036)))));
            end
          else
            begin
              reg3057 <= forvar3049[(2'h2):(1'h0)];
              reg3058 = (reg3059[(5'h17):(5'h11)] ?
                  ((wire42 ?
                      ($signed(reg3068) ?
                          (forvar3049 ?
                              reg3062 : reg3037) : (~&reg3057)) : {"C5pBwypBAFlDQtzOsxk6lDDH"}) ^~ reg3043) : ($unsigned(($unsigned(reg3069) ?
                          wire44 : {reg3051})) ?
                      wire3031[(3'h5):(1'h0)] : $unsigned($signed(reg3060))));
              reg3059 <= reg3047;
              for (forvar3060 = (1'h0); (forvar3060 < (1'h1)); forvar3060 = (forvar3060 + (1'h1)))
                begin
                  reg3061 = {($unsigned("0zdwwiNR9B0D8eJwboLK3B") >>> reg3058),
                      {$unsigned($unsigned((reg3057 ^ forvar3049))),
                          (({wire42, reg3036} ^ (!reg3053)) ?
                              (^~$signed(wire44)) : ((reg3051 || reg3069) ?
                                  (&reg3058) : (reg3065 || reg3054)))}};
                end
              reg3062 = (^reg3070[(1'h1):(1'h0)]);
              reg3063 = (~reg3064[(1'h0):(1'h0)]);
            end
        end
      for (forvar3071 = (1'h0); (forvar3071 < (3'h4)); forvar3071 = (forvar3071 + (1'h1)))
        begin
          reg3072 <= {(-$unsigned($unsigned(reg3044[(3'h4):(1'h1)])))};
          reg3073 = reg3059[(4'hf):(4'h9)];
          reg3074 <= {(~&("Mom" & (reg3072 & reg3041)))};
        end
    end
  assign wire3075 = reg3060[(3'h4):(2'h2)];
  module1146 modinst3077 (wire3076, clk, reg3074, reg3037, reg3035, reg3039, reg3054);
  module224 modinst3079 (wire3078, clk, reg3054, reg3070, reg3061, wire45);
  module435 modinst3081 (wire3080, clk, reg3047, reg3048, forvar3046, wire3076);
  module757 modinst3083 (wire3082, clk, reg3069, forvar3046, forvar3049, reg3037);
  always
    @(posedge clk) begin
      reg3084 = reg3035[(5'h12):(5'h11)];
    end
  module2592 modinst3086 (.wire2593(wire44), .wire2595(reg3062), .clk(clk), .wire2594(reg3041), .y(wire3085), .wire2596(reg3050));
  assign wire3087 = (~^"XQWu8X6Me4kKh");
  module2538 modinst3089 (wire3088, clk, wire3033, reg3053, wire42, wire3082, reg3066);
  always
    @(posedge clk) begin
      reg3090 <= "yvQ7mxSnLuAN1Q";
      reg3091 <= $unsigned(((forvar3057 <<< {"AYtMUKmQZGbI"}) ?
          ({forvar3046, "BNnBqbsA6G7OIq0QHoeWk"} ?
              (reg3042 == (^~(7'h45))) : (~|{reg3044, (8'ha6)})) : (+reg3072)));
      reg3092 <= (^~"xpNIr");
      reg3093 = reg3051;
    end
  assign wire3094 = reg3070;
  module76 modinst3096 (wire3095, clk, wire42, reg3090, reg3067, wire3080, reg3092);
  module2538 modinst3098 (.wire2541(wire42), .wire2542(reg3039), .wire2543(wire3087), .wire2539(reg3074), .y(wire3097), .clk(clk), .wire2540(reg3058));
  always
    @(posedge clk) begin
      reg3099 <= (+reg3045);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module48  (y, clk, wire52, wire51, wire50, wire49);
  output wire [(32'h615):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h19):(1'h0)] wire52;
  input wire [(5'h1a):(1'h0)] wire51;
  input wire signed [(5'h17):(1'h0)] wire50;
  input wire signed [(5'h10):(1'h0)] wire49;
  reg signed [(2'h3):(1'h0)] reg3030 = (1'h0);
  reg [(2'h2):(1'h0)] reg3029 = (1'h0);
  reg [(5'h19):(1'h0)] reg3028 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3027 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3026 = (1'h0);
  reg [(5'h17):(1'h0)] forvar3025 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3024 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3023 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3022 = (1'h0);
  reg [(3'h6):(1'h0)] reg3021 = (1'h0);
  reg [(3'h7):(1'h0)] reg3020 = (1'h0);
  reg [(4'hd):(1'h0)] reg3019 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg3018 = (1'h0);
  reg [(4'hc):(1'h0)] reg3017 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg3016 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3015 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3014 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3013 = (1'h0);
  reg [(5'h16):(1'h0)] forvar3012 = (1'h0);
  reg [(3'h4):(1'h0)] reg3011 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3010 = (1'h0);
  reg [(4'ha):(1'h0)] reg3009 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg3008 = (1'h0);
  reg [(4'hf):(1'h0)] reg3007 = (1'h0);
  wire [(5'h19):(1'h0)] wire3006;
  reg signed [(5'h15):(1'h0)] reg3005 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3004 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg3003 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire3001;
  wire signed [(4'h9):(1'h0)] wire3000;
  reg signed [(3'h6):(1'h0)] reg2999 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2998 = (1'h0);
  reg [(5'h18):(1'h0)] reg2997 = (1'h0);
  reg [(2'h3):(1'h0)] reg2996 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2995 = (1'h0);
  reg [(4'h9):(1'h0)] reg2994 = (1'h0);
  reg [(5'h18):(1'h0)] reg2993 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2992 = (1'h0);
  reg [(3'h7):(1'h0)] reg2991 = (1'h0);
  reg [(4'ha):(1'h0)] reg2990 = (1'h0);
  reg [(4'he):(1'h0)] forvar2989 = (1'h0);
  reg [(3'h7):(1'h0)] reg2988 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2987 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2986 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2985 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2984 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2983 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar2982 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2981 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2980 = (1'h0);
  reg [(4'he):(1'h0)] reg2979 = (1'h0);
  reg [(5'h10):(1'h0)] reg2978 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2977 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2976 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2975 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2974 = (1'h0);
  reg [(3'h5):(1'h0)] reg2973 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2972 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2971 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2970 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2969 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2968 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2967 = (1'h0);
  reg [(5'h15):(1'h0)] reg2966 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2965 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2964 = (1'h0);
  reg [(5'h14):(1'h0)] reg2963 = (1'h0);
  reg [(4'hb):(1'h0)] reg2962 = (1'h0);
  reg [(5'h12):(1'h0)] reg2961 = (1'h0);
  reg [(2'h2):(1'h0)] reg2960 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2956 = (1'h0);
  reg [(3'h4):(1'h0)] reg2959 = (1'h0);
  reg [(5'h12):(1'h0)] reg2958 = (1'h0);
  reg [(5'h19):(1'h0)] reg2957 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2956 = (1'h0);
  reg [(4'h9):(1'h0)] reg2955 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2954 = (1'h0);
  reg [(5'h14):(1'h0)] reg2953 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2952 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2951 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2950 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2949 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2948 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2947 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2946 = (1'h0);
  reg [(4'hf):(1'h0)] reg2945 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2944 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2943 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar2942 = (1'h0);
  reg [(3'h7):(1'h0)] reg2941 = (1'h0);
  reg [(5'h18):(1'h0)] reg2940 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2939 = (1'h0);
  reg [(5'h12):(1'h0)] reg2938 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2937 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar2936 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2935 = (1'h0);
  wire [(5'h1a):(1'h0)] wire2919;
  wire signed [(5'h10):(1'h0)] wire53;
  wire [(5'h16):(1'h0)] wire2921;
  reg signed [(5'h15):(1'h0)] reg2923 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2924 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2925 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2926 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2927 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2928 = (1'h0);
  wire [(5'h13):(1'h0)] wire2929;
  wire signed [(2'h2):(1'h0)] wire2930;
  wire signed [(5'h15):(1'h0)] wire2932;
  wire signed [(5'h11):(1'h0)] wire2933;
  assign y = {reg3030,
                 reg3029,
                 reg3028,
                 reg3027,
                 reg3026,
                 forvar3025,
                 forvar3024,
                 reg3023,
                 reg3022,
                 reg3021,
                 reg3020,
                 reg3019,
                 reg3018,
                 reg3017,
                 reg3016,
                 forvar3015,
                 reg3014,
                 reg3013,
                 forvar3012,
                 reg3011,
                 forvar3010,
                 reg3009,
                 reg3008,
                 reg3007,
                 wire3006,
                 reg3005,
                 reg3004,
                 reg3003,
                 wire3001,
                 wire3000,
                 reg2999,
                 reg2998,
                 reg2997,
                 reg2996,
                 forvar2995,
                 reg2994,
                 reg2993,
                 reg2992,
                 reg2991,
                 reg2990,
                 forvar2989,
                 reg2988,
                 reg2987,
                 forvar2986,
                 forvar2985,
                 reg2984,
                 reg2983,
                 forvar2982,
                 reg2981,
                 reg2980,
                 reg2979,
                 reg2978,
                 reg2977,
                 reg2976,
                 reg2975,
                 reg2974,
                 reg2973,
                 forvar2972,
                 reg2971,
                 reg2970,
                 forvar2969,
                 reg2968,
                 reg2967,
                 reg2966,
                 reg2965,
                 reg2964,
                 reg2963,
                 reg2962,
                 reg2961,
                 reg2960,
                 forvar2956,
                 reg2959,
                 reg2958,
                 reg2957,
                 reg2956,
                 reg2955,
                 reg2954,
                 reg2953,
                 reg2952,
                 forvar2951,
                 reg2950,
                 reg2949,
                 forvar2948,
                 reg2947,
                 reg2946,
                 reg2945,
                 reg2944,
                 forvar2943,
                 forvar2942,
                 reg2941,
                 reg2940,
                 forvar2939,
                 reg2938,
                 reg2937,
                 forvar2936,
                 reg2935,
                 wire2919,
                 wire53,
                 wire2921,
                 reg2923,
                 reg2924,
                 reg2925,
                 forvar2926,
                 reg2927,
                 reg2928,
                 wire2929,
                 wire2930,
                 wire2932,
                 wire2933,
                 (1'h0)};
  assign wire53 = (wire49 ?
                      $unsigned({(wire52 | wire52[(2'h2):(1'h0)]),
                          (wire49 > {wire51})}) : $signed(wire49));
  module54 modinst2920 (.wire58(wire53), .wire59(wire51), .y(wire2919), .wire55(wire52), .clk(clk), .wire57(wire50), .wire56(wire49));
  module2349 modinst2922 (wire2921, clk, wire51, wire2919, wire52, wire49);
  always
    @(posedge clk) begin
      reg2923 <= wire49;
      reg2924 = $signed("6b1vprfW5E80HBrtC0rs");
      reg2925 = $unsigned((reg2923[(4'hb):(2'h3)] == "RpwwfsrBxPig87"));
      for (forvar2926 = (1'h0); (forvar2926 < (3'h5)); forvar2926 = (forvar2926 + (1'h1)))
        begin
          reg2927 <= forvar2926[(2'h2):(2'h2)];
          reg2928 <= reg2927[(5'h15):(5'h13)];
        end
    end
  assign wire2929 = "1xUgDab8z";
  module690 modinst2931 (.clk(clk), .wire692(wire51), .y(wire2930), .wire691(reg2927), .wire694(wire2921), .wire693(wire2929));
  assign wire2932 = reg2924[(4'h8):(3'h7)];
  module1947 modinst2934 (wire2933, clk, wire51, wire2932, reg2923, wire53, wire2919);
  always
    @(posedge clk) begin
      reg2935 <= ($unsigned($signed($unsigned($signed(forvar2926)))) ?
          $signed($unsigned((reg2928 ^~ ((7'h48) ?
              reg2925 : wire2932)))) : (~&(|$signed((wire2933 ?
              wire2932 : wire2919)))));
    end
  always
    @(posedge clk) begin
      for (forvar2936 = (1'h0); (forvar2936 < (2'h3)); forvar2936 = (forvar2936 + (1'h1)))
        begin
          reg2937 <= {$unsigned(reg2925[(5'h10):(4'h9)])};
          reg2938 <= $signed((~reg2927[(4'hf):(1'h1)]));
        end
      for (forvar2939 = (1'h0); (forvar2939 < (2'h2)); forvar2939 = (forvar2939 + (1'h1)))
        begin
          reg2940 <= $unsigned(((8'hb2) != wire52));
          reg2941 <= $signed((-{$signed(wire53)}));
          for (forvar2942 = (1'h0); (forvar2942 < (2'h3)); forvar2942 = (forvar2942 + (1'h1)))
            begin
              for (forvar2943 = (1'h0); (forvar2943 < (1'h0)); forvar2943 = (forvar2943 + (1'h1)))
                begin
                  reg2944 <= forvar2939[(3'h6):(2'h3)];
                  reg2945 = (wire2919[(2'h2):(1'h0)] ?
                      {"ORWQ10TfpD",
                          ((wire51 ? "cJKN" : $signed(wire2921)) ?
                              (^wire2919[(1'h0):(1'h0)]) : {(^wire2932),
                                  $signed(wire50)})} : ($signed(({wire2933,
                                  wire2929} ?
                              wire49 : forvar2939[(4'hd):(2'h3)])) ?
                          (|"d") : ((|(reg2927 ?
                              wire49 : reg2928)) >= $signed("w"))));
                  reg2946 <= (("JlewU" - $signed("hs2GQNw88WmVlXUudz")) ?
                      reg2938 : ("K5Gzcx" && (-"U6Id6fzgEVx9EAz")));
                  reg2947 = reg2925[(4'h9):(3'h6)];
                end
              for (forvar2948 = (1'h0); (forvar2948 < (3'h5)); forvar2948 = (forvar2948 + (1'h1)))
                begin
                  reg2949 <= forvar2939;
                end
              reg2950 <= wire50;
              for (forvar2951 = (1'h0); (forvar2951 < (3'h4)); forvar2951 = (forvar2951 + (1'h1)))
                begin
                  reg2952 <= (8'hb7);
                  reg2953 = ($unsigned(((&$unsigned(reg2944)) ?
                      $signed($unsigned(reg2946)) : {(-reg2946),
                          {reg2947}})) != reg2925[(5'h11):(3'h7)]);
                end
              reg2954 <= wire2921[(4'he):(4'he)];
              reg2955 <= $signed((forvar2936 ?
                  $signed({(forvar2943 && wire2929)}) : wire2929));
            end
          if ($unsigned($unsigned(forvar2943)))
            begin
              reg2956 <= ("2YF0h4pAN6WB" ?
                  {(8'hae),
                      (+(forvar2943[(5'h12):(4'h8)] || (reg2938 ?
                          wire2929 : wire2930)))} : reg2927[(1'h0):(1'h0)]);
              reg2957 <= ({reg2947[(3'h4):(3'h4)]} > (8'haa));
              reg2958 <= "6iQc";
              reg2959 <= (-"82XYyIhqEsVPBtykk");
            end
          else
            begin
              for (forvar2956 = (1'h0); (forvar2956 < (1'h1)); forvar2956 = (forvar2956 + (1'h1)))
                begin
                  reg2957 = ((reg2938 ? reg2954 : forvar2936[(3'h5):(2'h3)]) ?
                      (+reg2938[(5'h12):(1'h1)]) : reg2959[(2'h2):(1'h0)]);
                  reg2958 <= "u4B1JmLylZvCDkS7a8FqW";
                end
              reg2959 <= ((~^forvar2948[(4'ha):(3'h7)]) << {"XXfymI1",
                  (^~($unsigned(reg2924) ?
                      $signed(forvar2942) : $unsigned(reg2954)))});
              if ({"5mbHWwUO3ZsUW7H"})
                begin
                  reg2960 <= "gfW86xv";
                  reg2961 <= $unsigned(wire2919);
                  reg2962 <= $unsigned((($unsigned(reg2927[(5'h17):(2'h2)]) ?
                      {(forvar2926 || wire2919)} : $unsigned($signed(wire52))) - $signed($unsigned($signed(forvar2951)))));
                  reg2963 = (~$signed($unsigned(reg2959)));
                end
              else
                begin
                  reg2960 <= (~$signed($unsigned($unsigned($signed(forvar2939)))));
                  reg2961 = $unsigned(wire49[(4'hd):(3'h7)]);
                  reg2962 <= $signed((^~(reg2963[(4'hd):(2'h2)] ^~ {wire2932[(2'h2):(1'h0)]})));
                  reg2963 <= ("p" >> $signed((forvar2956 * "HIGYlHPEbrRV6XLl")));
                end
              reg2964 <= (~^{forvar2939, $unsigned({(+(8'hb6))})});
              reg2965 <= $signed($signed($signed(((~|reg2958) <= (~&reg2961)))));
              reg2966 <= ((forvar2926[(2'h3):(1'h1)] ?
                  (7'h4a) : (forvar2939 && $unsigned((+reg2961)))) == $unsigned(forvar2948));
            end
        end
      reg2967 <= wire2930[(2'h2):(1'h1)];
      reg2968 <= ((reg2947[(1'h1):(1'h1)] == $unsigned(reg2946)) + reg2957[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      for (forvar2969 = (1'h0); (forvar2969 < (2'h2)); forvar2969 = (forvar2969 + (1'h1)))
        begin
          reg2970 <= wire2921[(4'ha):(4'ha)];
          reg2971 <= reg2950;
        end
      for (forvar2972 = (1'h0); (forvar2972 < (1'h0)); forvar2972 = (forvar2972 + (1'h1)))
        begin
          reg2973 = (reg2944[(4'ha):(1'h1)] == "rNZuuaMmWPBLH8oU");
          reg2974 <= (($signed((~reg2965[(2'h2):(1'h1)])) != {(+(wire49 | reg2959)),
              "hglKEoBfx4fZMUlMTmYUxGTp3"}) >> $signed(reg2968[(1'h0):(1'h0)]));
          reg2975 <= (reg2960[(1'h0):(1'h0)] <<< wire2919[(4'hf):(4'hd)]);
          reg2976 <= (wire49 ~^ ($signed((^"nM1Ny")) ~^ forvar2969));
          reg2977 <= (reg2944 >= $unsigned(reg2955[(3'h5):(3'h4)]));
          reg2978 <= "VOTUiMcuNJMIemNfdbMP08";
        end
      reg2979 <= (!forvar2951);
      reg2980 <= $unsigned({(~|$signed($unsigned(reg2959)))});
      reg2981 = reg2966[(3'h6):(3'h6)];
    end
  always
    @(posedge clk) begin
      for (forvar2982 = (1'h0); (forvar2982 < (2'h3)); forvar2982 = (forvar2982 + (1'h1)))
        begin
          reg2983 <= "LhM";
        end
      reg2984 <= reg2965[(2'h2):(2'h2)];
      for (forvar2985 = (1'h0); (forvar2985 < (1'h0)); forvar2985 = (forvar2985 + (1'h1)))
        begin
          for (forvar2986 = (1'h0); (forvar2986 < (2'h2)); forvar2986 = (forvar2986 + (1'h1)))
            begin
              reg2987 = "nVMJvqL93Iw";
              reg2988 = $unsigned((((^reg2974) | (~&(reg2980 ?
                  reg2927 : reg2957))) ^ reg2949[(3'h5):(1'h1)]));
              for (forvar2989 = (1'h0); (forvar2989 < (2'h3)); forvar2989 = (forvar2989 + (1'h1)))
                begin
                  reg2990 <= ((~&$unsigned("hzHHnC5MN8k4SholsYMa")) >>> $unsigned(reg2967));
                  reg2991 = "OFZw1sluh";
                  reg2992 <= $unsigned((((7'h41) >>> ($signed((8'ha5)) ?
                          (~^reg2987) : {reg2952})) ?
                      ("T9K2Q0AK5WOCxaJG7a07PI4J" >= $unsigned((!reg2927))) : (^$signed("HHNtszcRsdziav"))));
                end
              reg2993 = "QBggDoQ";
              reg2994 = wire2919[(1'h0):(1'h0)];
              for (forvar2995 = (1'h0); (forvar2995 < (1'h0)); forvar2995 = (forvar2995 + (1'h1)))
                begin
                  reg2996 = (((-"hWrgyBxCPA9") ?
                          $signed("1zHdGIY0Cal2VC") : "e25xvC7i8upNC5lyRf7") ?
                      $signed((^{$signed(reg2940),
                          "teZP5KT"})) : (~^$signed("O7YSbq52ab06pI3yAn4nBsI")));
                  reg2997 <= (^~($signed("o4XSIJgF8LeWW") ^ (($unsigned(reg2970) > $unsigned(reg2945)) ?
                      reg2956 : $signed((reg2960 && reg2977)))));
                  reg2998 <= (&(reg2954[(4'ha):(3'h7)] | "0RdiTfwwWGwLM9vXxa"));
                  reg2999 <= ($unsigned(("6" < ({reg2963,
                      reg2994} ^~ (8'haf)))) | ((~^(7'h44)) ?
                      ($signed((reg2958 ?
                          reg2923 : reg2962)) - $signed($signed(reg2928))) : (~reg2962[(3'h5):(2'h3)])));
                end
            end
        end
    end
  assign wire3000 = $signed($unsigned((+$unsigned({wire52}))));
  module2349 modinst3002 (wire3001, clk, wire52, reg2946, reg2976, reg2923);
  always
    @(posedge clk) begin
      reg3003 <= $signed($signed(wire50[(5'h13):(4'hf)]));
      reg3004 <= reg2956;
      reg3005 = ("VMXdlznm8r7QaaXMxdmqkp7" ? wire2929 : reg2953[(3'h6):(3'h5)]);
    end
  assign wire3006 = "8OCu7WpS";
  always
    @(posedge clk) begin
      reg3007 <= reg2924;
      reg3008 <= $unsigned(($signed((+"dmD8k")) ?
          reg2954 : {(reg2984[(2'h2):(1'h0)] >= forvar2948[(3'h7):(1'h1)])}));
      reg3009 = $unsigned(reg2953[(4'hd):(4'hc)]);
      for (forvar3010 = (1'h0); (forvar3010 < (2'h2)); forvar3010 = (forvar3010 + (1'h1)))
        begin
          reg3011 <= reg2997;
          for (forvar3012 = (1'h0); (forvar3012 < (3'h5)); forvar3012 = (forvar3012 + (1'h1)))
            begin
              reg3013 = $unsigned((("AfRYwCJsuf915dMa8" ?
                  (forvar2985[(1'h1):(1'h1)] ~^ (reg2996 ?
                      reg2952 : reg2954)) : $unsigned((~^reg2925))) - reg2944[(3'h7):(3'h4)]));
              reg3014 <= (((reg2960 ?
                  {$unsigned(reg2965),
                      $unsigned(reg2952)} : reg2975) * $signed("LpmdZ0p")) <<< forvar2926[(1'h0):(1'h0)]);
              for (forvar3015 = (1'h0); (forvar3015 < (1'h0)); forvar3015 = (forvar3015 + (1'h1)))
                begin
                  reg3016 <= reg3004[(3'h4):(1'h0)];
                  reg3017 <= (|(~&"c"));
                  reg3018 = $signed($unsigned((+reg2960)));
                  reg3019 <= (~|$signed(reg3004));
                  reg3020 <= (&$signed($signed(($signed(reg2990) ?
                      (~&wire3000) : ((8'ha2) ? forvar3010 : reg2935)))));
                  reg3021 <= "ExcXLLorHTXy8e91afkHIA";
                end
              reg3022 <= {("h4ywa6N5sFTITERHp" - reg3005[(3'h7):(2'h3)])};
            end
          reg3023 <= reg2997;
          for (forvar3024 = (1'h0); (forvar3024 < (1'h0)); forvar3024 = (forvar3024 + (1'h1)))
            begin
              for (forvar3025 = (1'h0); (forvar3025 < (1'h1)); forvar3025 = (forvar3025 + (1'h1)))
                begin
                  reg3026 <= {$unsigned("AUFo7mAmcM6")};
                end
              reg3027 <= (forvar3015 ?
                  wire53[(4'ha):(4'ha)] : $signed(((^{reg2938, forvar3010}) ?
                      {reg2949} : {$signed(wire2932), reg2941})));
            end
          reg3028 = forvar2942;
        end
      reg3029 <= reg2937;
      reg3030 <= (($signed(("" ?
          {(8'h9c), reg2987} : (~&reg2962))) & $signed(((+forvar2969) ?
          reg2962[(1'h1):(1'h0)] : reg2996[(2'h2):(1'h0)]))) || $signed(($unsigned((reg2980 + reg2980)) ?
          ($unsigned(wire53) < reg2935[(1'h0):(1'h0)]) : $unsigned(forvar3024))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module54  (y, clk, wire59, wire58, wire57, wire56, wire55);
  output wire [(32'h3c6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire59;
  input wire signed [(3'h7):(1'h0)] wire58;
  input wire [(5'h17):(1'h0)] wire57;
  input wire [(5'h10):(1'h0)] wire56;
  input wire signed [(5'h19):(1'h0)] wire55;
  reg [(5'h1a):(1'h0)] reg2918 = (1'h0);
  reg [(5'h10):(1'h0)] reg2917 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2916 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2915 = (1'h0);
  reg [(5'h15):(1'h0)] reg2914 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2913 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2912 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2911 = (1'h0);
  reg [(5'h17):(1'h0)] reg2910 = (1'h0);
  reg [(5'h16):(1'h0)] reg2909 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2908 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2907 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2906 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2905 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2904 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2903 = (1'h0);
  reg [(5'h19):(1'h0)] reg2902 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2901 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2900 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2899 = (1'h0);
  reg [(5'h18):(1'h0)] reg2898 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2897 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2896 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2895 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2894 = (1'h0);
  reg [(3'h6):(1'h0)] reg2893 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2892 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2891 = (1'h0);
  reg [(3'h6):(1'h0)] reg2890 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2889 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2888 = (1'h0);
  reg [(5'h16):(1'h0)] reg2887 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2886 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2885 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2884 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2883 = (1'h0);
  reg [(4'he):(1'h0)] reg2882 = (1'h0);
  reg [(5'h10):(1'h0)] reg2881 = (1'h0);
  reg [(5'h12):(1'h0)] reg2880 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2879 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2878 = (1'h0);
  reg [(4'he):(1'h0)] reg2877 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2876 = (1'h0);
  reg [(5'h13):(1'h0)] reg2875 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2874 = (1'h0);
  wire [(4'ha):(1'h0)] wire2872;
  wire [(5'h16):(1'h0)] wire2871;
  reg [(5'h12):(1'h0)] reg2870 = (1'h0);
  reg [(4'h9):(1'h0)] reg2869 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2868 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2867 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2866 = (1'h0);
  reg [(5'h11):(1'h0)] reg2865 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2864 = (1'h0);
  wire [(5'h18):(1'h0)] wire2863;
  wire [(5'h19):(1'h0)] wire2862;
  wire signed [(4'hc):(1'h0)] wire2860;
  wire signed [(5'h10):(1'h0)] wire60;
  assign y = {reg2918,
                 reg2917,
                 reg2916,
                 reg2915,
                 reg2914,
                 reg2913,
                 forvar2912,
                 forvar2911,
                 reg2910,
                 reg2909,
                 reg2908,
                 forvar2907,
                 reg2906,
                 reg2905,
                 reg2904,
                 reg2903,
                 reg2902,
                 reg2901,
                 reg2900,
                 forvar2899,
                 reg2898,
                 forvar2897,
                 forvar2896,
                 reg2895,
                 reg2894,
                 reg2893,
                 reg2892,
                 reg2891,
                 reg2890,
                 forvar2889,
                 reg2888,
                 reg2887,
                 forvar2886,
                 reg2885,
                 reg2884,
                 reg2883,
                 reg2882,
                 reg2881,
                 reg2880,
                 reg2879,
                 forvar2878,
                 reg2877,
                 reg2876,
                 reg2875,
                 reg2874,
                 wire2872,
                 wire2871,
                 reg2870,
                 reg2869,
                 reg2868,
                 reg2867,
                 reg2866,
                 reg2865,
                 reg2864,
                 wire2863,
                 wire2862,
                 wire2860,
                 wire60,
                 (1'h0)};
  assign wire60 = $unsigned($signed($unsigned("S6npbPoAwcwtZ")));
  module61 modinst2861 (.wire63(wire55), .wire64(wire60), .y(wire2860), .clk(clk), .wire65(wire57), .wire62(wire59));
  assign wire2862 = wire56;
  assign wire2863 = (~^{($unsigned(wire2862) ?
                            $unsigned($signed(wire2862)) : "iRi2yY0TUQpCrSF3llJON")});
  always
    @(posedge clk) begin
      reg2864 = {{(~|$signed((8'ha3))), (!(~^(7'h4e)))}};
      reg2865 <= wire56[(1'h0):(1'h0)];
      reg2866 = (~^$signed(("QwohZZv9wlc2xYXEwEhXH8q1" ?
          (^"FXd3CWK7IlbSRVnw") : "ttNNNSfVlYXGIBGi")));
    end
  always
    @(posedge clk) begin
      reg2867 <= $unsigned($signed(wire2863[(4'he):(3'h5)]));
      reg2868 <= $unsigned((8'ha9));
    end
  always
    @(posedge clk) begin
      reg2869 = (wire58[(1'h1):(1'h1)] ?
          ((^"sT") ?
              (((-reg2864) - "1yK") ?
                  {"IQt2W8wM",
                      (reg2865 ^ wire2860)} : $unsigned($unsigned(wire60))) : (({wire59,
                          wire60} ?
                      (|wire2862) : $signed((8'ha2))) ?
                  $unsigned("r") : wire59[(4'he):(4'hb)])) : (^~wire2862));
      reg2870 <= $unsigned($signed(wire58));
    end
  assign wire2871 = $signed(reg2869[(3'h7):(1'h1)]);
  module61 modinst2873 (wire2872, clk, wire60, wire2860, wire2862, reg2870);
  always
    @(posedge clk) begin
      reg2874 <= ($unsigned(((-$signed(reg2869)) >> ((~reg2870) ?
          reg2866[(4'hf):(1'h0)] : $unsigned(wire59)))) <= "TQbCYV");
      reg2875 <= $signed(((((wire58 == wire58) ?
              $signed(wire58) : "wPugCKn3mCo") < $unsigned(wire59[(4'h9):(4'h8)])) ?
          wire60[(4'h8):(3'h7)] : (reg2865 & ($signed(reg2865) ?
              {(8'hbe), (8'ha2)} : (8'hb0)))));
      reg2876 <= $signed($unsigned(wire2860));
      reg2877 <= wire2863;
      for (forvar2878 = (1'h0); (forvar2878 < (1'h1)); forvar2878 = (forvar2878 + (1'h1)))
        begin
          reg2879 <= wire56[(4'hb):(4'h8)];
          reg2880 <= $unsigned((7'h42));
          reg2881 <= ({$signed("S2"), "u73L4wJKWN"} ?
              {$unsigned((^((8'haf) ? reg2879 : reg2880))),
                  {$signed(((8'hb1) ? wire2860 : reg2864)),
                      $unsigned({reg2865, wire57})}} : "1trqP4YMwu4JNX4AR9U");
          reg2882 = ($signed($unsigned($signed(((8'ha0) || reg2880)))) << $signed(reg2870));
          reg2883 <= $signed({reg2880, wire55[(2'h3):(2'h2)]});
          reg2884 = wire56;
        end
      if ({$unsigned((~&((^~reg2874) ?
              reg2865[(1'h1):(1'h1)] : "52FgJgSqpGfF1DJ7e6UlTS"))),
          ($unsigned(reg2884[(3'h6):(2'h3)]) << (({reg2864} ?
              {(8'hb9)} : $signed(reg2875)) * wire55[(2'h3):(2'h3)]))})
        begin
          reg2885 = {(8'hb9)};
          for (forvar2886 = (1'h0); (forvar2886 < (2'h2)); forvar2886 = (forvar2886 + (1'h1)))
            begin
              reg2887 <= (reg2870[(4'ha):(4'h8)] ?
                  $signed(("3I10nuHLLYSmhKVBY6o" != reg2876)) : $signed((^~((-reg2877) << reg2865))));
            end
          reg2888 <= $signed((^(&(|(forvar2886 >>> reg2883)))));
        end
      else
        begin
          reg2885 <= "RbRxY2mSI49eUe";
          for (forvar2886 = (1'h0); (forvar2886 < (3'h4)); forvar2886 = (forvar2886 + (1'h1)))
            begin
              reg2887 <= reg2876;
              reg2888 = (~(wire59 ?
                  reg2884[(1'h0):(1'h0)] : reg2880[(3'h4):(2'h2)]));
            end
          for (forvar2889 = (1'h0); (forvar2889 < (2'h2)); forvar2889 = (forvar2889 + (1'h1)))
            begin
              reg2890 <= "mDc4LstzrcsldEGkKvwe97DQ";
              reg2891 <= $signed("cQ124dU6V4uqYfS75");
              reg2892 = (^(~&"1U5YcbYDTiBlDee"));
            end
        end
    end
  always
    @(posedge clk) begin
      reg2893 = reg2877[(2'h2):(1'h0)];
      reg2894 <= ((^~reg2888) & ($signed({$unsigned(forvar2886),
              $unsigned((8'haa))}) ?
          $unsigned("MLP4BLL5Wz18") : $unsigned(reg2891)));
      reg2895 = $signed($unsigned("n"));
      for (forvar2896 = (1'h0); (forvar2896 < (1'h0)); forvar2896 = (forvar2896 + (1'h1)))
        begin
          for (forvar2897 = (1'h0); (forvar2897 < (2'h2)); forvar2897 = (forvar2897 + (1'h1)))
            begin
              reg2898 = "ClGw7EOn9PQ7NvySpGVa";
              for (forvar2899 = (1'h0); (forvar2899 < (1'h1)); forvar2899 = (forvar2899 + (1'h1)))
                begin
                  reg2900 <= reg2880;
                  reg2901 <= "UrG9";
                  reg2902 <= ($signed($unsigned($signed($unsigned(reg2866)))) ~^ $signed(reg2864[(4'h8):(3'h5)]));
                end
            end
          reg2903 <= ($signed(reg2900) ?
              reg2880 : {(-wire2862[(2'h3):(1'h1)])});
          reg2904 = reg2902[(5'h14):(3'h6)];
        end
    end
  always
    @(posedge clk) begin
      reg2905 <= (wire2871 ? reg2890[(2'h2):(2'h2)] : reg2903);
      reg2906 <= reg2888[(5'h10):(2'h2)];
      for (forvar2907 = (1'h0); (forvar2907 < (1'h0)); forvar2907 = (forvar2907 + (1'h1)))
        begin
          reg2908 <= (8'ha5);
          reg2909 <= (+(forvar2889 >> (wire58 ?
              wire2872[(4'h8):(3'h4)] : "7ZlCZfKWqPtQRJdH")));
          reg2910 <= $unsigned((~&"mH8RJSJvEl4FNZGXK3WaQSnyd"));
          for (forvar2911 = (1'h0); (forvar2911 < (1'h1)); forvar2911 = (forvar2911 + (1'h1)))
            begin
              for (forvar2912 = (1'h0); (forvar2912 < (2'h3)); forvar2912 = (forvar2912 + (1'h1)))
                begin
                  reg2913 = $signed($unsigned("RyXgtxfoMK8BU7aWqFi4o0Htd"));
                  reg2914 <= reg2903;
                  reg2915 = (reg2876[(2'h2):(1'h1)] >> "wXnkeT");
                end
              reg2916 <= "LnyCWsQy71nxCC4aOCOXPsMA";
            end
          reg2917 <= (reg2909[(4'hc):(2'h3)] <= (^~(wire57 ?
              ((wire60 > (7'h40)) | {reg2883}) : ((forvar2896 ?
                  reg2877 : reg2910) > (wire2862 ? (7'h44) : reg2903)))));
          reg2918 = (~^(8'ha9));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module61  (y, clk, wire65, wire64, wire63, wire62);
  output wire [(32'h57a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire65;
  input wire [(4'hc):(1'h0)] wire64;
  input wire [(5'h19):(1'h0)] wire63;
  input wire signed [(5'h10):(1'h0)] wire62;
  wire signed [(4'h9):(1'h0)] wire2859;
  wire [(2'h3):(1'h0)] wire2857;
  reg [(5'h1a):(1'h0)] reg2856 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2855 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2854 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2853 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2852 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2851 = (1'h0);
  reg [(3'h4):(1'h0)] reg2850 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2849 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2848 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2847 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2846 = (1'h0);
  reg [(3'h5):(1'h0)] reg2845 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2844 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2843 = (1'h0);
  reg [(5'h19):(1'h0)] reg2842 = (1'h0);
  wire signed [(4'he):(1'h0)] wire2838;
  wire [(5'h18):(1'h0)] wire2806;
  wire [(5'h14):(1'h0)] wire2804;
  wire [(3'h4):(1'h0)] wire1936;
  reg [(5'h17):(1'h0)] reg661 = (1'h0);
  wire [(5'h16):(1'h0)] wire207;
  reg [(5'h18):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar74 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg72 = (1'h0);
  reg [(4'hc):(1'h0)] reg71 = (1'h0);
  reg [(5'h15):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar69 = (1'h0);
  reg [(5'h19):(1'h0)] reg68 = (1'h0);
  reg [(5'h1a):(1'h0)] reg67 = (1'h0);
  reg [(5'h19):(1'h0)] reg66 = (1'h0);
  reg signed [(4'he):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg210 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg211 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg212 = (1'h0);
  wire [(2'h3):(1'h0)] wire213;
  reg signed [(5'h19):(1'h0)] reg214 = (1'h0);
  reg [(5'h17):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg216 = (1'h0);
  wire [(5'h13):(1'h0)] wire659;
  wire [(5'h18):(1'h0)] wire1938;
  reg [(5'h15):(1'h0)] reg1939 = (1'h0);
  reg [(5'h15):(1'h0)] reg1940 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1941 = (1'h0);
  reg [(5'h13):(1'h0)] reg1942 = (1'h0);
  reg [(4'ha):(1'h0)] reg1943 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1944 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1945 = (1'h0);
  reg [(5'h13):(1'h0)] reg1946 = (1'h0);
  wire [(5'h19):(1'h0)] wire2802;
  reg signed [(5'h19):(1'h0)] reg2808 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2809 = (1'h0);
  reg [(5'h14):(1'h0)] reg2810 = (1'h0);
  reg [(3'h5):(1'h0)] reg2811 = (1'h0);
  reg [(4'hc):(1'h0)] reg2812 = (1'h0);
  reg [(3'h5):(1'h0)] reg2813 = (1'h0);
  wire [(5'h13):(1'h0)] wire2814;
  reg signed [(5'h11):(1'h0)] forvar2815 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2816 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2817 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2818 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2819 = (1'h0);
  reg [(3'h4):(1'h0)] reg2820 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2821 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2822 = (1'h0);
  reg [(5'h15):(1'h0)] reg2823 = (1'h0);
  reg [(5'h13):(1'h0)] forvar2824 = (1'h0);
  reg [(5'h13):(1'h0)] reg2825 = (1'h0);
  reg [(5'h12):(1'h0)] reg2826 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2827 = (1'h0);
  reg [(4'ha):(1'h0)] reg2828 = (1'h0);
  reg [(5'h13):(1'h0)] reg2829 = (1'h0);
  reg [(3'h5):(1'h0)] reg2830 = (1'h0);
  reg [(5'h19):(1'h0)] reg2831 = (1'h0);
  reg [(5'h17):(1'h0)] reg2832 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2833 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2834 = (1'h0);
  reg [(5'h13):(1'h0)] reg2835 = (1'h0);
  wire [(4'h8):(1'h0)] wire2836;
  wire [(5'h12):(1'h0)] wire2840;
  assign y = {wire2859,
                 wire2857,
                 reg2856,
                 reg2855,
                 reg2854,
                 reg2853,
                 reg2852,
                 forvar2851,
                 reg2850,
                 reg2849,
                 reg2848,
                 reg2847,
                 reg2846,
                 reg2845,
                 reg2844,
                 forvar2843,
                 reg2842,
                 wire2838,
                 wire2806,
                 wire2804,
                 wire1936,
                 reg661,
                 wire207,
                 reg75,
                 forvar74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 forvar69,
                 reg68,
                 reg67,
                 reg66,
                 reg209,
                 reg210,
                 reg211,
                 reg212,
                 wire213,
                 reg214,
                 reg215,
                 reg216,
                 wire659,
                 wire1938,
                 reg1939,
                 reg1940,
                 reg1941,
                 reg1942,
                 reg1943,
                 forvar1944,
                 reg1945,
                 reg1946,
                 wire2802,
                 reg2808,
                 forvar2809,
                 reg2810,
                 reg2811,
                 reg2812,
                 reg2813,
                 wire2814,
                 forvar2815,
                 forvar2816,
                 reg2817,
                 reg2818,
                 forvar2819,
                 reg2820,
                 reg2821,
                 reg2822,
                 reg2823,
                 forvar2824,
                 reg2825,
                 reg2826,
                 reg2827,
                 reg2828,
                 reg2829,
                 reg2830,
                 reg2831,
                 reg2832,
                 reg2833,
                 reg2834,
                 reg2835,
                 wire2836,
                 wire2840,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg66 <= $signed($unsigned($signed($unsigned((wire62 + (7'h45))))));
      reg67 <= $unsigned(wire65[(1'h0):(1'h0)]);
      reg68 <= $unsigned((~|"QR8"));
      for (forvar69 = (1'h0); (forvar69 < (1'h1)); forvar69 = (forvar69 + (1'h1)))
        begin
          reg70 = "x";
          reg71 <= (8'hb1);
          reg72 = "xouvvWgNA";
          reg73 <= {wire64[(3'h5):(2'h2)], reg72};
          for (forvar74 = (1'h0); (forvar74 < (1'h0)); forvar74 = (forvar74 + (1'h1)))
            begin
              reg75 <= "zQdhaqxmdAiDE";
            end
        end
    end
  module76 modinst208 (.wire77(forvar74), .y(wire207), .wire78(reg67), .wire79(reg70), .clk(clk), .wire81(wire63), .wire80(reg72));
  always
    @(posedge clk) begin
      reg209 <= {"8LSV2V2nuqM1V5zW", reg70[(4'he):(3'h4)]};
      reg210 <= (~|"HElaeUpKWugQxVGzeRWsg");
      reg211 <= (forvar74[(1'h0):(1'h0)] ?
          wire207[(4'hf):(4'ha)] : $signed("BLMhsgPCp7Y"));
    end
  always
    @(posedge clk) begin
      reg212 <= $unsigned({reg67, (reg75 | reg71)});
    end
  assign wire213 = (-$unsigned(((!$signed(wire62)) >= ($unsigned((8'hab)) >>> $unsigned(reg212)))));
  always
    @(posedge clk) begin
      reg214 <= "BbqREnFb";
      reg215 <= (reg73[(1'h1):(1'h0)] ^ {(^~($unsigned(wire207) > (reg73 ?
              forvar74 : forvar69)))});
      reg216 <= ($signed($unsigned("tTbhvCtttTI5")) <<< reg72);
    end
  module217 modinst660 (.wire221(reg72), .wire218(wire64), .y(wire659), .wire220(forvar69), .clk(clk), .wire222(reg75), .wire219(wire207));
  always
    @(posedge clk) begin
      reg661 = wire65;
    end
  module662 modinst1937 (.wire667(reg210), .clk(clk), .wire665(reg214), .wire666(reg68), .y(wire1936), .wire663(forvar74), .wire664(reg216));
  assign wire1938 = reg71;
  always
    @(posedge clk) begin
      reg1939 = (wire1936 == "1m7D0zEE6TGVg3IPFJCrCgmto");
      reg1940 = (^(~|(8'ha1)));
      reg1941 = (7'h4d);
      reg1942 = $unsigned((+(($signed(reg1939) ~^ (reg214 & reg210)) ?
          "4l6krw" : reg75)));
      reg1943 = $signed($signed(("NPFL" ?
          $signed((^~reg72)) : $unsigned(((7'h44) <<< reg73)))));
      for (forvar1944 = (1'h0); (forvar1944 < (2'h3)); forvar1944 = (forvar1944 + (1'h1)))
        begin
          reg1945 <= (~reg210[(1'h0):(1'h0)]);
          reg1946 <= reg71;
        end
    end
  module1947 modinst2803 (wire2802, clk, reg1945, reg661, wire207, wire65, reg67);
  module2298 modinst2805 (.wire2302(reg210), .y(wire2804), .wire2300(wire659), .wire2301(reg1945), .wire2299(reg1941), .clk(clk));
  module1953 modinst2807 (.wire1954(reg211), .wire1955(reg1940), .y(wire2806), .wire1958(reg1941), .wire1957(reg71), .wire1956(reg216), .clk(clk));
  always
    @(posedge clk) begin
      reg2808 = (~|({"9GbccO"} ? (~reg66) : $signed(wire1938[(5'h10):(1'h1)])));
      for (forvar2809 = (1'h0); (forvar2809 < (3'h4)); forvar2809 = (forvar2809 + (1'h1)))
        begin
          reg2810 = $unsigned((($signed((!reg73)) ^ reg1942) ~^ "4D"));
        end
      reg2811 <= $unsigned((+(-{wire1938, reg73})));
      reg2812 <= $unsigned((wire1938[(1'h0):(1'h0)] ?
          forvar1944[(3'h4):(2'h3)] : (~|((!(7'h4e)) ?
              "3FOsqOvqgSJGxag7" : {reg211}))));
      reg2813 <= $signed("sJlf67Ubcx1");
    end
  assign wire2814 = reg215[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar2815 = (1'h0); (forvar2815 < (2'h2)); forvar2815 = (forvar2815 + (1'h1)))
        begin
          for (forvar2816 = (1'h0); (forvar2816 < (1'h1)); forvar2816 = (forvar2816 + (1'h1)))
            begin
              reg2817 = {(~(reg2808[(5'h17):(5'h12)] ?
                      ($unsigned((8'ha3)) ?
                          $unsigned(wire659) : (!reg70)) : $unsigned(reg70[(4'h8):(3'h5)]))),
                  (|(~&reg215))};
              reg2818 <= $signed(wire213);
              for (forvar2819 = (1'h0); (forvar2819 < (3'h5)); forvar2819 = (forvar2819 + (1'h1)))
                begin
                  reg2820 <= reg2811;
                  reg2821 <= {reg209[(3'h7):(3'h6)],
                      {$unsigned(({(8'ha8)} ? $unsigned(reg214) : forvar2809)),
                          $signed(reg2808)}};
                  reg2822 <= ($signed(reg1945[(3'h6):(2'h2)]) ^~ (reg2821 ?
                      (~^"DpyUOS73dXr") : reg1942[(4'hf):(2'h2)]));
                end
              reg2823 = (^~{{("TNUK1quo8kr0Jikhwp03Y" ?
                          $signed(forvar2816) : (~(8'hb4))),
                      $signed("1AiNVC97C")},
                  {"oiYpBBZpvFzH"}});
              for (forvar2824 = (1'h0); (forvar2824 < (2'h3)); forvar2824 = (forvar2824 + (1'h1)))
                begin
                  reg2825 <= reg1942;
                  reg2826 <= ($unsigned(reg214[(4'he):(4'ha)]) ?
                      (~^reg1945) : (~(($signed(reg1942) - (wire64 ?
                          (8'haa) : reg1941)) << $unsigned((wire63 <= reg661)))));
                  reg2827 <= ($unsigned(wire62[(3'h7):(1'h1)]) ?
                      $unsigned($unsigned({(7'h42),
                          $unsigned(reg2820)})) : $signed((~^reg2811)));
                end
              reg2828 = ($signed({reg2826, "hfzm5bvp37fg7OLere"}) ?
                  $unsigned((("qKP" <= (forvar2819 ?
                      reg1941 : (8'hb7))) <= (reg2813 ?
                      ((7'h4e) - wire659) : (wire64 >> forvar2815)))) : "m");
            end
          reg2829 <= "8hTpIJx6h6rv1i";
          reg2830 <= ((~forvar2819) ?
              $unsigned($signed(wire2802[(3'h4):(2'h3)])) : reg1946[(4'ha):(4'h8)]);
          reg2831 <= (^~((^~wire63[(4'hd):(4'hd)]) ?
              $signed(((^(8'h9c)) ^ (~^(8'hac)))) : "ExcfKxf9"));
          reg2832 = (7'h48);
          reg2833 <= wire207[(4'hf):(1'h1)];
        end
      reg2834 <= reg66[(3'h6):(1'h0)];
      reg2835 <= $signed($unsigned(((-(reg2818 ? wire65 : reg211)) ?
          {reg75[(4'hd):(4'h8)]} : {(wire1936 ? reg210 : forvar1944),
              $signed(reg2823)})));
    end
  module2707 modinst2837 (.wire2709(wire2806), .wire2708(reg214), .wire2710(reg2834), .clk(clk), .wire2711(wire207), .y(wire2836), .wire2712(forvar2824));
  module1146 modinst2839 (.wire1150(reg2810), .clk(clk), .wire1147(reg66), .wire1148(reg2832), .wire1151(wire63), .wire1149(reg2818), .y(wire2838));
  module127 modinst2841 (.wire132(reg1939), .clk(clk), .y(wire2840), .wire130(reg2808), .wire129(reg66), .wire128(reg2831), .wire131(reg68));
  always
    @(posedge clk) begin
      reg2842 = wire2838[(3'h4):(1'h1)];
      for (forvar2843 = (1'h0); (forvar2843 < (3'h5)); forvar2843 = (forvar2843 + (1'h1)))
        begin
          reg2844 <= "uVSpF5UsWz20WHNJr5dLzaT";
          reg2845 = $signed(reg2844);
          reg2846 = ($signed("DGlq1un1YalXFRMempf7yh") <= "KTM8fGUwwwJ1z8RioAvHBpm");
          reg2847 <= $signed((8'hbf));
          reg2848 <= (+((~|((forvar74 ? wire1938 : reg2835) ?
                  ((7'h48) >= wire2806) : "")) ?
              (forvar69[(3'h6):(3'h4)] << ($unsigned(reg2834) ?
                  reg215[(4'hf):(4'he)] : reg2821[(5'h16):(4'hf)])) : "rFv"));
          reg2849 <= "dQ79adJBA";
        end
      reg2850 <= (wire65[(4'hb):(3'h6)] << (reg2845 >>> {(-{reg2813}),
          (reg2812 ? $unsigned(reg214) : wire2838)}));
      for (forvar2851 = (1'h0); (forvar2851 < (2'h3)); forvar2851 = (forvar2851 + (1'h1)))
        begin
          reg2852 <= (~("VfEmm70No8GQ4PZrT" ?
              ((&"C5EfF4lfZTtJ") ? reg1943 : "cGnu2scmHSm0SzI") : reg209));
          reg2853 <= $unsigned({($signed($signed(forvar2851)) ^~ reg2821[(4'hf):(1'h1)])});
          reg2854 <= {reg2831[(3'h6):(3'h4)], reg1940};
          reg2855 <= wire65[(1'h1):(1'h1)];
        end
      reg2856 <= $unsigned(wire64[(2'h2):(2'h2)]);
    end
  module881 modinst2858 (wire2857, clk, wire62, reg70, reg1946, reg2842);
  assign wire2859 = (&reg215[(3'h7):(2'h3)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1947
#( parameter param2801 = ((+(^(^~((8'h9c) ? (8'ha7) : (8'hb6))))) ? ((~((!(7'h4d)) * ((8'hbd) & (7'h41)))) ? {(((8'had) <<< (8'ha0)) ? ((8'hb6) != (8'hb3)) : ((8'hbc) ^ (8'hbb))), (((7'h40) ? (8'had) : (7'h43)) ? {(7'h4e)} : ((7'h41) ? (8'had) : (8'ha7)))} : (~|(^((8'ha3) ? (7'h4b) : (8'hb0))))) : ((-(!((8'ha3) >= (8'hb2)))) << {(^((8'hbd) ? (8'h9f) : (7'h44)))})) )
(y, clk, wire1952, wire1951, wire1950, wire1949, wire1948);
  output wire [(32'h3f6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire1952;
  input wire [(5'h15):(1'h0)] wire1951;
  input wire [(5'h15):(1'h0)] wire1950;
  input wire signed [(5'h10):(1'h0)] wire1949;
  input wire signed [(5'h1a):(1'h0)] wire1948;
  wire [(2'h2):(1'h0)] wire2800;
  reg [(4'he):(1'h0)] reg2799 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2798 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2797 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2796 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire2705;
  wire [(3'h6):(1'h0)] wire2689;
  wire [(5'h12):(1'h0)] wire2006;
  reg signed [(5'h17):(1'h0)] reg2008 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2009 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2010 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2011 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2012 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2013 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2014 = (1'h0);
  reg [(4'hc):(1'h0)] reg2015 = (1'h0);
  reg [(5'h15):(1'h0)] reg2016 = (1'h0);
  reg [(5'h15):(1'h0)] reg2017 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2018 = (1'h0);
  reg [(5'h19):(1'h0)] forvar2019 = (1'h0);
  reg [(3'h4):(1'h0)] reg2020 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2021 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2022 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2023 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2024 = (1'h0);
  reg [(5'h16):(1'h0)] reg2025 = (1'h0);
  reg [(4'h9):(1'h0)] reg2026 = (1'h0);
  reg [(4'ha):(1'h0)] reg2027 = (1'h0);
  reg [(5'h13):(1'h0)] reg2010 = (1'h0);
  reg [(5'h14):(1'h0)] reg2011 = (1'h0);
  reg [(2'h3):(1'h0)] reg2018 = (1'h0);
  reg [(4'hc):(1'h0)] reg2019 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2020 = (1'h0);
  wire [(4'hf):(1'h0)] wire2101;
  wire signed [(5'h10):(1'h0)] wire2103;
  wire signed [(3'h7):(1'h0)] wire2104;
  reg signed [(4'hc):(1'h0)] reg2105 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2106 = (1'h0);
  reg [(2'h3):(1'h0)] reg2107 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2108 = (1'h0);
  reg [(4'h9):(1'h0)] reg2109 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2110 = (1'h0);
  wire [(3'h6):(1'h0)] wire2111;
  wire signed [(5'h19):(1'h0)] wire2225;
  wire [(5'h17):(1'h0)] wire2280;
  wire signed [(5'h18):(1'h0)] wire2282;
  wire [(4'hf):(1'h0)] wire2283;
  reg signed [(4'hc):(1'h0)] forvar2284 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2285 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2286 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2287 = (1'h0);
  reg [(5'h10):(1'h0)] reg2288 = (1'h0);
  reg [(5'h19):(1'h0)] reg2289 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2290 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2291 = (1'h0);
  reg [(5'h19):(1'h0)] reg2292 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2293 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2294 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2295 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2296 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2297 = (1'h0);
  wire [(5'h13):(1'h0)] wire2347;
  wire signed [(3'h5):(1'h0)] wire2531;
  reg signed [(5'h15):(1'h0)] reg2533 = (1'h0);
  reg [(4'hb):(1'h0)] reg2534 = (1'h0);
  reg [(5'h13):(1'h0)] reg2535 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2536 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2537 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire2590;
  wire signed [(3'h6):(1'h0)] wire2794;
  assign y = {wire2800,
                 reg2799,
                 reg2798,
                 reg2797,
                 reg2796,
                 wire2705,
                 wire2689,
                 wire2006,
                 reg2008,
                 reg2009,
                 forvar2010,
                 forvar2011,
                 reg2012,
                 reg2013,
                 reg2014,
                 reg2015,
                 reg2016,
                 reg2017,
                 forvar2018,
                 forvar2019,
                 reg2020,
                 reg2021,
                 reg2022,
                 reg2023,
                 reg2024,
                 reg2025,
                 reg2026,
                 reg2027,
                 reg2010,
                 reg2011,
                 reg2018,
                 reg2019,
                 forvar2020,
                 wire2101,
                 wire2103,
                 wire2104,
                 reg2105,
                 reg2106,
                 reg2107,
                 reg2108,
                 reg2109,
                 reg2110,
                 wire2111,
                 wire2225,
                 wire2280,
                 wire2282,
                 wire2283,
                 forvar2284,
                 reg2285,
                 forvar2286,
                 forvar2287,
                 reg2288,
                 reg2289,
                 reg2290,
                 reg2291,
                 reg2292,
                 reg2293,
                 reg2294,
                 reg2295,
                 reg2296,
                 reg2297,
                 wire2347,
                 wire2531,
                 reg2533,
                 reg2534,
                 reg2535,
                 reg2536,
                 reg2537,
                 wire2590,
                 wire2794,
                 (1'h0)};
  module1953 modinst2007 (wire2006, clk, wire1949, wire1951, wire1952, wire1950, wire1948);
  always
    @(posedge clk) begin
      if (wire1949)
        begin
          reg2008 = (wire1949 ?
              "XNgV7u8dVO4fXRiITW" : $unsigned($unsigned("qtUAAARkBPXSwPZ")));
          reg2009 = wire1950[(4'hd):(4'hb)];
          for (forvar2010 = (1'h0); (forvar2010 < (1'h1)); forvar2010 = (forvar2010 + (1'h1)))
            begin
              for (forvar2011 = (1'h0); (forvar2011 < (1'h0)); forvar2011 = (forvar2011 + (1'h1)))
                begin
                  reg2012 <= (!$signed((8'had)));
                  reg2013 <= $signed((+$unsigned((8'ha4))));
                  reg2014 <= {"mqAuvDsDwia"};
                end
              reg2015 <= (reg2008[(5'h17):(3'h6)] - $unsigned("KM"));
              reg2016 <= forvar2010[(5'h10):(4'ha)];
              reg2017 <= $signed(wire2006[(3'h4):(1'h0)]);
            end
          for (forvar2018 = (1'h0); (forvar2018 < (2'h3)); forvar2018 = (forvar2018 + (1'h1)))
            begin
              for (forvar2019 = (1'h0); (forvar2019 < (2'h2)); forvar2019 = (forvar2019 + (1'h1)))
                begin
                  reg2020 <= ($unsigned("SCBi2yUaLGgRPT7Rv0yST6") << reg2013[(1'h0):(1'h0)]);
                  reg2021 <= reg2013;
                  reg2022 = "ad0pSOUn96Gxu";
                  reg2023 = (+$unsigned(forvar2011[(2'h3):(2'h2)]));
                  reg2024 = $unsigned(wire1952[(3'h6):(3'h6)]);
                end
              reg2025 <= (((((reg2015 ?
                          reg2021 : reg2009) ^ reg2021) << "rDyfIcbC29NCiXhpdUhdrh") ?
                      reg2017[(4'hd):(1'h0)] : wire2006) ?
                  $unsigned("BOme4ADuJRLSWP0vkGtCku") : ("CpPXocz5u2" ?
                      ($signed((reg2021 ?
                          wire1948 : (8'haa))) ^ wire1949[(4'h8):(1'h1)]) : (&wire1948[(3'h7):(2'h3)])));
              reg2026 <= reg2021;
              reg2027 <= ("lC" <<< reg2020);
            end
        end
      else
        begin
          reg2008 <= (forvar2018 ?
              reg2021[(1'h1):(1'h1)] : ((((reg2016 | forvar2019) ^ {reg2014}) ?
                  reg2022 : forvar2019) << (~^(|(+reg2015)))));
          reg2009 <= (|(+(~|$signed(wire1948))));
          if ((+(wire1948[(4'hd):(3'h4)] ?
              {$unsigned((reg2008 >> (8'hbb))),
                  reg2020[(1'h0):(1'h0)]} : reg2022)))
            begin
              reg2010 <= {$signed($signed({$unsigned(reg2012),
                      $signed(reg2026)}))};
              if (reg2012[(3'h5):(2'h3)])
                begin
                  reg2011 = $signed((+"JyUDR"));
                  reg2012 <= wire2006;
                  reg2013 <= $unsigned($signed(reg2013));
                  reg2014 = forvar2010;
                  reg2015 <= (wire1948[(5'h18):(1'h0)] ?
                      "YaDdT0vsIyAW18pSxmuGrVTdD" : reg2026[(1'h1):(1'h1)]);
                end
              else
                begin
                  reg2011 = ("VzeF" & reg2023);
                  reg2012 <= {reg2008, (8'hab)};
                  reg2013 <= (($signed(wire1950[(4'ha):(4'h8)]) ?
                          {reg2013[(1'h1):(1'h1)]} : $signed("O6QAWp3ImosuRbrFRSONNWF")) ?
                      (forvar2018 ?
                          (({reg2009} & $unsigned(reg2017)) ?
                              reg2015 : forvar2018[(1'h1):(1'h0)]) : (-{(reg2009 << wire1951),
                              (wire1949 << reg2017)})) : (~($signed((forvar2018 ?
                              reg2012 : reg2008)) ?
                          $signed(wire1948[(1'h1):(1'h0)]) : forvar2019)));
                  reg2014 <= reg2021[(3'h7):(3'h7)];
                end
              if ($unsigned((wire1948 <= forvar2019)))
                begin
                  reg2016 <= $unsigned(reg2009[(4'ha):(1'h1)]);
                  reg2017 <= $unsigned("nGTwX8XYPywEHzy1bF0p");
                  reg2018 <= $signed(($unsigned($unsigned("CfesgHn8MgA")) ?
                      ((|reg2023) ?
                          ($signed(reg2024) || (forvar2018 && forvar2019)) : $signed(forvar2019)) : (-"")));
                end
              else
                begin
                  reg2016 <= "9CTKLQO6JP";
                  reg2017 <= (&$signed(($unsigned((|(8'hae))) | $unsigned(wire1951))));
                  reg2018 <= (reg2012[(3'h4):(3'h4)] ~^ "O");
                end
              reg2019 = (reg2014[(1'h0):(1'h0)] ?
                  $signed({(~(!(7'h42)))}) : $unsigned("QrSWnqys5TMe"));
              for (forvar2020 = (1'h0); (forvar2020 < (1'h1)); forvar2020 = (forvar2020 + (1'h1)))
                begin
                  reg2021 <= forvar2011[(3'h4):(2'h3)];
                  reg2022 <= forvar2011[(4'hd):(3'h6)];
                  reg2023 <= (($unsigned("BAoYsyLEu5gFChAg") ?
                      "3MFNfvxFJUHHxy" : {reg2008}) << ({"0FHW2ZOtW28n3"} ?
                      (7'h4d) : $unsigned(reg2014)));
                  reg2024 = $unsigned(reg2017[(2'h3):(2'h3)]);
                  reg2025 = forvar2019;
                  reg2026 = "tZJXTTWq2Hk1caTzKBbcKg";
                end
              reg2027 <= $signed(reg2021);
            end
          else
            begin
              reg2010 <= ($unsigned($unsigned(((&reg2013) & (reg2021 ?
                  (7'h44) : (7'h43))))) < reg2011);
              for (forvar2011 = (1'h0); (forvar2011 < (1'h1)); forvar2011 = (forvar2011 + (1'h1)))
                begin
                  reg2012 <= reg2015;
                  reg2013 = forvar2010[(5'h11):(4'he)];
                end
            end
        end
    end
  module2028 modinst2102 (wire2101, clk, reg2009, reg2026, reg2017, reg2016);
  assign wire2103 = forvar2018[(1'h1):(1'h1)];
  assign wire2104 = ((reg2009 ^ ((forvar2018[(1'h0):(1'h0)] == (reg2016 ~^ wire1950)) & $unsigned((reg2013 << (8'hb2))))) == forvar2018);
  always
    @(posedge clk) begin
      reg2105 = (~&$unsigned($unsigned(reg2011)));
      reg2106 <= $signed((~|(reg2019 ?
          $unsigned((reg2020 ? (8'ha5) : (7'h43))) : reg2024[(2'h2):(1'h0)])));
      reg2107 <= ((^{({forvar2011, (8'hb1)} ?
              reg2013 : reg2016)}) >>> reg2023[(3'h7):(3'h4)]);
      reg2108 = (8'ha0);
      reg2109 <= reg2106[(5'h15):(5'h14)];
      reg2110 <= (|$signed((~|$unsigned($signed(wire1950)))));
    end
  assign wire2111 = (((reg2015 >> reg2018[(1'h0):(1'h0)]) ?
                            "rZsmWMGylLum9UadovefHwn3y" : ($signed(reg2017[(4'hd):(2'h3)]) ^ $unsigned((~&wire1951)))) ?
                        $unsigned(((-"xfEDPsp9zSkDip233pMlHXMp") ?
                            "" : wire1948)) : $signed(reg2018));
  module2112 modinst2226 (.y(wire2225), .wire2115(wire1951), .wire2116(reg2015), .wire2113(reg2110), .clk(clk), .wire2114(forvar2011));
  module2227 modinst2281 (.wire2228(reg2015), .wire2230(wire2103), .wire2231(forvar2010), .wire2229(wire1948), .clk(clk), .y(wire2280));
  assign wire2282 = ((~^$signed((^~(forvar2019 <= wire1951)))) - forvar2011[(1'h1):(1'h1)]);
  assign wire2283 = reg2015[(4'hc):(3'h4)];
  always
    @(posedge clk) begin
      for (forvar2284 = (1'h0); (forvar2284 < (1'h1)); forvar2284 = (forvar2284 + (1'h1)))
        begin
          reg2285 <= $signed(((~|((reg2027 | reg2017) ?
              $unsigned(wire2103) : {reg2024})) ^ ({$signed((8'ha7))} != ($unsigned(reg2027) ?
              (reg2017 >= reg2015) : $signed(reg2017)))));
          for (forvar2286 = (1'h0); (forvar2286 < (1'h1)); forvar2286 = (forvar2286 + (1'h1)))
            begin
              for (forvar2287 = (1'h0); (forvar2287 < (2'h3)); forvar2287 = (forvar2287 + (1'h1)))
                begin
                  reg2288 <= wire1948[(5'h10):(5'h10)];
                  reg2289 = (~{{(|(reg2008 ? (7'h43) : wire1950)),
                          $signed(wire2283[(2'h3):(1'h0)])}});
                  reg2290 <= ("JONxaHatvOsNSkZMfSGcd9" && $signed(((~|(!(8'hac))) ?
                      ($signed(wire2006) ?
                          (wire1951 ? (8'hba) : reg2289) : (reg2107 ?
                              forvar2284 : reg2015)) : (forvar2011 ?
                          ((8'h9f) ?
                              forvar2011 : (8'h9c)) : $signed(reg2106)))));
                  reg2291 <= $signed("W7DvEiDbnZq1E");
                  reg2292 = wire1952[(2'h2):(1'h0)];
                  reg2293 <= (($signed("TTM1a71GXCTOx") ?
                          ("oRsk50B" ?
                              ((-(8'hbe)) + forvar2286) : "2e") : $signed(reg2014)) ?
                      (($signed(((8'ha9) ?
                              reg2012 : wire2103)) * {forvar2011}) ?
                          $unsigned({(reg2107 < reg2105)}) : ($unsigned(reg2108) ?
                              $unsigned({reg2289}) : $signed(reg2105[(3'h5):(3'h4)]))) : reg2290);
                end
              reg2294 <= ((~|(reg2292[(4'hb):(3'h7)] ?
                  (^reg2024) : $signed((reg2019 ?
                      reg2021 : reg2011)))) && $signed($unsigned((reg2027[(4'h8):(3'h5)] ?
                  $unsigned(forvar2019) : reg2026[(2'h3):(2'h2)]))));
              reg2295 <= "4fJSG46e3Y43G";
              reg2296 <= reg2292;
            end
          reg2297 = ((7'h49) >= wire2104[(1'h0):(1'h0)]);
        end
    end
  module2298 modinst2348 (wire2347, clk, wire2283, forvar2010, reg2297, wire2282);
  module2349 modinst2532 (wire2531, clk, reg2297, reg2288, reg2289, reg2010);
  always
    @(posedge clk) begin
      reg2533 <= ($unsigned(($unsigned((reg2296 ? reg2107 : (8'h9e))) ?
              $unsigned(forvar2018) : $unsigned("03tuPsYSVBBU6Bc72uByvF"))) ?
          (~|$signed(forvar2019)) : (~^$signed($unsigned((reg2290 >>> reg2292)))));
      reg2534 <= $unsigned(reg2021[(4'hb):(3'h4)]);
      reg2535 <= {(+reg2009)};
      reg2536 <= $signed($unsigned((wire2531 <= ({reg2295, reg2290} ?
          (~^reg2020) : $signed(reg2294)))));
      reg2537 <= ({(($unsigned(wire1952) + {wire2282, wire2111}) ?
              reg2535[(4'hd):(3'h6)] : (~^(reg2289 ?
                  (8'hb0) : reg2108)))} != ({""} >>> reg2294[(1'h0):(1'h0)]));
    end
  module2538 modinst2591 (.y(wire2590), .wire2541(forvar2284), .wire2540(wire2101), .wire2539(reg2011), .wire2542(wire1951), .wire2543(forvar2011), .clk(clk));
  module2592 modinst2690 (.wire2596(reg2019), .wire2595(wire2225), .y(wire2689), .clk(clk), .wire2594(wire2280), .wire2593(wire2101));
  module2691 modinst2706 (.wire2693(wire2006), .wire2692(reg2012), .wire2696(reg2014), .y(wire2705), .clk(clk), .wire2694(wire2590), .wire2695(reg2537));
  module2707 modinst2795 (.wire2712(reg2106), .wire2709(reg2025), .clk(clk), .wire2708(forvar2019), .y(wire2794), .wire2711(reg2296), .wire2710(wire2225));
  always
    @(posedge clk) begin
      reg2796 <= reg2106;
    end
  always
    @(posedge clk) begin
      reg2797 = ($signed((((|reg2110) ?
          (reg2008 ?
              wire2282 : wire2111) : (reg2012 >= (8'haa))) << forvar2284)) + $signed((reg2018[(1'h1):(1'h1)] ?
          $unsigned("ZozsoJnVfW9Rx5LTCzIxH9") : reg2535[(4'he):(4'h8)])));
      reg2798 <= $signed((($unsigned((forvar2010 ? reg2105 : (8'hbd))) ?
          "4ZDzXDn" : reg2285[(2'h2):(1'h1)]) ^~ reg2107));
      reg2799 <= ((+(~|(reg2017 | ((8'ha9) ?
          reg2534 : (7'h42))))) >> ($unsigned($signed($unsigned(reg2008))) ^ (~^{{(8'haf)},
          $signed(reg2797)})));
    end
  assign wire2800 = reg2294;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module662
#( parameter param1934 = (|(!(!(((8'ha9) <<< (7'h4d)) ? {(8'ha3)} : ((8'hab) ? (7'h46) : (7'h44))))))
, parameter param1935 = (param1934 >= (&(((^param1934) < {param1934}) ? ((param1934 ? (8'hbd) : (8'h9e)) ^~ (param1934 ? param1934 : param1934)) : {(param1934 + param1934)}))) )
(y, clk, wire663, wire664, wire665, wire666, wire667);
  output wire [(32'h9d8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire663;
  input wire [(5'h13):(1'h0)] wire664;
  input wire [(5'h18):(1'h0)] wire665;
  input wire signed [(4'hb):(1'h0)] wire666;
  input wire [(5'h14):(1'h0)] wire667;
  wire [(4'hb):(1'h0)] wire1932;
  reg signed [(5'h10):(1'h0)] reg1752 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1751 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1750 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1744 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1742 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1736 = (1'h0);
  reg [(5'h18):(1'h0)] reg1745 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1749 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1748 = (1'h0);
  reg [(4'hf):(1'h0)] reg1747 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1746 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1745 = (1'h0);
  reg [(5'h14):(1'h0)] reg1744 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1743 = (1'h0);
  reg [(5'h12):(1'h0)] reg1742 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1741 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1740 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1739 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1738 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1737 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1736 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1735 = (1'h0);
  reg [(5'h17):(1'h0)] reg1734 = (1'h0);
  reg [(5'h12):(1'h0)] reg1733 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1732 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1731 = (1'h0);
  reg [(5'h11):(1'h0)] reg1730 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1729 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1728 = (1'h0);
  reg [(3'h4):(1'h0)] reg1727 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1700 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1726 = (1'h0);
  reg [(4'hd):(1'h0)] reg1725 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1724 = (1'h0);
  reg [(4'hf):(1'h0)] reg1723 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1722 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1721 = (1'h0);
  reg [(3'h6):(1'h0)] reg1720 = (1'h0);
  reg [(4'h9):(1'h0)] reg1719 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1718 = (1'h0);
  reg [(3'h7):(1'h0)] reg1717 = (1'h0);
  reg [(5'h11):(1'h0)] reg1716 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1715 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1714 = (1'h0);
  reg [(4'hb):(1'h0)] reg1713 = (1'h0);
  reg [(5'h17):(1'h0)] reg1712 = (1'h0);
  reg [(4'hb):(1'h0)] reg1711 = (1'h0);
  reg [(5'h19):(1'h0)] reg1710 = (1'h0);
  reg [(5'h13):(1'h0)] reg1709 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1708 = (1'h0);
  reg [(4'hf):(1'h0)] reg1707 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1706 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1705 = (1'h0);
  reg [(5'h18):(1'h0)] reg1704 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1703 = (1'h0);
  reg [(3'h7):(1'h0)] reg1702 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1701 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1700 = (1'h0);
  reg [(5'h19):(1'h0)] reg1699 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1698 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1697 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1696 = (1'h0);
  reg [(4'ha):(1'h0)] reg1695 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1694 = (1'h0);
  reg [(4'h8):(1'h0)] reg1693 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1692 = (1'h0);
  reg [(4'hf):(1'h0)] reg1691 = (1'h0);
  reg [(5'h18):(1'h0)] reg1690 = (1'h0);
  reg [(5'h14):(1'h0)] reg1689 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1688 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1687 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1686 = (1'h0);
  reg [(5'h18):(1'h0)] reg1685 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1684 = (1'h0);
  reg [(5'h17):(1'h0)] reg1683 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1682 = (1'h0);
  reg [(4'h9):(1'h0)] reg1681 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1680 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1679 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1678 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1677 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1676 = (1'h0);
  reg [(5'h14):(1'h0)] reg1675 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1674 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1673 = (1'h0);
  reg [(4'h9):(1'h0)] reg1672 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1671 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1670 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1669 = (1'h0);
  reg [(4'hf):(1'h0)] reg1668 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1667 = (1'h0);
  wire [(4'hb):(1'h0)] wire1666;
  wire [(5'h11):(1'h0)] wire1372;
  wire [(5'h15):(1'h0)] wire668;
  wire [(5'h18):(1'h0)] wire669;
  reg signed [(5'h12):(1'h0)] forvar670 = (1'h0);
  reg [(5'h17):(1'h0)] forvar671 = (1'h0);
  reg [(5'h1a):(1'h0)] reg672 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg673 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg674 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg675 = (1'h0);
  reg [(5'h13):(1'h0)] reg676 = (1'h0);
  reg [(5'h18):(1'h0)] reg677 = (1'h0);
  reg signed [(4'he):(1'h0)] reg678 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg679 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg680 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg681 = (1'h0);
  reg [(5'h17):(1'h0)] reg682 = (1'h0);
  reg [(4'he):(1'h0)] reg683 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg684 = (1'h0);
  reg [(5'h16):(1'h0)] reg685 = (1'h0);
  reg [(4'hf):(1'h0)] reg686 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg687 = (1'h0);
  reg [(5'h17):(1'h0)] reg688 = (1'h0);
  wire [(4'he):(1'h0)] wire689;
  wire [(5'h12):(1'h0)] wire755;
  wire [(3'h6):(1'h0)] wire868;
  reg signed [(5'h15):(1'h0)] reg870 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar871 = (1'h0);
  reg [(5'h17):(1'h0)] reg872 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar873 = (1'h0);
  reg [(3'h7):(1'h0)] reg874 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg875 = (1'h0);
  reg [(5'h15):(1'h0)] reg876 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg877 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar878 = (1'h0);
  reg [(4'hf):(1'h0)] reg879 = (1'h0);
  reg [(5'h19):(1'h0)] reg880 = (1'h0);
  wire [(5'h11):(1'h0)] wire943;
  reg signed [(5'h17):(1'h0)] reg945 = (1'h0);
  reg [(5'h19):(1'h0)] reg946 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar947 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar948 = (1'h0);
  reg [(5'h18):(1'h0)] reg949 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg950 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg951 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg952 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg953 = (1'h0);
  reg [(4'h8):(1'h0)] reg954 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar955 = (1'h0);
  reg [(4'hc):(1'h0)] reg956 = (1'h0);
  wire signed [(4'he):(1'h0)] wire1144;
  reg signed [(4'hc):(1'h0)] reg1374 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1375 = (1'h0);
  reg [(5'h14):(1'h0)] reg1376 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1377 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1378 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1379 = (1'h0);
  reg [(4'hc):(1'h0)] reg1380 = (1'h0);
  reg [(4'h9):(1'h0)] reg1381 = (1'h0);
  reg [(5'h10):(1'h0)] reg1382 = (1'h0);
  wire [(4'hd):(1'h0)] wire1443;
  wire signed [(4'hd):(1'h0)] wire1445;
  wire signed [(4'ha):(1'h0)] wire1550;
  wire [(3'h6):(1'h0)] wire1552;
  wire [(3'h6):(1'h0)] wire1553;
  wire [(5'h1a):(1'h0)] wire1664;
  assign y = {wire1932,
                 reg1752,
                 reg1751,
                 reg1750,
                 forvar1744,
                 forvar1742,
                 reg1736,
                 reg1745,
                 reg1749,
                 reg1748,
                 reg1747,
                 reg1746,
                 forvar1745,
                 reg1744,
                 reg1743,
                 reg1742,
                 reg1741,
                 reg1740,
                 reg1739,
                 reg1738,
                 reg1737,
                 forvar1736,
                 forvar1735,
                 reg1734,
                 reg1733,
                 reg1732,
                 forvar1731,
                 reg1730,
                 reg1729,
                 forvar1728,
                 reg1727,
                 reg1700,
                 reg1726,
                 reg1725,
                 reg1724,
                 reg1723,
                 reg1722,
                 reg1721,
                 reg1720,
                 reg1719,
                 reg1718,
                 reg1717,
                 reg1716,
                 forvar1715,
                 forvar1714,
                 reg1713,
                 reg1712,
                 reg1711,
                 reg1710,
                 reg1709,
                 reg1708,
                 reg1707,
                 reg1706,
                 forvar1705,
                 reg1704,
                 forvar1703,
                 reg1702,
                 reg1701,
                 forvar1700,
                 reg1699,
                 reg1698,
                 reg1697,
                 reg1696,
                 reg1695,
                 reg1694,
                 reg1693,
                 forvar1692,
                 reg1691,
                 reg1690,
                 reg1689,
                 reg1688,
                 forvar1687,
                 forvar1686,
                 reg1685,
                 forvar1684,
                 reg1683,
                 reg1682,
                 reg1681,
                 reg1680,
                 forvar1679,
                 reg1678,
                 reg1677,
                 reg1676,
                 reg1675,
                 reg1674,
                 reg1673,
                 reg1672,
                 reg1671,
                 reg1670,
                 reg1669,
                 reg1668,
                 forvar1667,
                 wire1666,
                 wire1372,
                 wire668,
                 wire669,
                 forvar670,
                 forvar671,
                 reg672,
                 reg673,
                 reg674,
                 reg675,
                 reg676,
                 reg677,
                 reg678,
                 reg679,
                 reg680,
                 reg681,
                 reg682,
                 reg683,
                 reg684,
                 reg685,
                 reg686,
                 reg687,
                 reg688,
                 wire689,
                 wire755,
                 wire868,
                 reg870,
                 forvar871,
                 reg872,
                 forvar873,
                 reg874,
                 reg875,
                 reg876,
                 reg877,
                 forvar878,
                 reg879,
                 reg880,
                 wire943,
                 reg945,
                 reg946,
                 forvar947,
                 forvar948,
                 reg949,
                 reg950,
                 reg951,
                 reg952,
                 reg953,
                 reg954,
                 forvar955,
                 reg956,
                 wire1144,
                 reg1374,
                 reg1375,
                 reg1376,
                 forvar1377,
                 forvar1378,
                 reg1379,
                 reg1380,
                 reg1381,
                 reg1382,
                 wire1443,
                 wire1445,
                 wire1550,
                 wire1552,
                 wire1553,
                 wire1664,
                 (1'h0)};
  assign wire668 = "J657vaVpedANV";
  assign wire669 = ((~|"o7HEMdKMNV8iphc4Awp") ?
                       "yccVU4f1" : (^~wire663[(1'h1):(1'h1)]));
  always
    @(posedge clk) begin
      for (forvar670 = (1'h0); (forvar670 < (2'h2)); forvar670 = (forvar670 + (1'h1)))
        begin
          for (forvar671 = (1'h0); (forvar671 < (1'h0)); forvar671 = (forvar671 + (1'h1)))
            begin
              reg672 <= (^~$unsigned($signed(wire663[(4'hc):(4'ha)])));
              reg673 <= (wire665[(3'h5):(1'h1)] ?
                  "cTHIfyx6ztPICbtTp5" : $unsigned((|$signed($signed(forvar671)))));
              reg674 = $signed(reg672);
              reg675 <= "xAvT";
              reg676 = wire669;
            end
          reg677 <= ((+$unsigned(($unsigned(wire667) == ((7'h45) ?
              (8'h9f) : reg676)))) << "KK2TfiXQ2EpryHqZdmwtcLC52");
          reg678 = wire666[(4'h9):(3'h4)];
        end
      reg679 = "YCfXpJruV4PXiFUfQVToiKmB";
      reg680 <= {($signed($signed((^reg677))) ?
              $signed($unsigned({(8'hb4)})) : reg673),
          forvar671[(4'hc):(1'h0)]};
      reg681 <= "nY9QQeopK1yYe";
      reg682 <= ((7'h4e) ^~ (wire663 | (((~^wire664) ?
              ((7'h42) && forvar670) : reg679[(1'h0):(1'h0)]) ?
          $signed($unsigned(reg675)) : ((reg676 >>> wire664) ^~ $unsigned((8'ha2))))));
      reg683 <= (~^({($unsigned(reg681) != (wire666 + wire667))} == reg674[(4'hd):(3'h4)]));
    end
  always
    @(posedge clk) begin
      reg684 <= {{$signed(("7" ? $unsigned(reg678) : reg675)),
              $signed((!reg681))},
          (8'hba)};
      reg685 <= ((+(~^reg675[(2'h2):(1'h0)])) ?
          wire664[(3'h6):(3'h4)] : reg683);
      reg686 <= reg675;
      reg687 <= (($unsigned($signed((7'h4a))) < $unsigned($unsigned("zOSWzFJHU9Rm"))) ?
          ($signed($signed(reg675[(1'h0):(1'h0)])) ?
              ($unsigned(reg673[(4'ha):(4'h9)]) ?
                  ((wire667 < reg680) ?
                      wire665[(2'h2):(1'h1)] : reg679[(5'h14):(5'h14)]) : reg674[(4'hd):(3'h7)]) : (~&(~{reg679}))) : $signed((7'h41)));
      reg688 <= (7'h47);
    end
  assign wire689 = reg684[(3'h7):(3'h5)];
  module690 modinst756 (wire755, clk, reg685, wire666, wire665, wire668);
  module757 modinst869 (.wire759(wire664), .y(wire868), .wire758(wire689), .wire760(reg682), .wire761(reg686), .clk(clk));
  always
    @(posedge clk) begin
      reg870 <= $unsigned(reg675[(1'h1):(1'h1)]);
      for (forvar871 = (1'h0); (forvar871 < (2'h2)); forvar871 = (forvar871 + (1'h1)))
        begin
          reg872 <= $unsigned((reg676 ? (8'ha8) : forvar670[(4'hf):(1'h0)]));
          for (forvar873 = (1'h0); (forvar873 < (2'h3)); forvar873 = (forvar873 + (1'h1)))
            begin
              reg874 = $unsigned((8'hbc));
              reg875 <= (reg686[(1'h1):(1'h0)] | {(((8'hb4) ?
                          $unsigned(reg675) : $unsigned(forvar873)) ?
                      ("pgp65Qfv4SbNZX1aAV7alXBWS" ?
                          (forvar671 | reg685) : reg872[(1'h1):(1'h1)]) : wire868),
                  "9JFXG9W21g480DEGis"});
              reg876 = {(reg688 && reg674),
                  $unsigned(($signed((reg686 < reg682)) | ("M7rbMt" ^ (wire868 || reg874))))};
              reg877 <= $unsigned({"S3c6UMBsl3PFoLv", (8'hb3)});
              for (forvar878 = (1'h0); (forvar878 < (1'h1)); forvar878 = (forvar878 + (1'h1)))
                begin
                  reg879 <= (~|wire665);
                end
              reg880 <= reg686[(4'hc):(4'h8)];
            end
        end
    end
  module881 modinst944 (.wire882(reg677), .clk(clk), .wire884(reg876), .y(wire943), .wire885(wire667), .wire883(reg676));
  always
    @(posedge clk) begin
      reg945 <= (~&"");
      reg946 <= (reg874 > wire667);
      for (forvar947 = (1'h0); (forvar947 < (1'h0)); forvar947 = (forvar947 + (1'h1)))
        begin
          for (forvar948 = (1'h0); (forvar948 < (1'h1)); forvar948 = (forvar948 + (1'h1)))
            begin
              if ((reg880 ?
                  (-$signed((~^$signed((8'hb7))))) : ((((reg945 == reg872) ?
                          $unsigned(reg673) : "2TPdY8CRA3vaJ2LTChJ12") ^~ forvar948) ?
                      (+(((8'haf) ? wire668 : reg688) ?
                          ((8'hae) - reg876) : (^~reg946))) : $unsigned(((forvar947 >>> reg683) & (wire943 << reg685))))))
                begin
                  reg949 <= $signed((+$unsigned(reg681)));
                  reg950 = $signed((~wire868));
                  reg951 <= "mUPgmzMgsLM0LbdTYfmF";
                  reg952 <= $unsigned(("eh" ?
                      (reg684 + $signed((wire755 + reg874))) : $unsigned("doPc3WlYmYG7pR70EnC2CK")));
                end
              else
                begin
                  reg949 <= ((8'hba) ~^ reg672);
                  reg950 <= (~reg870[(4'hf):(3'h7)]);
                end
            end
        end
      reg953 <= "wTF4dvvhWJwHkJCSoIi";
      reg954 <= reg874;
      for (forvar955 = (1'h0); (forvar955 < (3'h4)); forvar955 = (forvar955 + (1'h1)))
        begin
          reg956 <= reg683[(4'hc):(2'h3)];
        end
    end
  module957 modinst1145 (wire1144, clk, reg681, forvar671, reg688, reg870, reg953);
  module1146 modinst1373 (wire1372, clk, reg880, wire668, forvar878, reg674, reg877);
  always
    @(posedge clk) begin
      reg1374 <= $unsigned(reg949[(4'hc):(4'ha)]);
      reg1375 <= reg877[(4'h9):(4'h9)];
      reg1376 <= "x";
      for (forvar1377 = (1'h0); (forvar1377 < (3'h4)); forvar1377 = (forvar1377 + (1'h1)))
        begin
          for (forvar1378 = (1'h0); (forvar1378 < (3'h5)); forvar1378 = (forvar1378 + (1'h1)))
            begin
              reg1379 <= $signed((forvar955 ?
                  (((^~(8'ha5)) ?
                      reg949 : reg688) ^ reg879[(3'h6):(2'h2)]) : ("DX13Z76G0kl637" == ((7'h47) != reg874[(3'h4):(1'h1)]))));
              reg1380 <= reg684;
              reg1381 <= (^~forvar1378);
            end
          reg1382 <= reg673[(4'h8):(3'h4)];
        end
    end
  module1383 modinst1444 (.wire1384(wire755), .wire1385(reg688), .clk(clk), .wire1386(reg870), .wire1387(reg683), .y(wire1443));
  assign wire1445 = "uSvoXu0uSEZRT";
  module1446 modinst1551 (wire1550, clk, reg1376, forvar955, reg951, reg687);
  assign wire1552 = $unsigned($unsigned($signed({$unsigned(reg677)})));
  assign wire1553 = (^"GGu");
  module1554 modinst1665 (wire1664, clk, wire1443, reg675, wire1372, reg678, wire663);
  assign wire1666 = wire1443;
  always
    @(posedge clk) begin
      for (forvar1667 = (1'h0); (forvar1667 < (1'h1)); forvar1667 = (forvar1667 + (1'h1)))
        begin
          reg1668 <= $unsigned((~(&(7'h4a))));
          reg1669 <= $signed(($signed($unsigned("FWvhmkBr5w4y")) ?
              (&{(~wire943),
                  (+wire1144)}) : $signed($signed("kdoLygKrkHOlH"))));
          reg1670 = (8'haa);
          reg1671 = {reg682,
              {(("1pNiA" * "8zYGf") ?
                      $unsigned({reg1670}) : $unsigned((forvar1378 ?
                          forvar671 : reg872)))}};
          reg1672 <= "Lkf";
          reg1673 <= $signed((((~(forvar670 && (8'hb1))) ^~ ($unsigned((8'ha5)) ?
                  reg1381 : "s")) ?
              (+reg673[(4'hb):(1'h1)]) : reg949[(4'hc):(2'h2)]));
        end
      reg1674 <= "q61PzNLbkNuuWN4hTSVxDH8";
      reg1675 <= reg672[(3'h5):(1'h1)];
      reg1676 <= $signed(($signed({$unsigned(wire666), (reg953 < wire868)}) ?
          (^$unsigned((reg675 ? forvar671 : reg1675))) : ((8'hbc) < (((7'h40) ?
              wire1445 : forvar871) | (~&wire665)))));
      reg1677 = (((|$unsigned($unsigned(reg875))) > (~reg952[(5'h11):(4'ha)])) & (|$signed(reg674)));
      reg1678 = ($signed("f7iTzqq35z4xd17Vl") || {wire868, forvar955});
    end
  always
    @(posedge clk) begin
      for (forvar1679 = (1'h0); (forvar1679 < (1'h1)); forvar1679 = (forvar1679 + (1'h1)))
        begin
          reg1680 <= (!$unsigned($unsigned((forvar871 << (^reg1375)))));
          reg1681 <= {($unsigned((+(~|wire1144))) >= $unsigned($signed(reg945[(1'h0):(1'h0)])))};
          reg1682 <= ((reg682 ^ ((forvar1667[(3'h7):(3'h5)] ?
                      "" : $unsigned(reg1675)) ?
                  ((^~(8'h9c)) - ((7'h4e) >>> forvar1377)) : (reg870[(4'h9):(3'h4)] ?
                      (reg1381 + reg872) : {forvar873, reg1678}))) ?
              $signed($signed(reg1673[(5'h15):(2'h2)])) : (reg673[(3'h7):(3'h7)] ?
                  forvar1378[(5'h16):(4'hd)] : wire663[(4'hb):(3'h6)]));
          reg1683 <= (wire1666[(3'h7):(1'h0)] | ($unsigned($unsigned($unsigned(wire868))) < {reg682}));
        end
    end
  always
    @(posedge clk) begin
      for (forvar1684 = (1'h0); (forvar1684 < (2'h2)); forvar1684 = (forvar1684 + (1'h1)))
        begin
          reg1685 <= "T1BVB9GiMR9dklHsw";
          for (forvar1686 = (1'h0); (forvar1686 < (1'h1)); forvar1686 = (forvar1686 + (1'h1)))
            begin
              for (forvar1687 = (1'h0); (forvar1687 < (1'h1)); forvar1687 = (forvar1687 + (1'h1)))
                begin
                  reg1688 <= (wire1372[(1'h1):(1'h1)] ?
                      $signed({$unsigned(reg688[(4'hc):(4'hb)]),
                          forvar1684[(2'h2):(1'h1)]}) : reg683);
                  reg1689 <= (~forvar1687);
                  reg1690 <= $unsigned(reg880);
                end
            end
          reg1691 <= reg1380[(3'h7):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar1692 = (1'h0); (forvar1692 < (2'h3)); forvar1692 = (forvar1692 + (1'h1)))
        begin
          reg1693 <= reg678;
          reg1694 <= $unsigned("crs2XS");
          reg1695 <= reg874[(2'h2):(2'h2)];
          reg1696 <= "8bls8k8BE";
          reg1697 <= (^reg870[(1'h1):(1'h1)]);
          reg1698 <= (reg687 ?
              (^~$unsigned($unsigned(((7'h48) ? reg874 : (7'h44))))) : (8'ha5));
        end
      if (((+($signed($signed(reg950)) ?
          reg877[(4'h9):(3'h5)] : $signed((wire1553 == reg952)))) * wire868))
        begin
          reg1699 <= "10UYqSxHyNUIaQKli9wQBpBp";
          for (forvar1700 = (1'h0); (forvar1700 < (1'h1)); forvar1700 = (forvar1700 + (1'h1)))
            begin
              reg1701 = (~&(+reg684));
              reg1702 <= reg684;
              for (forvar1703 = (1'h0); (forvar1703 < (2'h3)); forvar1703 = (forvar1703 + (1'h1)))
                begin
                  reg1704 <= $signed(((!((reg1669 >>> reg1673) ?
                      (wire665 ?
                          reg684 : reg686) : (forvar1687 ^~ (7'h44)))) == reg1671));
                end
              for (forvar1705 = (1'h0); (forvar1705 < (1'h1)); forvar1705 = (forvar1705 + (1'h1)))
                begin
                  reg1706 = {$unsigned("OLkI3esgDvVg"),
                      (reg950 ?
                          (((reg1688 <<< wire665) ~^ (!forvar871)) ?
                              "fZ5ourtEYKc8tOD4ACUKVN" : (!(wire1666 ?
                                  (8'h9d) : (7'h42)))) : "x1R7NN7")};
                  reg1707 <= reg675[(1'h0):(1'h0)];
                  reg1708 = (~^reg1691[(3'h5):(1'h1)]);
                  reg1709 <= $unsigned("");
                  reg1710 <= $signed(wire1445[(1'h0):(1'h0)]);
                  reg1711 <= (!$signed(({"4pV7YYNV0gC6aXBhs"} ?
                      $signed($signed(reg1681)) : reg1693[(1'h1):(1'h1)])));
                end
              reg1712 = (^~reg945);
              reg1713 <= ((($signed(reg1382[(1'h1):(1'h0)]) ?
                      ((reg1685 ?
                          reg877 : reg1690) >>> $signed(reg1697)) : reg1711) < ($signed("PlkpnMcfmW9") | reg1681[(2'h2):(2'h2)])) ?
                  wire943[(4'h9):(4'h9)] : ($signed((reg1697 ?
                      forvar1705 : (^forvar1705))) <= (wire755[(4'hb):(3'h5)] ?
                      $unsigned({reg1681, reg682}) : $signed((!reg874)))));
            end
          for (forvar1714 = (1'h0); (forvar1714 < (3'h4)); forvar1714 = (forvar1714 + (1'h1)))
            begin
              for (forvar1715 = (1'h0); (forvar1715 < (1'h0)); forvar1715 = (forvar1715 + (1'h1)))
                begin
                  reg1716 <= (^$unsigned((wire755 ?
                      $signed({reg876}) : {reg1696[(5'h14):(3'h7)],
                          {reg1690, reg875}})));
                  reg1717 = reg680[(1'h1):(1'h1)];
                  reg1718 <= ((&$signed(reg1675[(5'h11):(4'h8)])) ?
                      "X0p2V0oBKqpo7uyMHV" : (|{(7'h48)}));
                  reg1719 <= $unsigned("");
                  reg1720 = $signed(($unsigned("dly7ngRFupsekd1") == $unsigned("bAGLJmVKNuS5wJG")));
                  reg1721 <= $unsigned($unsigned($unsigned(reg946)));
                end
              reg1722 <= reg1711;
              reg1723 = wire665[(3'h5):(3'h5)];
              reg1724 <= $signed((~^(~&reg1701)));
              reg1725 <= ($signed("BJM") ?
                  (^~$unsigned($signed(((8'ha9) ?
                      forvar1692 : reg952)))) : (+(~|reg1676)));
            end
          reg1726 = "Obup";
        end
      else
        begin
          reg1699 <= "nH7aGEMA0QiJUlWs9z6LV";
          reg1700 <= forvar1377[(4'hc):(4'hb)];
        end
      reg1727 <= (-(8'hb4));
      for (forvar1728 = (1'h0); (forvar1728 < (2'h2)); forvar1728 = (forvar1728 + (1'h1)))
        begin
          reg1729 = "Oa";
          reg1730 = $unsigned({(~|$signed("Y"))});
          for (forvar1731 = (1'h0); (forvar1731 < (1'h0)); forvar1731 = (forvar1731 + (1'h1)))
            begin
              reg1732 <= ($unsigned((^~reg1723)) ?
                  reg1381 : ((^~forvar1684[(1'h1):(1'h0)]) && (("8kF1mt9nKhU30XoGuNHmApF" << "U7") ?
                      reg1695 : "Q3of6TKHRERJukVp5DW7VLXH")));
            end
          reg1733 = "1SDAkPZSziLtqE5o";
          reg1734 = forvar1728;
        end
      if (($unsigned(reg674) ? "tIrNmrSJeqU6AA6lwfu7NMrv" : (~|"WDp5e")))
        begin
          for (forvar1735 = (1'h0); (forvar1735 < (2'h3)); forvar1735 = (forvar1735 + (1'h1)))
            begin
              for (forvar1736 = (1'h0); (forvar1736 < (3'h5)); forvar1736 = (forvar1736 + (1'h1)))
                begin
                  reg1737 <= "6xOw97A0AidNGQu50dE";
                  reg1738 = reg1724;
                  reg1739 <= {((8'hae) ?
                          ({reg946[(4'hd):(3'h5)], $signed(reg676)} ?
                              "LSPuGRbZDJTzp0k" : reg870[(5'h10):(3'h7)]) : "DxxSqoiNN3dQ")};
                  reg1740 = (($signed(({reg1689} > "Fz96JltdbfgtKEQ")) ^~ "VksVmwRk1t") | forvar1692);
                end
            end
          reg1741 <= $signed(reg1672[(1'h1):(1'h0)]);
          reg1742 <= $signed(reg1739);
          reg1743 = (~&{reg1734[(5'h15):(5'h12)], (~(~^$unsigned(wire868)))});
          reg1744 <= wire667;
          if ($unsigned((8'hac)))
            begin
              for (forvar1745 = (1'h0); (forvar1745 < (3'h4)); forvar1745 = (forvar1745 + (1'h1)))
                begin
                  reg1746 = $unsigned("DVAqUwX7eCGbatr");
                  reg1747 <= (reg870[(3'h4):(2'h3)] >>> "U1C");
                end
              reg1748 <= $unsigned("M7iob");
              reg1749 <= reg1737;
            end
          else
            begin
              reg1745 <= ("tsCwGLA2Qbr8" ?
                  $unsigned($signed(forvar873[(3'h6):(3'h6)])) : reg1671);
            end
        end
      else
        begin
          for (forvar1735 = (1'h0); (forvar1735 < (1'h0)); forvar1735 = (forvar1735 + (1'h1)))
            begin
              reg1736 = reg1689[(3'h4):(1'h0)];
              reg1737 <= ($unsigned("yvJrdhWoTYap6BirRaad") ?
                  reg1727 : reg1677[(5'h16):(5'h13)]);
              reg1738 <= forvar1745[(5'h16):(5'h12)];
            end
          reg1739 <= wire666[(3'h7):(3'h6)];
          reg1740 <= $unsigned({reg879, wire1553[(3'h6):(3'h4)]});
          reg1741 <= $unsigned(wire667);
          for (forvar1742 = (1'h0); (forvar1742 < (1'h1)); forvar1742 = (forvar1742 + (1'h1)))
            begin
              reg1743 <= ((reg1668[(4'hf):(4'h9)] ?
                      $signed(reg950) : "JtQnxIfUW32") ?
                  $signed((|(~^wire1445))) : $signed($unsigned((&$unsigned(reg1376)))));
              for (forvar1744 = (1'h0); (forvar1744 < (2'h3)); forvar1744 = (forvar1744 + (1'h1)))
                begin
                  reg1745 <= reg1739[(4'ha):(3'h4)];
                  reg1746 <= {$signed((($signed(reg1745) && (^~reg1720)) * ($unsigned(wire1553) > "xJmU6K96IE1fui3VfREErO"))),
                      reg1713};
                end
              reg1747 = $signed("");
            end
        end
      reg1750 = {("ewkOHbyfCydwivN" ?
              $signed((^$signed(reg1672))) : forvar1692),
          "os"};
    end
  always
    @(posedge clk) begin
      reg1751 <= {(~&reg879[(3'h5):(2'h2)])};
      reg1752 <= "cyQcMlRSq2dUEJwT7gwcnl";
    end
  module1753 modinst1933 (wire1932, clk, reg949, forvar1700, reg1724, reg672);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module217
#( parameter param657 = ((({(7'h45), ((7'h41) && (7'h44))} ? (((7'h43) ? (8'ha1) : (7'h4d)) - ((8'ha8) && (8'hb8))) : {((8'h9d) <<< (8'ha9)), ((8'had) > (8'hba))}) ? (~({(8'hb5), (8'hbd)} ? ((8'hbb) ? (8'hbf) : (8'ha6)) : ((8'hb3) < (8'hb0)))) : {((~&(8'h9c)) + ((7'h42) == (8'hbd))), (-{(8'haa), (8'hb4)})}) | ((~&(&((7'h4e) ? (8'hba) : (7'h49)))) >= (((8'hba) ? {(8'hac), (7'h4b)} : ((8'hbc) ? (7'h43) : (8'ha8))) ? (-(8'hae)) : (((8'hba) ? (8'h9c) : (8'ha9)) && (|(8'h9f))))))
, parameter param658 = (~^param657) )
(y, clk, wire222, wire221, wire220, wire219, wire218);
  output wire [(32'h256):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire222;
  input wire signed [(5'h12):(1'h0)] wire221;
  input wire signed [(5'h11):(1'h0)] wire220;
  input wire [(4'hb):(1'h0)] wire219;
  input wire signed [(4'hc):(1'h0)] wire218;
  reg [(5'h16):(1'h0)] reg656 = (1'h0);
  reg [(5'h16):(1'h0)] reg655 = (1'h0);
  reg [(4'hc):(1'h0)] reg654 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg653 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg652 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg651 = (1'h0);
  reg [(4'hc):(1'h0)] reg650 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg649 = (1'h0);
  reg [(5'h13):(1'h0)] reg648 = (1'h0);
  reg [(4'h9):(1'h0)] reg647 = (1'h0);
  reg signed [(4'he):(1'h0)] reg646 = (1'h0);
  reg [(5'h10):(1'h0)] reg645 = (1'h0);
  reg [(5'h18):(1'h0)] reg644 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar643 = (1'h0);
  wire signed [(5'h19):(1'h0)] wire641;
  wire signed [(3'h5):(1'h0)] wire491;
  wire [(4'h9):(1'h0)] wire489;
  reg [(5'h1a):(1'h0)] reg434 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg433 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg432 = (1'h0);
  reg signed [(4'he):(1'h0)] reg431 = (1'h0);
  reg [(5'h1a):(1'h0)] reg430 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg429 = (1'h0);
  reg [(5'h17):(1'h0)] reg428 = (1'h0);
  reg [(3'h7):(1'h0)] reg427 = (1'h0);
  reg [(4'h8):(1'h0)] forvar426 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg425 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg424 = (1'h0);
  reg [(4'hc):(1'h0)] reg423 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg422 = (1'h0);
  reg [(5'h10):(1'h0)] reg421 = (1'h0);
  reg [(2'h2):(1'h0)] reg420 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar419 = (1'h0);
  reg [(4'hc):(1'h0)] forvar418 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg417 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar416 = (1'h0);
  reg [(2'h2):(1'h0)] reg415 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg414 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg413 = (1'h0);
  reg [(5'h13):(1'h0)] reg412 = (1'h0);
  reg [(4'h8):(1'h0)] reg411 = (1'h0);
  reg [(4'hc):(1'h0)] reg410 = (1'h0);
  reg [(5'h11):(1'h0)] reg409 = (1'h0);
  reg [(2'h3):(1'h0)] reg408 = (1'h0);
  wire [(2'h3):(1'h0)] wire406;
  wire [(4'hb):(1'h0)] wire223;
  assign y = {reg656,
                 reg655,
                 reg654,
                 reg653,
                 reg652,
                 reg651,
                 reg650,
                 reg649,
                 reg648,
                 reg647,
                 reg646,
                 reg645,
                 reg644,
                 forvar643,
                 wire641,
                 wire491,
                 wire489,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 forvar426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 forvar419,
                 forvar418,
                 reg417,
                 forvar416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 wire406,
                 wire223,
                 (1'h0)};
  assign wire223 = (^wire222[(4'hc):(3'h6)]);
  module224 modinst407 (.wire226(wire222), .wire227(wire220), .y(wire406), .wire225(wire221), .clk(clk), .wire228(wire219));
  always
    @(posedge clk) begin
      reg408 <= (~&"vCB");
      reg409 <= $unsigned("dC7g9IKScaI");
      reg410 <= $unsigned(("oPUW" >> ((+wire406[(1'h0):(1'h0)]) ?
          ((wire223 < reg409) >= $unsigned(wire218)) : {(wire222 > wire406)})));
      reg411 <= {(wire223[(2'h3):(1'h0)] ?
              (~^$unsigned((^wire221))) : (($signed(wire406) < $unsigned(reg410)) ?
                  (~&(wire218 ? (8'haa) : wire223)) : reg408[(1'h0):(1'h0)]))};
      reg412 <= reg410;
      reg413 <= wire222[(4'ha):(1'h1)];
    end
  always
    @(posedge clk) begin
      reg414 <= "EW2GtF88dP49N3s8e";
      reg415 <= $signed(($signed(reg409[(5'h10):(4'h8)]) && "hbMNpxiSioeExb2uP"));
      for (forvar416 = (1'h0); (forvar416 < (1'h1)); forvar416 = (forvar416 + (1'h1)))
        begin
          reg417 <= "RwyGf2MkDbrK";
          for (forvar418 = (1'h0); (forvar418 < (2'h2)); forvar418 = (forvar418 + (1'h1)))
            begin
              for (forvar419 = (1'h0); (forvar419 < (1'h1)); forvar419 = (forvar419 + (1'h1)))
                begin
                  reg420 <= "lK5tB9";
                  reg421 <= (((!(forvar419 * {wire221,
                      reg420})) | "6MhzyGuLT") <<< forvar419[(3'h5):(1'h1)]);
                  reg422 <= (~&(+reg420));
                  reg423 <= (reg415[(1'h0):(1'h0)] ?
                      $signed(forvar418) : wire221[(4'h8):(3'h6)]);
                  reg424 = $signed((reg411 ?
                      reg417 : {$unsigned(reg412),
                          ({reg412, reg423} ?
                              "vMgbDWZD6BHwYaFu0TE94" : (reg411 ?
                                  wire406 : reg423))}));
                end
              reg425 <= "G";
              for (forvar426 = (1'h0); (forvar426 < (3'h5)); forvar426 = (forvar426 + (1'h1)))
                begin
                  reg427 <= ($signed($signed($unsigned((reg408 != reg424)))) ?
                      (~(({wire222, reg411} ?
                              wire219[(4'h9):(1'h0)] : "gN9w39qGIHHb") ?
                          ($unsigned((7'h4d)) ?
                              (wire219 && reg420) : $unsigned(wire219)) : ((forvar426 != (8'hb2)) ^ (~&reg421)))) : wire222);
                end
            end
          reg428 <= {((reg427[(1'h0):(1'h0)] ?
                  (8'hbb) : (reg424 ^ {(8'hb7)})) | reg415)};
        end
      reg429 <= $unsigned("OlBpqGEHnKkqUqDqJqPUZC5");
      reg430 = (wire219 == (|$signed(wire223)));
      reg431 = $unsigned(($signed(($signed(wire222) ?
          $unsigned(reg410) : $signed(reg430))) < $unsigned(("duEd" >> (~|(8'hbf))))));
    end
  always
    @(posedge clk) begin
      reg432 <= reg429[(2'h3):(1'h1)];
      reg433 <= $signed((((^~reg421) && $signed("TxghMqlEVs")) ?
          (!wire223) : (~&$signed((forvar426 >>> reg425)))));
      reg434 = (("GPFCMAylS6gK4LTe" ?
          $unsigned("74rS") : wire223[(2'h3):(1'h0)]) > "D2Ce4s0qqCpwWX");
    end
  module435 modinst490 (wire489, clk, wire218, reg413, reg422, reg425);
  assign wire491 = (8'ha8);
  module492 modinst642 (.wire495(forvar416), .wire496(wire220), .y(wire641), .wire493(reg423), .wire494(reg417), .clk(clk));
  always
    @(posedge clk) begin
      for (forvar643 = (1'h0); (forvar643 < (2'h2)); forvar643 = (forvar643 + (1'h1)))
        begin
          reg644 <= "PAhwTWnTI8nDLbr3QoW";
        end
      reg645 = $signed(forvar426);
      reg646 <= $unsigned($unsigned($unsigned({((8'hae) ? reg425 : reg421),
          reg410})));
      reg647 <= ("k5nApJws7KrKN7" >>> ({((forvar419 ? (8'hba) : (8'hab)) ?
              (reg422 ?
                  forvar418 : reg645) : ((8'haa) | reg433))} & {($signed(reg427) + "RBTvEXO13Pfbw9bBS4tZuocon"),
          "IbASnkFyOfAZFk"}));
      reg648 <= $unsigned(reg414[(5'h15):(1'h0)]);
      reg649 = reg422[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg650 <= reg421[(5'h10):(4'hb)];
    end
  always
    @(posedge clk) begin
      reg651 = $signed((+$signed("GZb6iXnU0hpW4o9cUgBDUOe")));
      reg652 <= (&{$unsigned({{wire218}, (~|(7'h46))})});
      reg653 <= {(|$signed(reg433[(4'ha):(2'h2)])),
          (wire223 * $unsigned((reg421[(4'h9):(2'h2)] ?
              $signed(reg420) : "5pq5kCs7eesSMpp")))};
      reg654 = (~(reg415[(1'h1):(1'h1)] | ($signed((+(7'h47))) ?
          ($unsigned(reg413) ?
              reg415[(1'h1):(1'h0)] : wire489) : $signed((reg431 ?
              reg434 : reg432)))));
      reg655 <= wire218;
      reg656 <= $signed(($signed($unsigned($unsigned(reg425))) ?
          {"D5vuRxGDt8X2dbhc"} : (forvar416 << ($unsigned(reg429) ^ ((8'ha3) ?
              reg408 : wire641)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module76  (y, clk, wire77, wire78, wire79, wire80, wire81);
  output wire [(32'h3e1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire77;
  input wire signed [(5'h16):(1'h0)] wire78;
  input wire [(5'h11):(1'h0)] wire79;
  input wire [(5'h13):(1'h0)] wire80;
  input wire signed [(5'h12):(1'h0)] wire81;
  reg signed [(5'h16):(1'h0)] reg206 = (1'h0);
  reg [(4'h9):(1'h0)] reg205 = (1'h0);
  reg [(4'hf):(1'h0)] reg204 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg202 = (1'h0);
  reg [(4'hb):(1'h0)] forvar201 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg200 = (1'h0);
  reg [(3'h6):(1'h0)] reg199 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire198;
  reg signed [(5'h16):(1'h0)] reg197 = (1'h0);
  reg [(4'hb):(1'h0)] reg196 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg195 = (1'h0);
  reg [(4'hc):(1'h0)] reg194 = (1'h0);
  reg [(5'h11):(1'h0)] reg193 = (1'h0);
  reg [(4'h9):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg190 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar189 = (1'h0);
  reg [(3'h7):(1'h0)] forvar188 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg187 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg185 = (1'h0);
  reg [(4'h9):(1'h0)] forvar184 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg183 = (1'h0);
  reg [(5'h18):(1'h0)] reg182 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar181 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire82;
  reg [(4'hf):(1'h0)] reg83 = (1'h0);
  reg [(5'h1a):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar85 = (1'h0);
  reg [(4'he):(1'h0)] reg86 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar87 = (1'h0);
  reg [(5'h11):(1'h0)] forvar88 = (1'h0);
  reg signed [(4'he):(1'h0)] reg89 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg90 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar91 = (1'h0);
  reg [(4'hb):(1'h0)] reg92 = (1'h0);
  reg [(4'hb):(1'h0)] reg93 = (1'h0);
  reg [(4'he):(1'h0)] reg94 = (1'h0);
  reg [(4'he):(1'h0)] reg95 = (1'h0);
  reg [(5'h13):(1'h0)] reg96 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg97 = (1'h0);
  reg [(4'hf):(1'h0)] reg98 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg99 = (1'h0);
  reg [(3'h6):(1'h0)] reg100 = (1'h0);
  wire [(3'h6):(1'h0)] wire101;
  wire signed [(3'h5):(1'h0)] wire102;
  wire signed [(5'h17):(1'h0)] wire103;
  reg signed [(3'h5):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg106 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar105 = (1'h0);
  reg [(4'ha):(1'h0)] forvar106 = (1'h0);
  reg [(5'h10):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar109 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg110 = (1'h0);
  reg [(4'hd):(1'h0)] reg111 = (1'h0);
  reg [(4'hb):(1'h0)] reg112 = (1'h0);
  reg [(5'h17):(1'h0)] forvar113 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg114 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar115 = (1'h0);
  reg [(5'h17):(1'h0)] forvar116 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg117 = (1'h0);
  reg [(2'h2):(1'h0)] reg118 = (1'h0);
  reg [(4'ha):(1'h0)] reg119 = (1'h0);
  wire signed [(5'h16):(1'h0)] wire120;
  reg [(4'hc):(1'h0)] reg121 = (1'h0);
  reg [(2'h3):(1'h0)] reg122 = (1'h0);
  reg [(3'h7):(1'h0)] reg123 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg124 = (1'h0);
  reg [(3'h5):(1'h0)] reg125 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire126;
  wire signed [(5'h15):(1'h0)] wire179;
  assign y = {reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 forvar201,
                 reg200,
                 reg199,
                 wire198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 forvar189,
                 forvar188,
                 reg187,
                 reg186,
                 reg185,
                 forvar184,
                 reg183,
                 reg182,
                 forvar181,
                 wire82,
                 reg83,
                 reg84,
                 forvar85,
                 reg86,
                 forvar87,
                 forvar88,
                 reg89,
                 reg90,
                 forvar91,
                 reg92,
                 reg93,
                 reg94,
                 reg95,
                 reg96,
                 reg97,
                 reg98,
                 reg99,
                 reg100,
                 wire101,
                 wire102,
                 wire103,
                 reg104,
                 reg105,
                 reg106,
                 forvar105,
                 forvar106,
                 reg107,
                 reg108,
                 forvar109,
                 reg110,
                 reg111,
                 reg112,
                 forvar113,
                 reg114,
                 forvar115,
                 forvar116,
                 reg117,
                 reg118,
                 reg119,
                 wire120,
                 reg121,
                 reg122,
                 reg123,
                 reg124,
                 reg125,
                 wire126,
                 wire179,
                 (1'h0)};
  assign wire82 = wire80;
  always
    @(posedge clk) begin
      reg83 = ((&(!(((8'hbb) >= wire79) ? $signed((8'hb3)) : "ZJuTsMbU5"))) ?
          $unsigned((wire81 >> ($signed(wire81) >= wire80))) : "SaGK8");
      reg84 <= wire78[(5'h14):(4'hb)];
      for (forvar85 = (1'h0); (forvar85 < (2'h3)); forvar85 = (forvar85 + (1'h1)))
        begin
          reg86 <= ((forvar85[(2'h3):(1'h1)] << (|"")) || "qt3aWXgk");
        end
      for (forvar87 = (1'h0); (forvar87 < (3'h5)); forvar87 = (forvar87 + (1'h1)))
        begin
          for (forvar88 = (1'h0); (forvar88 < (3'h5)); forvar88 = (forvar88 + (1'h1)))
            begin
              reg89 <= reg84[(5'h19):(2'h2)];
              reg90 <= "D";
              for (forvar91 = (1'h0); (forvar91 < (1'h0)); forvar91 = (forvar91 + (1'h1)))
                begin
                  reg92 <= $unsigned($unsigned(reg90));
                  reg93 <= $signed(wire82);
                  reg94 <= ("g3OI7eEgLvltKVAD" ?
                      $signed($signed(wire79)) : reg90[(3'h5):(2'h2)]);
                  reg95 = $signed("LXXq38BwnAdfI1E");
                  reg96 <= "Xk3fHbWlBIF2k1qbAvu7KX";
                  reg97 = $unsigned($unsigned(forvar91));
                end
              reg98 <= forvar88[(2'h2):(2'h2)];
              reg99 <= $unsigned($signed({{(reg86 ? wire82 : reg86),
                      "ESRHiap"}}));
            end
          reg100 <= (+((|reg99[(2'h3):(1'h0)]) ? {(8'ha3)} : (~&reg96)));
        end
    end
  assign wire101 = "E8T61xS92ylgmcey4qRD";
  assign wire102 = ("UZcgEVR" || "TFf4riP91zEzq0w0C");
  assign wire103 = (({wire101, wire102[(1'h1):(1'h0)]} ~^ {({reg95, reg98} ?
                               (wire79 ? reg86 : forvar91) : (^~(8'hb1))),
                           $signed($unsigned(reg94))}) ?
                       (~((-$unsigned(reg89)) ?
                           $signed("Knwg91ZcquCq2b") : "4H")) : (7'h42));
  always
    @(posedge clk) begin
      if ("bBhx3Oicr")
        begin
          reg104 <= wire77[(1'h1):(1'h1)];
          reg105 <= $signed(reg98[(1'h1):(1'h1)]);
          reg106 <= "iT3";
        end
      else
        begin
          reg104 <= (($unsigned((reg86[(3'h4):(1'h1)] - (+reg93))) ?
                  $signed($unsigned(wire81)) : wire103[(4'ha):(3'h4)]) ?
              $unsigned("xUixPoKvyHQieZlXgM") : $signed((($signed(reg83) ?
                      reg89 : (reg83 ? (7'h47) : reg86)) ?
                  "" : $unsigned("WLzJDKFgeIB"))));
          for (forvar105 = (1'h0); (forvar105 < (1'h1)); forvar105 = (forvar105 + (1'h1)))
            begin
              for (forvar106 = (1'h0); (forvar106 < (3'h5)); forvar106 = (forvar106 + (1'h1)))
                begin
                  reg107 = (reg90 ? reg84[(5'h15):(5'h13)] : $unsigned(reg95));
                end
              reg108 <= (~$signed($unsigned(((+(7'h48)) != (wire101 >> wire77)))));
            end
          for (forvar109 = (1'h0); (forvar109 < (3'h5)); forvar109 = (forvar109 + (1'h1)))
            begin
              reg110 = wire81;
              reg111 <= ((-("OwVI29Wy7vkPb06LT" ?
                      reg108 : (~|forvar105[(4'h8):(3'h7)]))) ?
                  $signed((&"t")) : $signed((reg104[(1'h1):(1'h1)] ?
                      ((wire102 <= wire81) ?
                          reg99[(2'h3):(1'h1)] : reg98) : {(reg107 ?
                              wire101 : (8'hb4)),
                          (reg96 * reg98)})));
              reg112 = (($unsigned((((7'h46) << wire102) ?
                      $unsigned(wire103) : (reg111 ^ reg94))) ?
                  (wire82[(1'h1):(1'h1)] == (^~"N8A")) : ((~$signed(wire82)) ?
                      "ZtRU3hUJkmKb" : ((forvar88 ?
                          reg105 : forvar109) < forvar106))) ^ reg110);
              for (forvar113 = (1'h0); (forvar113 < (2'h2)); forvar113 = (forvar113 + (1'h1)))
                begin
                  reg114 <= $signed(((8'hab) ?
                      $signed((((8'ha5) ?
                          wire81 : wire103) * (8'hbb))) : (!$unsigned(reg94))));
                end
            end
          for (forvar115 = (1'h0); (forvar115 < (3'h4)); forvar115 = (forvar115 + (1'h1)))
            begin
              for (forvar116 = (1'h0); (forvar116 < (3'h5)); forvar116 = (forvar116 + (1'h1)))
                begin
                  reg117 <= $signed(reg94);
                end
            end
        end
      reg118 <= "2cf1ZC4pEJEd4r";
      reg119 <= $unsigned((((forvar105[(3'h6):(3'h6)] ?
                  (|forvar91) : (!reg104)) ?
              ((-forvar88) ?
                  $unsigned(reg83) : (+(7'h47))) : (reg117[(3'h6):(3'h6)] <<< {reg105})) ?
          reg114[(5'h17):(5'h11)] : $unsigned((wire80 > (reg92 <= reg108)))));
    end
  assign wire120 = $unsigned((forvar85 ?
                       forvar109[(2'h2):(2'h2)] : $signed($unsigned($unsigned(reg84)))));
  always
    @(posedge clk) begin
      reg121 <= ($unsigned($signed("f0ppb7tJyEwmPyJXML")) ?
          forvar113[(4'hf):(2'h3)] : $unsigned("yLnpxQQbSQZGtH"));
      reg122 <= ("2pF8bseJo" ?
          (("8zfIzpHGJ3UIy" >> ($signed(reg106) & {(7'h41)})) - ($unsigned((~&forvar116)) >>> $unsigned($signed((8'ha2))))) : (8'hbe));
      reg123 = $signed(((|{reg98, wire77}) != forvar85));
      reg124 <= forvar85[(2'h3):(1'h1)];
      reg125 <= "i3h5FDqItfPkL22f9EvLr9rHA";
    end
  assign wire126 = ($signed(forvar91[(3'h6):(3'h5)]) > "GheRIKdUe4xvEdD87yu4ZNTI");
  module127 modinst180 (wire179, clk, reg111, reg86, forvar113, reg96, forvar85);
  always
    @(posedge clk) begin
      for (forvar181 = (1'h0); (forvar181 < (3'h4)); forvar181 = (forvar181 + (1'h1)))
        begin
          reg182 <= reg104;
        end
      reg183 <= $signed($signed("OPf2ZpXsWSELmC4J"));
      for (forvar184 = (1'h0); (forvar184 < (2'h3)); forvar184 = (forvar184 + (1'h1)))
        begin
          reg185 = $signed("mJlDI");
          reg186 <= $signed(wire79);
          reg187 <= "oFMbFRDbMG6SBiiD2P";
        end
      for (forvar188 = (1'h0); (forvar188 < (3'h5)); forvar188 = (forvar188 + (1'h1)))
        begin
          for (forvar189 = (1'h0); (forvar189 < (2'h3)); forvar189 = (forvar189 + (1'h1)))
            begin
              reg190 <= {forvar184[(2'h3):(1'h1)]};
              reg191 = wire79;
              reg192 <= "dmaWJXwhg";
            end
          reg193 <= "I3Nlh33paRtwuPpy4MB5r";
          reg194 <= $unsigned(forvar115[(5'h10):(5'h10)]);
          reg195 <= ((reg114[(5'h14):(5'h14)] != $signed($signed((reg186 | wire78)))) ?
              ($signed("8NUBZ8RywKl9iJ") ?
                  {reg93} : ($unsigned($unsigned(reg182)) < wire78[(4'h8):(3'h7)])) : forvar105);
          reg196 <= reg185[(5'h17):(4'hd)];
          reg197 <= $unsigned((!({(reg195 >>> forvar181)} | (((8'h9d) ?
                  (7'h49) : wire103) ?
              forvar109[(5'h10):(2'h3)] : reg182[(1'h0):(1'h0)]))));
        end
    end
  assign wire198 = reg99;
  always
    @(posedge clk) begin
      reg199 = ((($signed((~|wire120)) >= {wire179, $signed(forvar184)}) ?
              "fWbsqyxO" : "4Yy2kSRu0") ?
          (+"UAZ14MtgnJwNp5LrK2at") : reg100);
      reg200 = reg106[(2'h3):(1'h0)];
      for (forvar201 = (1'h0); (forvar201 < (3'h4)); forvar201 = (forvar201 + (1'h1)))
        begin
          reg202 <= (!"OOAKHkvn1aJdBJCeGWMW");
          reg203 = (((reg106[(4'hf):(3'h7)] ?
                  ((~^(8'ha3)) ? $signed(reg121) : (~(7'h42))) : {{reg202},
                      forvar88[(4'hc):(4'h9)]}) ?
              (($unsigned((7'h44)) ?
                      ((8'hb8) ? forvar181 : (8'hba)) : (reg95 + forvar106)) ?
                  "slQtyHsWIDw" : $unsigned($unsigned(reg100))) : reg90[(4'h9):(3'h6)]) ^~ $signed({(&((8'ha5) ?
                  reg199 : wire79)),
              reg107}));
          reg204 <= $unsigned({(^$signed((reg191 == wire126))), "uXeA"});
        end
      reg205 = {reg197};
      reg206 = "V9NsVPmrEeCR";
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module127
#( parameter param178 = ((^~((8'ha0) * ((^(7'h41)) - (7'h4a)))) | (({((8'hb1) ? (8'hbd) : (8'ha2))} >> (8'hb3)) ? {(((8'ha8) || (8'hb5)) ^ ((8'h9f) + (8'ha0))), (((8'hb2) ? (8'hb2) : (8'ha5)) ? {(8'ha4), (8'hb3)} : ((7'h4b) ? (7'h4a) : (7'h42)))} : (^{((7'h4c) ? (7'h49) : (7'h49)), ((8'h9e) ? (8'ha0) : (8'hb3))}))) )
(y, clk, wire132, wire131, wire130, wire129, wire128);
  output wire [(32'h280):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire132;
  input wire [(3'h6):(1'h0)] wire131;
  input wire [(4'ha):(1'h0)] wire130;
  input wire [(4'hb):(1'h0)] wire129;
  input wire signed [(4'hd):(1'h0)] wire128;
  reg [(4'he):(1'h0)] reg177 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar176 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg175 = (1'h0);
  reg [(5'h11):(1'h0)] reg174 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg172 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg171 = (1'h0);
  reg [(3'h6):(1'h0)] reg170 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg168 = (1'h0);
  reg [(3'h6):(1'h0)] reg167 = (1'h0);
  reg [(5'h12):(1'h0)] reg166 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg165 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg164 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar163 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg162 = (1'h0);
  reg [(5'h15):(1'h0)] forvar161 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar160 = (1'h0);
  reg [(4'h8):(1'h0)] reg159 = (1'h0);
  reg [(5'h19):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg157 = (1'h0);
  reg [(3'h7):(1'h0)] reg156 = (1'h0);
  reg [(5'h17):(1'h0)] reg155 = (1'h0);
  reg [(3'h6):(1'h0)] reg154 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar153 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg152 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg150 = (1'h0);
  reg [(5'h1a):(1'h0)] reg149 = (1'h0);
  reg [(4'hb):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar147 = (1'h0);
  reg [(2'h2):(1'h0)] forvar146 = (1'h0);
  reg [(4'hc):(1'h0)] reg145 = (1'h0);
  reg [(4'hc):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg142 = (1'h0);
  reg [(4'hf):(1'h0)] reg141 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg140 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg139 = (1'h0);
  wire [(5'h1a):(1'h0)] wire138;
  reg [(5'h15):(1'h0)] reg137 = (1'h0);
  reg [(2'h3):(1'h0)] reg136 = (1'h0);
  reg [(4'hd):(1'h0)] forvar135 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg134 = (1'h0);
  wire [(4'h8):(1'h0)] wire133;
  assign y = {reg177,
                 forvar176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 forvar163,
                 reg162,
                 forvar161,
                 forvar160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 forvar153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 forvar147,
                 forvar146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 wire138,
                 reg137,
                 reg136,
                 forvar135,
                 reg134,
                 wire133,
                 (1'h0)};
  assign wire133 = $unsigned($signed("olVD8Fn6mDWlWTToe5HKnhLe"));
  always
    @(posedge clk) begin
      reg134 <= ((((!{wire129, wire132}) ?
              {(wire133 - wire128), $signed(wire133)} : ($unsigned(wire132) ?
                  wire128 : (^wire133))) * wire131) ?
          wire129 : $unsigned((({wire131, wire128} == {(8'hb8)}) ?
              wire132[(2'h3):(1'h1)] : ("BNr" ^~ "mhsNqnEM"))));
      for (forvar135 = (1'h0); (forvar135 < (1'h1)); forvar135 = (forvar135 + (1'h1)))
        begin
          reg136 = (^~$unsigned((+$unsigned("V"))));
          reg137 <= ((~|(!wire128)) >= $unsigned(wire128[(4'h9):(3'h5)]));
        end
    end
  assign wire138 = $signed(wire128);
  always
    @(posedge clk) begin
      reg139 <= (~^(|(({forvar135} ? reg136 : (~(8'hb1))) ?
          ((wire133 ? wire130 : (7'h4b)) ?
              $signed(wire138) : (+wire138)) : (~|$unsigned((7'h40))))));
    end
  always
    @(posedge clk) begin
      reg140 <= ($signed($signed($unsigned((reg139 ? wire131 : wire130)))) ?
          wire131[(2'h3):(2'h3)] : "MXaGIM");
      reg141 <= wire131;
    end
  always
    @(posedge clk) begin
      reg142 <= ($signed("svr6dr9T") ?
          $unsigned($unsigned($unsigned((-reg134)))) : (!{reg139}));
      reg143 = {reg141[(3'h7):(3'h4)]};
    end
  always
    @(posedge clk) begin
      reg144 <= (!$unsigned({((8'h9d) + (~reg143)), reg141}));
    end
  always
    @(posedge clk) begin
      reg145 <= (-(reg141[(1'h1):(1'h1)] + (((~&reg136) ^ (wire129 != reg137)) != wire128[(1'h0):(1'h0)])));
      for (forvar146 = (1'h0); (forvar146 < (1'h0)); forvar146 = (forvar146 + (1'h1)))
        begin
          for (forvar147 = (1'h0); (forvar147 < (1'h1)); forvar147 = (forvar147 + (1'h1)))
            begin
              reg148 <= "Kp4Zuxy2NKoLw3vP0pVcKs6q";
              reg149 <= (~|{$unsigned((~^reg134[(1'h1):(1'h1)]))});
              reg150 <= reg141[(3'h6):(3'h4)];
              reg151 <= wire138;
              reg152 <= {forvar147,
                  ({("ZmgNViK1tzKb5KlsEZ" ?
                              (forvar146 ? reg145 : forvar147) : reg136),
                          $unsigned($unsigned((7'h42)))} ?
                      ($unsigned(reg136) != (reg151 > $signed(reg149))) : reg144[(3'h4):(1'h1)])};
              for (forvar153 = (1'h0); (forvar153 < (2'h3)); forvar153 = (forvar153 + (1'h1)))
                begin
                  reg154 <= $unsigned($signed($unsigned((8'hb8))));
                  reg155 <= forvar153;
                  reg156 <= {((^$unsigned({reg144, (8'hb9)})) ?
                          wire131[(3'h6):(2'h2)] : $unsigned($signed(wire131[(3'h5):(1'h1)]))),
                      "9umXgGpk1BB1UhJFObcSeyTXm"};
                  reg157 <= $signed(reg148);
                  reg158 <= (^wire129[(4'h9):(1'h0)]);
                end
            end
          reg159 <= (&$signed($unsigned((reg143[(2'h2):(1'h0)] ?
              (reg156 ? wire130 : reg144) : $unsigned(reg134)))));
          for (forvar160 = (1'h0); (forvar160 < (3'h4)); forvar160 = (forvar160 + (1'h1)))
            begin
              for (forvar161 = (1'h0); (forvar161 < (2'h2)); forvar161 = (forvar161 + (1'h1)))
                begin
                  reg162 <= ("a9gnWdnE3C9siHyFUtqXni2" ?
                      $unsigned($unsigned($unsigned("8OBiKRHYQ0QVVWKSC11nXDi"))) : "Er1uemIxmgACBNtW");
                end
              for (forvar163 = (1'h0); (forvar163 < (2'h2)); forvar163 = (forvar163 + (1'h1)))
                begin
                  reg164 <= ("rGPudm" ? (!(8'hbd)) : reg158[(4'hd):(4'h8)]);
                  reg165 = $unsigned(($unsigned(reg152) != {(~&$signed(reg159))}));
                end
              if ((8'hb9))
                begin
                  reg166 = ((8'hac) ~^ (&(reg164[(3'h7):(2'h3)] ?
                      forvar153[(5'h14):(1'h0)] : ($unsigned(reg165) ?
                          $signed(reg134) : reg134[(1'h0):(1'h0)]))));
                  reg167 <= $unsigned((7'h45));
                  reg168 <= (reg157[(1'h1):(1'h1)] != $unsigned({{(reg142 ?
                              reg150 : reg159),
                          (^reg162)},
                      ({wire130} ? (reg149 ~^ reg134) : {(7'h49), wire138})}));
                end
              else
                begin
                  reg166 = wire133;
                  reg167 <= reg134;
                  reg168 <= "vnYhJ";
                end
              reg169 <= (reg166 & (8'hb7));
              reg170 <= $unsigned($signed(reg144[(3'h5):(1'h1)]));
              reg171 <= ((&$unsigned(reg141[(4'h9):(3'h7)])) ?
                  forvar147 : $unsigned($unsigned("3ao1xXmry4rdAzoJ2moot")));
            end
          reg172 <= {reg154, "1e7aGMC"};
        end
      reg173 <= reg144[(4'h9):(4'h9)];
      reg174 = $unsigned(forvar160[(5'h13):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg175 <= "rDpn2ymFYZvxZ85Bq";
      for (forvar176 = (1'h0); (forvar176 < (1'h0)); forvar176 = (forvar176 + (1'h1)))
        begin
          reg177 <= $signed($signed((~^(~|reg142))));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module492
#( parameter param639 = (~|(((((8'hb8) ? (8'haa) : (7'h41)) ? ((7'h4c) ? (8'ha9) : (7'h48)) : (^~(8'hb9))) ? (&(~|(7'h44))) : (^((8'ha5) | (8'ha0)))) & (+({(8'ha2)} | ((8'hbd) ? (8'hbf) : (8'hb3))))))
, parameter param640 = param639 )
(y, clk, wire496, wire495, wire494, wire493);
  output wire [(32'h74e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire496;
  input wire [(5'h11):(1'h0)] wire495;
  input wire signed [(5'h10):(1'h0)] wire494;
  input wire [(4'hc):(1'h0)] wire493;
  reg [(5'h16):(1'h0)] reg638 = (1'h0);
  reg [(3'h7):(1'h0)] reg637 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg636 = (1'h0);
  reg signed [(4'he):(1'h0)] reg635 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg634 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg633 = (1'h0);
  reg [(5'h11):(1'h0)] reg632 = (1'h0);
  reg [(4'hd):(1'h0)] reg631 = (1'h0);
  reg [(4'hc):(1'h0)] reg630 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg629 = (1'h0);
  reg [(5'h16):(1'h0)] reg628 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg627 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg626 = (1'h0);
  reg [(4'h9):(1'h0)] forvar625 = (1'h0);
  reg [(4'hd):(1'h0)] reg624 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire623;
  reg [(3'h4):(1'h0)] reg622 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg621 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg620 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar619 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg618 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg617 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg616 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar615 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg614 = (1'h0);
  reg [(4'h9):(1'h0)] reg613 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg612 = (1'h0);
  reg [(3'h7):(1'h0)] reg611 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg610 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar609 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg608 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg607 = (1'h0);
  wire [(4'he):(1'h0)] wire606;
  wire [(5'h13):(1'h0)] wire605;
  reg [(4'hd):(1'h0)] reg604 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg603 = (1'h0);
  reg [(5'h16):(1'h0)] reg602 = (1'h0);
  reg [(3'h5):(1'h0)] reg601 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg600 = (1'h0);
  reg [(3'h6):(1'h0)] reg599 = (1'h0);
  reg [(4'h9):(1'h0)] reg598 = (1'h0);
  reg [(4'h9):(1'h0)] reg597 = (1'h0);
  reg [(4'hf):(1'h0)] reg596 = (1'h0);
  reg [(4'he):(1'h0)] reg595 = (1'h0);
  wire signed [(4'he):(1'h0)] wire594;
  wire signed [(4'h9):(1'h0)] wire593;
  wire [(5'h1a):(1'h0)] wire592;
  reg [(5'h1a):(1'h0)] reg591 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg590 = (1'h0);
  reg [(4'h8):(1'h0)] reg589 = (1'h0);
  reg [(3'h7):(1'h0)] reg588 = (1'h0);
  reg [(4'h9):(1'h0)] reg587 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg586 = (1'h0);
  reg [(2'h3):(1'h0)] reg585 = (1'h0);
  reg [(4'hb):(1'h0)] forvar584 = (1'h0);
  reg [(5'h17):(1'h0)] reg583 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg582 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg581 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire580;
  wire [(3'h6):(1'h0)] wire579;
  reg [(3'h7):(1'h0)] reg578 = (1'h0);
  reg [(3'h4):(1'h0)] reg577 = (1'h0);
  reg [(5'h12):(1'h0)] reg576 = (1'h0);
  wire [(5'h10):(1'h0)] wire575;
  wire [(2'h2):(1'h0)] wire574;
  reg [(3'h5):(1'h0)] reg573 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg572 = (1'h0);
  reg [(3'h6):(1'h0)] reg571 = (1'h0);
  reg [(4'hf):(1'h0)] reg570 = (1'h0);
  reg signed [(4'he):(1'h0)] reg569 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar568 = (1'h0);
  reg [(5'h11):(1'h0)] reg567 = (1'h0);
  reg [(5'h18):(1'h0)] reg566 = (1'h0);
  reg [(5'h10):(1'h0)] reg565 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg563 = (1'h0);
  reg [(3'h7):(1'h0)] reg562 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg561 = (1'h0);
  reg [(2'h3):(1'h0)] forvar560 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg559 = (1'h0);
  reg [(3'h6):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg557 = (1'h0);
  reg [(5'h16):(1'h0)] forvar556 = (1'h0);
  reg [(5'h17):(1'h0)] forvar555 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar554 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg553 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg552 = (1'h0);
  reg [(3'h5):(1'h0)] reg551 = (1'h0);
  reg [(4'ha):(1'h0)] reg550 = (1'h0);
  reg [(5'h12):(1'h0)] reg549 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg548 = (1'h0);
  reg [(5'h18):(1'h0)] reg547 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg546 = (1'h0);
  reg [(4'h9):(1'h0)] reg545 = (1'h0);
  reg [(5'h16):(1'h0)] reg544 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg543 = (1'h0);
  reg [(5'h12):(1'h0)] forvar542 = (1'h0);
  reg [(3'h5):(1'h0)] reg541 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg540 = (1'h0);
  reg [(3'h5):(1'h0)] reg539 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg538 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg537 = (1'h0);
  reg [(4'h8):(1'h0)] reg536 = (1'h0);
  reg [(4'hc):(1'h0)] forvar535 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg534 = (1'h0);
  reg [(5'h17):(1'h0)] reg533 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar531 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg526 = (1'h0);
  reg [(4'hc):(1'h0)] forvar525 = (1'h0);
  reg [(2'h2):(1'h0)] reg530 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg529 = (1'h0);
  reg [(2'h3):(1'h0)] reg528 = (1'h0);
  reg [(4'he):(1'h0)] reg527 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar526 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg525 = (1'h0);
  reg [(5'h14):(1'h0)] reg524 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar523 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg522 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg521 = (1'h0);
  reg [(3'h5):(1'h0)] reg520 = (1'h0);
  reg [(4'hf):(1'h0)] forvar519 = (1'h0);
  reg [(4'he):(1'h0)] reg518 = (1'h0);
  reg [(4'hf):(1'h0)] reg517 = (1'h0);
  reg [(3'h7):(1'h0)] reg516 = (1'h0);
  reg [(5'h1a):(1'h0)] reg515 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar514 = (1'h0);
  reg [(3'h7):(1'h0)] reg513 = (1'h0);
  wire [(5'h19):(1'h0)] wire512;
  wire signed [(5'h10):(1'h0)] wire511;
  reg signed [(5'h12):(1'h0)] reg510 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg509 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg508 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg507 = (1'h0);
  reg [(3'h7):(1'h0)] reg506 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg505 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar504 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg503 = (1'h0);
  reg [(5'h12):(1'h0)] reg502 = (1'h0);
  reg [(5'h19):(1'h0)] forvar501 = (1'h0);
  reg [(3'h6):(1'h0)] reg500 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg499 = (1'h0);
  reg [(5'h13):(1'h0)] reg498 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg497 = (1'h0);
  assign y = {reg638,
                 reg637,
                 reg636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 forvar625,
                 reg624,
                 wire623,
                 reg622,
                 reg621,
                 reg620,
                 forvar619,
                 reg618,
                 reg617,
                 reg616,
                 forvar615,
                 reg614,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 forvar609,
                 reg608,
                 reg607,
                 wire606,
                 wire605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 wire594,
                 wire593,
                 wire592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 reg586,
                 reg585,
                 forvar584,
                 reg583,
                 reg582,
                 reg581,
                 wire580,
                 wire579,
                 reg578,
                 reg577,
                 reg576,
                 wire575,
                 wire574,
                 reg573,
                 reg572,
                 reg571,
                 reg570,
                 reg569,
                 forvar568,
                 reg567,
                 reg566,
                 reg565,
                 reg564,
                 reg563,
                 reg562,
                 reg561,
                 forvar560,
                 reg559,
                 reg558,
                 reg557,
                 forvar556,
                 forvar555,
                 forvar554,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 reg543,
                 forvar542,
                 reg541,
                 reg540,
                 reg539,
                 reg538,
                 reg537,
                 reg536,
                 forvar535,
                 reg534,
                 reg533,
                 reg532,
                 forvar531,
                 reg526,
                 forvar525,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 forvar526,
                 reg525,
                 reg524,
                 forvar523,
                 reg522,
                 reg521,
                 reg520,
                 forvar519,
                 reg518,
                 reg517,
                 reg516,
                 reg515,
                 forvar514,
                 reg513,
                 wire512,
                 wire511,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 forvar504,
                 reg503,
                 reg502,
                 forvar501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg497 <= wire493;
      reg498 = ((^($signed(wire495[(5'h10):(4'hd)]) ?
              ($signed(wire493) != $unsigned(reg497)) : $unsigned("6EKvX7WG"))) ?
          (wire493 ?
              ((~^(reg497 ? (8'ha5) : wire493)) ^~ ($signed(reg497) ?
                  ((8'h9f) ?
                      wire494 : wire494) : reg497)) : wire496[(3'h7):(3'h7)]) : ((^~wire495) >= "Tsg09smq"));
      reg499 <= $signed($signed($unsigned((~^$unsigned(reg498)))));
    end
  always
    @(posedge clk) begin
      reg500 <= (("TQPYYPgWthoe9Q7EqR1p" ?
          wire493 : (~(|"PAGgoS1PFMv5kV"))) <<< wire493);
      for (forvar501 = (1'h0); (forvar501 < (2'h2)); forvar501 = (forvar501 + (1'h1)))
        begin
          reg502 <= $unsigned((wire493 ? $unsigned(wire494) : wire493));
          reg503 <= "FX6rP2AVXC2okxgr9637it9m";
          for (forvar504 = (1'h0); (forvar504 < (3'h5)); forvar504 = (forvar504 + (1'h1)))
            begin
              reg505 <= (~^{"fWRR7PhMzOEnwDwOOwXApdALG"});
              reg506 = ((8'hb4) ?
                  ((~|((^~wire493) ?
                          $unsigned(reg505) : $unsigned(forvar501))) ?
                      ((8'hba) - reg499[(1'h0):(1'h0)]) : $signed(reg505[(4'hc):(3'h5)])) : reg500);
              reg507 <= forvar501;
              reg508 <= reg498;
              reg509 <= "sHi92AlHbkS";
            end
          reg510 <= (((|"2yE2YIVwRRtVTZPPkFN") ~^ reg506) - ((reg497 & $unsigned(reg502[(1'h0):(1'h0)])) != ($signed((~&wire496)) ?
              reg505[(3'h7):(1'h1)] : $unsigned(forvar501))));
        end
    end
  assign wire511 = {forvar501};
  assign wire512 = reg508[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      reg513 <= (~&"RkIWQXq03");
    end
  always
    @(posedge clk) begin
      for (forvar514 = (1'h0); (forvar514 < (2'h3)); forvar514 = (forvar514 + (1'h1)))
        begin
          reg515 <= $signed(forvar504);
          reg516 <= (8'h9c);
          reg517 = "b9wmZUTXVMZQhL";
          reg518 <= reg498;
        end
      for (forvar519 = (1'h0); (forvar519 < (1'h0)); forvar519 = (forvar519 + (1'h1)))
        begin
          reg520 <= (!{$signed($signed({reg505}))});
        end
      reg521 = $signed({((|(~&reg509)) ^ $unsigned(reg507))});
      reg522 <= (8'ha9);
    end
  always
    @(posedge clk) begin
      for (forvar523 = (1'h0); (forvar523 < (2'h3)); forvar523 = (forvar523 + (1'h1)))
        begin
          if (("o" ?
              (&(-((^reg497) ?
                  (^~reg500) : "OIWcLLAp"))) : ($unsigned({$signed(reg517),
                      (reg513 ? (8'hbf) : reg513)}) ?
                  ($unsigned({reg513}) ?
                      reg516 : ((+forvar501) ?
                          $unsigned(forvar519) : reg498[(4'hf):(3'h5)])) : "0rtfBwSX3WHl1p")))
            begin
              reg524 = forvar501;
              reg525 <= "yQ7eB9hK3axq5nECWyyW";
              for (forvar526 = (1'h0); (forvar526 < (1'h0)); forvar526 = (forvar526 + (1'h1)))
                begin
                  reg527 = forvar504;
                  reg528 <= wire511;
                end
              reg529 <= "TyFdlKNCw";
              reg530 <= $signed((^~(($unsigned(wire493) ?
                      $signed(wire494) : forvar504) ?
                  $unsigned($unsigned(forvar519)) : $unsigned((8'hba)))));
            end
          else
            begin
              reg524 <= (reg521[(1'h0):(1'h0)] >= (|"4koergZ4"));
              for (forvar525 = (1'h0); (forvar525 < (1'h0)); forvar525 = (forvar525 + (1'h1)))
                begin
                  reg526 <= ({(^$unsigned({(8'hbb)})),
                      (~forvar526[(3'h6):(3'h4)])} > reg497[(4'h8):(3'h6)]);
                  reg527 <= forvar526[(2'h3):(2'h3)];
                  reg528 = "SFJBMHYJCdKGh2ULe4vS";
                  reg529 <= forvar523[(1'h1):(1'h0)];
                  reg530 = (~|reg513);
                end
              for (forvar531 = (1'h0); (forvar531 < (3'h5)); forvar531 = (forvar531 + (1'h1)))
                begin
                  reg532 <= reg500[(1'h1):(1'h0)];
                  reg533 <= "UGCtN51";
                end
              reg534 <= {{$unsigned("xSV9gaCC8N1XxqLL9XRYoEp2"),
                      ("ulgdvaOpo7Wc" ?
                          (~(reg510 ?
                              wire496 : reg517)) : $unsigned("26fvn7DtT6T"))},
                  wire493[(1'h0):(1'h0)]};
              for (forvar535 = (1'h0); (forvar535 < (1'h1)); forvar535 = (forvar535 + (1'h1)))
                begin
                  reg536 <= $signed(wire495);
                  reg537 <= reg516[(3'h4):(2'h3)];
                  reg538 <= $signed(reg507);
                  reg539 <= (-$unsigned(reg518));
                  reg540 <= "6BQXP5uVB";
                  reg541 <= $signed($signed((("1zoQ4DuLnlcryEOoFKC" ^~ (7'h4b)) ?
                      ({forvar535, wire493} >> wire494) : "LiNneB4ybL")));
                end
              for (forvar542 = (1'h0); (forvar542 < (1'h0)); forvar542 = (forvar542 + (1'h1)))
                begin
                  reg543 <= (reg520[(1'h0):(1'h0)] ^~ {reg497[(2'h2):(1'h0)],
                      ({((7'h48) == reg510)} ~^ ({wire512} ?
                          reg525 : "yFZZERz6"))});
                  reg544 <= (^"IxE1");
                  reg545 <= "2AuL";
                  reg546 <= reg540[(2'h3):(2'h2)];
                  reg547 <= "00mKBxOeOgFnMv";
                end
            end
          reg548 <= (forvar519[(3'h5):(3'h4)] ?
              ($signed(reg515[(5'h16):(4'hd)]) + $unsigned(($unsigned((8'hb6)) ^~ forvar526))) : "8sB");
          reg549 <= $signed(((~|reg525) ?
              forvar531 : ($unsigned($signed(reg547)) ?
                  (&reg505[(4'hf):(4'hd)]) : reg527)));
          reg550 <= "3dM9rOUrm5nmH6OdU";
          reg551 <= ((^(&(~^(~|reg499)))) ?
              wire493 : $signed(($signed($signed(wire511)) ?
                  wire495 : reg530)));
        end
      reg552 <= $unsigned("n");
      reg553 = {{$unsigned(($signed(forvar504) ?
                  $signed((8'ha8)) : (reg521 && wire495)))},
          reg541[(1'h0):(1'h0)]};
      for (forvar554 = (1'h0); (forvar554 < (2'h2)); forvar554 = (forvar554 + (1'h1)))
        begin
          for (forvar555 = (1'h0); (forvar555 < (2'h3)); forvar555 = (forvar555 + (1'h1)))
            begin
              for (forvar556 = (1'h0); (forvar556 < (2'h3)); forvar556 = (forvar556 + (1'h1)))
                begin
                  reg557 = $unsigned(forvar535);
                  reg558 <= $signed("lbLaYDM2WLuGp7");
                end
              reg559 <= wire511[(4'hb):(4'ha)];
              for (forvar560 = (1'h0); (forvar560 < (1'h1)); forvar560 = (forvar560 + (1'h1)))
                begin
                  reg561 <= ($unsigned("Pdxlt5HWl") <= {$signed((reg516 ?
                          (reg543 ? reg534 : reg559) : (~|wire494)))});
                  reg562 <= reg525[(4'hb):(4'hb)];
                  reg563 <= $unsigned(((^~$unsigned($signed(reg525))) ?
                      reg506 : $signed($signed({reg532, reg529}))));
                  reg564 = ((("c" ? reg550 : forvar525) ?
                      (reg548 ~^ $unsigned(reg521)) : ($signed({wire512,
                          reg562}) > {"gqJV6oRkvyeyP4SpsO"})) & $signed((&(~reg529))));
                end
              reg565 <= ((reg559[(4'ha):(3'h7)] ?
                  ((wire496 & (~|forvar556)) ?
                      ((reg527 ?
                          reg509 : reg534) <= reg533) : (~((7'h45) >> reg500))) : (forvar535 || (^~$signed(reg508)))) <= reg529);
              reg566 <= $unsigned((forvar555 | reg502));
              reg567 <= forvar555;
            end
          for (forvar568 = (1'h0); (forvar568 < (2'h3)); forvar568 = (forvar568 + (1'h1)))
            begin
              reg569 <= {(reg544 ^ reg559[(3'h6):(3'h6)])};
              reg570 <= (~|$unsigned(reg499));
              reg571 <= ((|($unsigned($signed(reg565)) ~^ (8'h9c))) > $unsigned(forvar542[(5'h11):(4'hc)]));
              reg572 <= (reg543[(4'hc):(4'hb)] ?
                  ($unsigned({$unsigned((7'h40)), $unsigned(reg538)}) ?
                      "Miwr" : $unsigned((8'ha6))) : reg513[(1'h0):(1'h0)]);
            end
        end
      reg573 <= (8'hb3);
    end
  assign wire574 = (reg498 ? $unsigned("BLLvoJFQx50RPkx") : forvar535);
  assign wire575 = ($signed($unsigned($unsigned((forvar554 ?
                       reg540 : forvar531)))) <= (!(reg548 ?
                       wire512[(5'h10):(1'h1)] : ($unsigned(reg532) && (reg569 ?
                           reg552 : reg522)))));
  always
    @(posedge clk) begin
      reg576 <= ("0XnEPI37HfAx4r4vwHJU36Zwy" == ("oTdb" ?
          reg543 : (+(~^((8'hac) ? reg571 : reg524)))));
      reg577 <= (!("sNBM1n3S7EddwJGASK1oY0mna" ?
          (|(8'hbb)) : (~^(reg522 ^ reg498))));
      reg578 <= {"3yDma"};
    end
  assign wire579 = "Ea0G";
  assign wire580 = (~|({{{reg550, reg536}, {wire493}}, reg508[(1'h1):(1'h1)]} ?
                       (((reg508 ?
                           wire579 : reg510) & $signed(forvar542)) < (+"Y6ea0VmPIvZQYUd1r7")) : ("ioRB9" ?
                           ("0NzcPLdB" + {forvar556,
                               reg521}) : $signed($signed(reg550)))));
  always
    @(posedge clk) begin
      reg581 <= reg538;
      reg582 <= $unsigned((reg525 ? (+reg534) : (~reg573[(1'h0):(1'h0)])));
    end
  always
    @(posedge clk) begin
      reg583 <= (|forvar556);
      for (forvar584 = (1'h0); (forvar584 < (2'h3)); forvar584 = (forvar584 + (1'h1)))
        begin
          reg585 <= $unsigned(($signed((reg518 <= (8'hb9))) ?
              ("HCScrG3yI7E2" ?
                  (8'hbe) : $signed($unsigned(reg549))) : $signed(reg541[(2'h3):(1'h0)])));
          reg586 <= $unsigned("yaXn883ExcQr");
          reg587 = "I0mT9B";
          reg588 = (~^$signed($unsigned($signed((8'ha9)))));
          reg589 <= "qPGaNVQUG0k";
          reg590 <= $unsigned(reg577[(2'h3):(2'h2)]);
        end
      reg591 <= (reg532 ?
          $signed((forvar555 | ((reg529 ?
              forvar514 : reg516) >= "CFtaPJfNEYWbTqNQZDyA"))) : "z8Ece1MSaF");
    end
  assign wire592 = forvar519;
  assign wire593 = "88";
  assign wire594 = {{"WdS9zq", (+$unsigned($signed(reg589)))}};
  always
    @(posedge clk) begin
      reg595 <= (~^({reg500[(2'h2):(1'h0)]} ?
          ((&$unsigned(forvar568)) >> $signed($unsigned(reg587))) : $signed("44YDGGsCfxFyVq4")));
      if ("seeCP")
        begin
          reg596 <= (($unsigned((reg571 ?
                  reg543[(3'h4):(1'h1)] : wire496)) >>> (((~^forvar531) ?
                  (forvar501 ?
                      wire494 : reg522) : (reg545 ^ reg539)) ~^ {{reg532},
                  "myRfTGylkp"})) ?
              ((~&(|$unsigned(reg573))) ~^ $unsigned("VDHOEZIFK")) : reg563);
        end
      else
        begin
          reg596 = $signed(wire496);
        end
      reg597 <= (8'ha6);
      reg598 <= reg597[(1'h1):(1'h0)];
      if ($signed($unsigned((wire580 || $signed(reg563)))))
        begin
          reg599 <= $signed($signed(reg513));
          reg600 <= "HdIOgDGd6u";
          reg601 <= forvar560;
          reg602 <= (({reg500} ?
                  {(~&reg576[(4'he):(4'he)])} : "0khwDOX866WMgI5E1") ?
              forvar501 : $unsigned($signed(($signed(reg570) > $unsigned(reg596)))));
          reg603 <= $unsigned((wire594 == $signed(((8'ha5) ?
              reg567 : wire594[(2'h2):(1'h0)]))));
          reg604 <= $unsigned(wire511);
        end
      else
        begin
          reg599 <= reg591[(2'h3):(2'h3)];
          reg600 <= {((^reg500[(3'h4):(1'h0)]) ^~ reg538)};
        end
    end
  assign wire605 = forvar556;
  assign wire606 = (|$unsigned(reg550));
  always
    @(posedge clk) begin
      reg607 <= reg500[(2'h3):(1'h1)];
      reg608 <= (!{$signed($unsigned(reg515)), "StdPKaayzlbibyw"});
      for (forvar609 = (1'h0); (forvar609 < (2'h2)); forvar609 = (forvar609 + (1'h1)))
        begin
          reg610 = $unsigned((reg564 ? "xKBYToarfL2fU0v9dcaXulo" : reg509));
          reg611 <= ($unsigned({$unsigned((~&reg517)),
                  ("A4CuTxvu" ? $signed(forvar519) : {(8'ha0)})}) ?
              $unsigned(((|$unsigned((8'ha6))) * reg572[(3'h5):(3'h5)])) : (reg558[(2'h2):(1'h0)] ?
                  ($unsigned(reg603[(3'h7):(3'h6)]) != ((^reg586) ?
                      {reg547} : (8'hb7))) : "4VkCfJ8"));
        end
      reg612 = (!forvar519[(3'h7):(2'h2)]);
      reg613 <= ($unsigned("5p") >> $unsigned((+($unsigned(wire493) >> ""))));
      reg614 <= "e3";
    end
  always
    @(posedge clk) begin
      for (forvar615 = (1'h0); (forvar615 < (3'h5)); forvar615 = (forvar615 + (1'h1)))
        begin
          reg616 <= $unsigned((7'h43));
          reg617 <= "zPVWizdDOaa2DB0S";
          reg618 <= ($signed((~|((reg498 ? (8'h9c) : reg586) ?
                  $unsigned(reg572) : "C2O6zZNVNHVShhTxTehA0N8dT"))) ?
              reg561[(1'h0):(1'h0)] : reg540);
          for (forvar619 = (1'h0); (forvar619 < (2'h2)); forvar619 = (forvar619 + (1'h1)))
            begin
              reg620 <= ((8'hb2) >= (~&reg562));
              reg621 = forvar554[(1'h1):(1'h0)];
              reg622 <= (8'hb3);
            end
        end
    end
  assign wire623 = forvar542;
  always
    @(posedge clk) begin
      reg624 <= forvar542[(3'h7):(1'h0)];
      for (forvar625 = (1'h0); (forvar625 < (2'h3)); forvar625 = (forvar625 + (1'h1)))
        begin
          reg626 <= ((!$signed(($unsigned((8'hb3)) ?
              $unsigned(reg613) : $unsigned(reg578)))) == forvar535);
          reg627 = "NH0v";
          reg628 <= reg590[(3'h6):(3'h5)];
          reg629 <= $signed((~^{$signed($unsigned(reg550)),
              ($unsigned(forvar514) + {reg497})}));
          reg630 <= reg621;
          reg631 <= reg538[(1'h1):(1'h1)];
        end
    end
  always
    @(posedge clk) begin
      reg632 <= ((reg528[(2'h3):(1'h1)] ?
          $unsigned((^~$unsigned(reg576))) : ((~^(reg570 << reg544)) | "I1wCJUbD2")) >> (!$unsigned(($signed((7'h45)) || $signed(reg550)))));
    end
  always
    @(posedge clk) begin
      reg633 <= ($signed(wire574) >> reg587);
      reg634 <= $signed($signed(reg595[(1'h1):(1'h0)]));
      reg635 <= ((reg530 ?
          (($signed(reg630) + reg561[(5'h13):(4'he)]) >= $unsigned("5SR7fMVKtaKG")) : $unsigned($signed($signed(forvar514)))) | reg585);
      reg636 = (~reg533);
      reg637 <= (($unsigned($unsigned($signed(reg573))) ?
              ((!"vFeXl7BTppNqNO7MC") ?
                  "TAP" : (|(reg617 ?
                      wire592 : reg541))) : (^~$signed(reg630[(3'h7):(3'h7)]))) ?
          reg561 : ((+"EKw9mQetyQNE4") ?
              (reg622 ?
                  $signed((&(8'hab))) : reg585[(2'h2):(1'h0)]) : $signed(reg499[(1'h1):(1'h1)])));
      reg638 = $signed(wire605);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module435  (y, clk, wire439, wire438, wire437, wire436);
  output wire [(32'h2eb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire439;
  input wire [(4'hf):(1'h0)] wire438;
  input wire signed [(2'h3):(1'h0)] wire437;
  input wire [(3'h5):(1'h0)] wire436;
  reg signed [(5'h18):(1'h0)] reg488 = (1'h0);
  reg [(3'h5):(1'h0)] reg487 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg486 = (1'h0);
  reg [(4'hd):(1'h0)] reg485 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg484 = (1'h0);
  reg [(5'h16):(1'h0)] forvar483 = (1'h0);
  reg [(5'h1a):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg481 = (1'h0);
  reg [(4'ha):(1'h0)] reg480 = (1'h0);
  reg [(5'h17):(1'h0)] reg479 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg477 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg476 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar475 = (1'h0);
  reg [(5'h19):(1'h0)] forvar474 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg473 = (1'h0);
  reg [(3'h4):(1'h0)] reg472 = (1'h0);
  reg [(4'hf):(1'h0)] reg471 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg470 = (1'h0);
  reg [(4'h9):(1'h0)] forvar469 = (1'h0);
  reg [(4'hb):(1'h0)] reg468 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire467;
  wire [(2'h3):(1'h0)] wire466;
  reg [(4'hc):(1'h0)] reg465 = (1'h0);
  reg [(3'h5):(1'h0)] reg464 = (1'h0);
  wire [(5'h14):(1'h0)] wire463;
  wire signed [(4'h9):(1'h0)] wire462;
  reg signed [(3'h7):(1'h0)] reg461 = (1'h0);
  reg [(5'h11):(1'h0)] reg460 = (1'h0);
  reg [(5'h15):(1'h0)] reg459 = (1'h0);
  reg [(5'h18):(1'h0)] reg458 = (1'h0);
  reg [(5'h17):(1'h0)] reg457 = (1'h0);
  reg [(4'h9):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg455 = (1'h0);
  wire [(5'h13):(1'h0)] wire454;
  reg [(5'h17):(1'h0)] reg453 = (1'h0);
  reg [(4'hb):(1'h0)] reg452 = (1'h0);
  reg [(3'h6):(1'h0)] reg451 = (1'h0);
  reg [(5'h19):(1'h0)] reg450 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg447 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg446 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar445 = (1'h0);
  reg [(5'h19):(1'h0)] reg444 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg443 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg442 = (1'h0);
  reg [(4'hd):(1'h0)] reg441 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg440 = (1'h0);
  assign y = {reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 forvar483,
                 reg482,
                 reg481,
                 reg480,
                 reg479,
                 reg478,
                 reg477,
                 reg476,
                 forvar475,
                 forvar474,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 forvar469,
                 reg468,
                 wire467,
                 wire466,
                 reg465,
                 reg464,
                 wire463,
                 wire462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 wire454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 reg447,
                 reg446,
                 forvar445,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg440 <= (wire436 >= "");
      reg441 = wire437[(2'h3):(1'h1)];
      reg442 <= $signed(wire439);
      reg443 = ("PnyK51LFx2XFBGl3DAaBX5l1" < {(^{$unsigned(wire437),
              (reg440 << wire437)})});
      reg444 = $signed($unsigned($signed(wire439[(1'h1):(1'h1)])));
      for (forvar445 = (1'h0); (forvar445 < (3'h4)); forvar445 = (forvar445 + (1'h1)))
        begin
          reg446 <= ((^$unsigned(reg442)) <<< {"5KWpuvcf2qp2kc2GRkfeAJf",
              (reg442 ?
                  reg443[(3'h5):(3'h4)] : {(reg442 ? reg441 : wire438),
                      reg440[(1'h1):(1'h0)]})});
          reg447 <= ((("LSm" > reg440[(4'ha):(3'h6)]) < $signed("RN3ISRDOd0UFHkdv")) + $unsigned($unsigned(forvar445)));
          reg448 <= (wire438 ?
              wire437[(1'h0):(1'h0)] : (wire437[(2'h3):(1'h1)] ?
                  {{{(8'ha6), wire439}}} : (7'h4e)));
          reg449 <= wire437;
          reg450 <= reg441[(4'h8):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      reg451 <= (~&"yCt");
      reg452 <= (reg447[(5'h12):(2'h3)] & (~{(^((8'hb1) && wire437)),
          $unsigned("mvkD811HJ")}));
      reg453 <= ((&($signed("ez8ISBesmvqScSWr") ?
          ($unsigned(reg450) ?
              wire439[(1'h0):(1'h0)] : "e8FgbwNY") : (^~$signed(wire436)))) < forvar445);
    end
  assign wire454 = reg452;
  always
    @(posedge clk) begin
      reg455 <= {$signed(reg446), $unsigned(reg446)};
    end
  always
    @(posedge clk) begin
      reg456 <= wire436[(1'h1):(1'h0)];
      reg457 <= $unsigned($unsigned(reg441[(4'ha):(2'h2)]));
      reg458 = (forvar445 ? "BFc1tKDAMeFZeU" : $unsigned("TMKd1s8g3SNTvx6"));
      reg459 = $unsigned(reg458[(3'h5):(3'h5)]);
      reg460 <= reg450[(5'h10):(4'ha)];
      reg461 = (wire436[(1'h0):(1'h0)] <= wire439);
    end
  assign wire462 = $signed((((^{reg443,
                           (8'ha8)}) >> "PZbMWLLVlbFKRvHD4MKVwhRD") ?
                       $unsigned(reg452[(4'hb):(3'h7)]) : $unsigned(("w4aOIRxhyqs" ~^ $unsigned(wire454)))));
  assign wire463 = $signed($signed(($unsigned((reg458 ^~ reg444)) && (&wire462[(3'h7):(3'h6)]))));
  always
    @(posedge clk) begin
      reg464 <= $unsigned({($unsigned($signed((7'h44))) || "13xCnZuJVnVbr50T6qhpU7"),
          (($unsigned(reg452) <<< (reg449 ?
              wire462 : wire436)) + $signed((|reg459)))});
      reg465 <= {(($unsigned($unsigned(wire439)) ?
              "Y2ZOYIytUBOy1lhA" : (|(wire462 <<< reg449))) <<< forvar445),
          (reg455[(4'hf):(4'h9)] ? reg440[(2'h2):(2'h2)] : reg464)};
    end
  assign wire466 = reg451[(2'h3):(2'h3)];
  assign wire467 = reg450;
  always
    @(posedge clk) begin
      if ((^$unsigned("12KmQ3AB3Z")))
        begin
          reg468 = $signed(wire437[(1'h0):(1'h0)]);
        end
      else
        begin
          reg468 <= (|$unsigned($signed("D7nk")));
        end
      for (forvar469 = (1'h0); (forvar469 < (1'h1)); forvar469 = (forvar469 + (1'h1)))
        begin
          reg470 <= "";
          reg471 <= reg441[(2'h2):(2'h2)];
          reg472 <= (reg460 ?
              $signed((reg440 || $signed(reg448))) : wire466[(2'h2):(1'h1)]);
          reg473 = (8'hb8);
          for (forvar474 = (1'h0); (forvar474 < (3'h4)); forvar474 = (forvar474 + (1'h1)))
            begin
              for (forvar475 = (1'h0); (forvar475 < (1'h0)); forvar475 = (forvar475 + (1'h1)))
                begin
                  reg476 <= "dmKQII6lO";
                  reg477 <= $signed((~&$unsigned({{reg472},
                      $unsigned(reg447)})));
                  reg478 = wire437;
                  reg479 <= ({(-(wire438 == (reg472 <= reg452)))} ?
                      $unsigned($signed((~&(8'hb0)))) : reg476);
                  reg480 <= "ffLCbinV";
                  reg481 <= reg442[(2'h3):(1'h0)];
                end
              reg482 <= (~|(+"lKZQlT3IkpQ9g7"));
              for (forvar483 = (1'h0); (forvar483 < (2'h2)); forvar483 = (forvar483 + (1'h1)))
                begin
                  reg484 <= {$signed("ZZ"), $signed(reg472)};
                end
              reg485 <= wire437[(2'h3):(2'h3)];
              reg486 <= $signed($unsigned((($signed(reg443) ?
                  (reg484 << forvar469) : (~&wire436)) ^ "XJKLwJBvhHa5tXem")));
            end
          reg487 = "S";
        end
      reg488 <= forvar483[(4'hc):(4'ha)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module224
#(parameter param404 = {(|{(^~(+(8'hb9)))})}, parameter param405 = param404)
(y, clk, wire228, wire227, wire226, wire225);
  output wire [(32'h9dd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire228;
  input wire signed [(5'h11):(1'h0)] wire227;
  input wire [(5'h13):(1'h0)] wire226;
  input wire signed [(5'h10):(1'h0)] wire225;
  reg [(5'h18):(1'h0)] reg403 = (1'h0);
  reg [(3'h6):(1'h0)] reg402 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg401 = (1'h0);
  reg [(4'hf):(1'h0)] reg400 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg399 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg398 = (1'h0);
  wire [(5'h15):(1'h0)] wire397;
  wire [(5'h17):(1'h0)] wire396;
  wire [(5'h1a):(1'h0)] wire395;
  reg [(3'h5):(1'h0)] reg391 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg394 = (1'h0);
  reg [(5'h11):(1'h0)] reg393 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg392 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar391 = (1'h0);
  reg [(5'h10):(1'h0)] reg390 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg389 = (1'h0);
  reg [(3'h4):(1'h0)] reg388 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg387 = (1'h0);
  reg [(5'h1a):(1'h0)] reg386 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg385 = (1'h0);
  reg [(4'hf):(1'h0)] reg384 = (1'h0);
  reg [(5'h19):(1'h0)] reg383 = (1'h0);
  reg [(3'h7):(1'h0)] reg382 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg381 = (1'h0);
  reg [(3'h6):(1'h0)] reg380 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg378 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg377 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg376 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg375 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar374 = (1'h0);
  reg [(2'h3):(1'h0)] forvar373 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg372 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg371 = (1'h0);
  reg [(2'h2):(1'h0)] reg370 = (1'h0);
  reg [(5'h13):(1'h0)] forvar369 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg368 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg366 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg365 = (1'h0);
  reg [(2'h3):(1'h0)] reg364 = (1'h0);
  wire [(5'h11):(1'h0)] wire363;
  reg [(5'h17):(1'h0)] reg362 = (1'h0);
  reg [(3'h6):(1'h0)] reg361 = (1'h0);
  reg [(3'h6):(1'h0)] forvar360 = (1'h0);
  reg [(4'hc):(1'h0)] reg359 = (1'h0);
  reg [(4'he):(1'h0)] reg358 = (1'h0);
  reg [(5'h17):(1'h0)] reg357 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg356 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg355 = (1'h0);
  reg [(2'h2):(1'h0)] forvar354 = (1'h0);
  reg [(5'h15):(1'h0)] reg353 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg352 = (1'h0);
  reg [(3'h4):(1'h0)] forvar351 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg350 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg349 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg348 = (1'h0);
  reg [(3'h6):(1'h0)] reg347 = (1'h0);
  reg [(5'h16):(1'h0)] reg346 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg345 = (1'h0);
  reg [(4'he):(1'h0)] reg344 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg343 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg342 = (1'h0);
  reg [(5'h19):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg340 = (1'h0);
  reg [(2'h3):(1'h0)] forvar339 = (1'h0);
  reg [(4'ha):(1'h0)] reg338 = (1'h0);
  reg [(4'hd):(1'h0)] reg337 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar336 = (1'h0);
  reg [(2'h2):(1'h0)] forvar335 = (1'h0);
  reg [(5'h11):(1'h0)] reg334 = (1'h0);
  reg [(5'h11):(1'h0)] reg333 = (1'h0);
  wire [(5'h15):(1'h0)] wire332;
  reg signed [(2'h2):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg330 = (1'h0);
  reg [(4'hc):(1'h0)] reg329 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg327 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar325 = (1'h0);
  reg [(4'hc):(1'h0)] forvar323 = (1'h0);
  reg [(5'h17):(1'h0)] reg321 = (1'h0);
  reg [(4'hf):(1'h0)] reg320 = (1'h0);
  reg [(4'hc):(1'h0)] reg326 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg325 = (1'h0);
  reg [(5'h16):(1'h0)] reg324 = (1'h0);
  reg [(5'h11):(1'h0)] reg323 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg322 = (1'h0);
  reg [(3'h7):(1'h0)] forvar321 = (1'h0);
  reg [(5'h14):(1'h0)] forvar320 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg319 = (1'h0);
  reg [(5'h16):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg317 = (1'h0);
  reg [(4'hd):(1'h0)] reg316 = (1'h0);
  reg [(5'h12):(1'h0)] reg315 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg314 = (1'h0);
  reg [(4'hb):(1'h0)] reg313 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar311 = (1'h0);
  reg [(5'h13):(1'h0)] reg310 = (1'h0);
  reg [(4'hb):(1'h0)] forvar309 = (1'h0);
  reg [(4'h9):(1'h0)] reg308 = (1'h0);
  reg [(5'h19):(1'h0)] reg307 = (1'h0);
  reg [(5'h14):(1'h0)] reg306 = (1'h0);
  reg [(4'hc):(1'h0)] reg305 = (1'h0);
  reg [(5'h10):(1'h0)] reg304 = (1'h0);
  reg [(5'h10):(1'h0)] forvar303 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg302 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar301 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg300 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar299 = (1'h0);
  reg [(3'h7):(1'h0)] reg298 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg297 = (1'h0);
  reg [(4'he):(1'h0)] forvar296 = (1'h0);
  reg [(4'ha):(1'h0)] reg295 = (1'h0);
  reg [(2'h2):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg293 = (1'h0);
  reg [(3'h6):(1'h0)] reg292 = (1'h0);
  reg [(4'hd):(1'h0)] reg291 = (1'h0);
  reg [(5'h19):(1'h0)] reg290 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg289 = (1'h0);
  reg [(5'h19):(1'h0)] reg288 = (1'h0);
  reg [(5'h11):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar286 = (1'h0);
  reg [(5'h19):(1'h0)] forvar285 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg284 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg283 = (1'h0);
  reg [(3'h4):(1'h0)] reg282 = (1'h0);
  reg [(4'hd):(1'h0)] reg281 = (1'h0);
  reg [(5'h19):(1'h0)] reg280 = (1'h0);
  reg [(4'h9):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg278 = (1'h0);
  reg [(3'h6):(1'h0)] reg277 = (1'h0);
  reg [(4'hc):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg275 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg274 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg273 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar272 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg271 = (1'h0);
  reg [(4'hf):(1'h0)] forvar270 = (1'h0);
  reg [(5'h11):(1'h0)] forvar269 = (1'h0);
  wire [(4'h9):(1'h0)] wire268;
  wire signed [(4'h9):(1'h0)] wire267;
  reg signed [(4'hd):(1'h0)] reg266 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg265 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire264;
  reg signed [(3'h4):(1'h0)] reg263 = (1'h0);
  reg [(5'h1a):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg261 = (1'h0);
  reg [(5'h17):(1'h0)] forvar260 = (1'h0);
  reg [(4'hc):(1'h0)] reg259 = (1'h0);
  reg [(4'hf):(1'h0)] reg258 = (1'h0);
  reg [(5'h18):(1'h0)] reg257 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg255 = (1'h0);
  reg [(5'h14):(1'h0)] reg254 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar252 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg251 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg250 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg249 = (1'h0);
  reg [(5'h17):(1'h0)] reg248 = (1'h0);
  reg [(4'h9):(1'h0)] reg247 = (1'h0);
  reg [(5'h15):(1'h0)] reg246 = (1'h0);
  reg [(5'h19):(1'h0)] reg245 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg244 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg243 = (1'h0);
  reg [(3'h4):(1'h0)] reg242 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg241 = (1'h0);
  reg signed [(4'he):(1'h0)] reg240 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg239 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar238 = (1'h0);
  reg [(4'he):(1'h0)] forvar237 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg236 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg235 = (1'h0);
  reg [(5'h13):(1'h0)] reg234 = (1'h0);
  reg [(4'h9):(1'h0)] reg233 = (1'h0);
  reg [(5'h10):(1'h0)] forvar232 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg230 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg229 = (1'h0);
  assign y = {reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 wire397,
                 wire396,
                 wire395,
                 reg391,
                 reg394,
                 reg393,
                 reg392,
                 forvar391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 forvar374,
                 forvar373,
                 reg372,
                 reg371,
                 reg370,
                 forvar369,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 wire363,
                 reg362,
                 reg361,
                 forvar360,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 forvar354,
                 reg353,
                 reg352,
                 forvar351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 forvar339,
                 reg338,
                 reg337,
                 forvar336,
                 forvar335,
                 reg334,
                 reg333,
                 wire332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 forvar325,
                 forvar323,
                 reg321,
                 reg320,
                 reg326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 forvar321,
                 forvar320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 forvar311,
                 reg310,
                 forvar309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 forvar303,
                 reg302,
                 forvar301,
                 reg300,
                 forvar299,
                 reg298,
                 reg297,
                 forvar296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 forvar286,
                 forvar285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 forvar272,
                 reg271,
                 forvar270,
                 forvar269,
                 wire268,
                 wire267,
                 reg266,
                 reg265,
                 wire264,
                 reg263,
                 reg262,
                 reg261,
                 forvar260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 forvar252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 forvar238,
                 forvar237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 forvar232,
                 reg231,
                 reg230,
                 reg229,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg229 <= wire227;
      reg230 = $signed(wire227[(5'h11):(4'hc)]);
      reg231 <= $signed(reg230[(1'h1):(1'h1)]);
      for (forvar232 = (1'h0); (forvar232 < (3'h5)); forvar232 = (forvar232 + (1'h1)))
        begin
          reg233 <= (~$unsigned((wire225[(4'hc):(4'hb)] ?
              ({reg231} & wire226[(4'ha):(1'h0)]) : (^$signed(reg231)))));
          reg234 <= wire228[(1'h1):(1'h0)];
          reg235 <= forvar232[(4'hb):(4'hb)];
          reg236 = {(reg231 || $signed((wire228[(3'h5):(3'h5)] ?
                  (reg231 ? reg233 : wire226) : (wire227 & reg235))))};
          for (forvar237 = (1'h0); (forvar237 < (1'h1)); forvar237 = (forvar237 + (1'h1)))
            begin
              for (forvar238 = (1'h0); (forvar238 < (2'h2)); forvar238 = (forvar238 + (1'h1)))
                begin
                  reg239 <= $signed($signed((~^(8'hbe))));
                end
              reg240 <= $signed($signed(reg239));
              reg241 <= {reg236[(2'h2):(1'h0)],
                  ("iTnnF" <= (((reg236 && wire225) != (reg239 ?
                          reg233 : wire226)) ?
                      ((|wire227) | (reg229 ?
                          reg230 : forvar238)) : ($signed(wire228) ?
                          "2nJ5IWvYdIKN821anbpuDw39" : (!wire228))))};
              if ($unsigned($unsigned(wire227)))
                begin
                  reg242 <= $signed($signed(forvar232));
                  reg243 <= (~$unsigned($unsigned({(reg242 ?
                          reg230 : reg241)})));
                  reg244 <= reg240[(2'h2):(2'h2)];
                  reg245 <= ("kB" > ($signed((reg240 ?
                          $signed(wire227) : reg231[(2'h2):(1'h1)])) ?
                      (reg242 ?
                          ($signed(wire226) ?
                              (reg234 >= reg231) : (wire228 <= wire225)) : reg242) : ""));
                end
              else
                begin
                  reg242 <= $signed((~reg231));
                  reg243 <= $unsigned(wire228);
                  reg244 <= (wire225[(5'h10):(5'h10)] == reg241);
                  reg245 = {reg233};
                end
              reg246 <= $unsigned($signed((("3Ri" >= $unsigned(reg243)) ?
                  $unsigned($signed(reg240)) : ($signed(reg233) - {reg236}))));
            end
          reg247 <= reg229[(2'h2):(1'h1)];
        end
    end
  always
    @(posedge clk) begin
      reg248 <= (reg229 + (^~({(reg243 ? reg233 : reg241), "keNfR7gpvDY"} ?
          (~^$unsigned(wire227)) : {"xHGX80wepT6K6FkbbTk1",
              (reg229 ? reg243 : wire225)})));
    end
  always
    @(posedge clk) begin
      reg249 <= $signed($signed((reg242[(1'h1):(1'h0)] < ($unsigned(reg245) ?
          $signed(wire225) : $signed((8'ha9))))));
      reg250 <= ((reg249[(2'h3):(1'h0)] ?
          $signed(reg231) : reg248[(5'h11):(3'h5)]) && reg246);
      reg251 <= $signed(reg229);
    end
  always
    @(posedge clk) begin
      for (forvar252 = (1'h0); (forvar252 < (2'h3)); forvar252 = (forvar252 + (1'h1)))
        begin
          reg253 <= ($unsigned(reg233[(1'h1):(1'h0)]) ?
              forvar238[(5'h19):(2'h3)] : reg249);
          reg254 <= "C";
          reg255 = $signed({"Oa0BuWLhC4rxkoq"});
          reg256 <= $unsigned(((reg246 - (~|reg240[(3'h6):(2'h2)])) && (reg246[(4'ha):(3'h4)] ^~ ($unsigned(reg254) ?
              $signed(reg242) : reg243[(2'h2):(1'h0)]))));
        end
      reg257 <= {reg243[(2'h3):(1'h0)]};
      reg258 <= reg245[(1'h1):(1'h1)];
      reg259 <= $unsigned($unsigned($unsigned((reg236[(4'ha):(3'h6)] ?
          reg247[(3'h7):(3'h4)] : "pwUgP"))));
      for (forvar260 = (1'h0); (forvar260 < (3'h4)); forvar260 = (forvar260 + (1'h1)))
        begin
          reg261 <= reg251;
          reg262 <= "Sg42gZNQ18";
        end
      reg263 <= "8ybxRagk95gwt3V11VOtx";
    end
  assign wire264 = (($signed("PQciGYI6M6Zll7n") ?
                           (~($unsigned(reg236) ?
                               {forvar238,
                                   reg247} : (reg262 ^~ wire228))) : ($unsigned($signed(reg230)) ?
                               ((!forvar232) ?
                                   (reg231 ?
                                       reg242 : reg258) : (^reg243)) : reg254[(4'h8):(3'h7)])) ?
                       ("fFWmkPkvPc" == reg258[(4'hc):(2'h3)]) : reg255);
  always
    @(posedge clk) begin
      reg265 <= $unsigned(($signed(reg233) << $unsigned("2rf980NZB")));
      reg266 <= "NHdiUyRRKx387qINyvZLl";
    end
  assign wire267 = ($unsigned($signed((8'hba))) - (((^~(wire227 & reg254)) + reg261) ?
                       ($signed("IVEg06SWeJan5TAcqTR") ?
                           reg233 : (!(+reg245))) : (|(reg253 ?
                           (~^reg265) : $unsigned(reg234)))));
  assign wire268 = {$unsigned($unsigned(reg242))};
  always
    @(posedge clk) begin
      for (forvar269 = (1'h0); (forvar269 < (1'h0)); forvar269 = (forvar269 + (1'h1)))
        begin
          for (forvar270 = (1'h0); (forvar270 < (1'h1)); forvar270 = (forvar270 + (1'h1)))
            begin
              reg271 <= reg250;
              for (forvar272 = (1'h0); (forvar272 < (3'h4)); forvar272 = (forvar272 + (1'h1)))
                begin
                  reg273 <= reg248[(5'h12):(2'h3)];
                  reg274 <= ((~^$unsigned((+(|reg230)))) >> reg255[(4'hf):(4'hf)]);
                  reg275 = $unsigned(({"8vMXWWqIytn23h45YbHEv",
                          $signed((&(8'hba)))} ?
                      ((-(reg266 ?
                          wire228 : reg239)) <<< {reg233[(1'h0):(1'h0)],
                          wire226}) : (!$signed($unsigned(reg271)))));
                  reg276 <= (((reg265[(4'hf):(3'h6)] >>> ((~^wire264) ?
                              reg247 : (reg248 ? reg243 : forvar269))) ?
                          "VVJx09OUuebXKfW4tH" : $signed(wire225)) ?
                      {(-"4VFX1NDRo5RRVhFWhvKmHMt"),
                          (reg255 ?
                              ($signed(reg233) ?
                                  reg242 : reg233) : $signed(reg257))} : ("OE1Q5La0oyPAfa" <<< "OpO0KbtiNtyfGwvOg"));
                  reg277 = "R9eOFx4XvQCECe9";
                  reg278 <= $unsigned($signed((reg276[(3'h4):(3'h4)] ?
                      ($unsigned((8'ha2)) | (^~reg246)) : reg244[(3'h6):(3'h6)])));
                end
            end
          reg279 = (7'h4b);
          reg280 = (^(+$signed(reg253)));
          reg281 <= forvar237[(4'hb):(4'h8)];
          reg282 <= reg250;
        end
      reg283 <= {(|(~|((reg235 ? (8'ha0) : wire225) ?
              (^~reg247) : (wire268 ^ reg251)))),
          ($unsigned($unsigned(forvar270[(4'he):(4'he)])) ?
              ("8WS1IFt82v7tTQ2iJEJLG" ?
                  reg246 : {$signed(forvar238)}) : (~|(|forvar269)))};
      reg284 <= (reg239 < (("Ke5vh" ?
              ($unsigned((8'hbb)) ? "AS9" : $signed(reg255)) : (^~reg229)) ?
          $signed($unsigned(reg249)) : "IHiD7Ly3cBN9"));
    end
  always
    @(posedge clk) begin
      for (forvar285 = (1'h0); (forvar285 < (3'h4)); forvar285 = (forvar285 + (1'h1)))
        begin
          for (forvar286 = (1'h0); (forvar286 < (3'h5)); forvar286 = (forvar286 + (1'h1)))
            begin
              reg287 <= "MlrPs6t0yl00D7gYXf5LcS";
              reg288 <= reg242;
              reg289 = ((8'ha1) >> {{$unsigned($signed(reg239)),
                      forvar285[(5'h16):(3'h7)]}});
              reg290 <= reg257[(5'h16):(4'hf)];
            end
        end
      reg291 <= reg247;
      reg292 <= $unsigned("lemmmZT2SLzHFuS");
      reg293 = ($unsigned(forvar270[(3'h5):(1'h1)]) ?
          (-reg290) : ((-"WsbvIB") < reg229));
      reg294 = ($signed(forvar260[(4'hb):(3'h4)]) ?
          {"n",
              $unsigned(reg281[(4'hc):(1'h0)])} : {"ClEFbvfQxNue99J6mvOOOyLg"});
      reg295 <= reg265;
    end
  always
    @(posedge clk) begin
      for (forvar296 = (1'h0); (forvar296 < (1'h0)); forvar296 = (forvar296 + (1'h1)))
        begin
          reg297 <= {$signed((~{"fQ", (wire228 ? reg277 : reg274)}))};
          reg298 <= (^~reg236);
          for (forvar299 = (1'h0); (forvar299 < (1'h0)); forvar299 = (forvar299 + (1'h1)))
            begin
              reg300 = reg276;
              for (forvar301 = (1'h0); (forvar301 < (3'h5)); forvar301 = (forvar301 + (1'h1)))
                begin
                  reg302 <= (reg244[(1'h1):(1'h0)] | "6dBqdlNenPwRKUX11");
                end
            end
          for (forvar303 = (1'h0); (forvar303 < (2'h2)); forvar303 = (forvar303 + (1'h1)))
            begin
              if ((reg297[(3'h6):(1'h0)] ?
                  $signed(reg242[(3'h4):(2'h2)]) : $unsigned($signed(({reg239} == $signed((8'ha3)))))))
                begin
                  reg304 <= (reg263 || (((~|$unsigned(wire227)) ?
                      {(^~(7'h47)),
                          forvar303[(3'h5):(1'h0)]} : $unsigned((reg229 ?
                          reg276 : wire268))) < ({(8'hab)} ? (8'hb6) : "r")));
                end
              else
                begin
                  reg304 <= $signed((^~reg297));
                  reg305 <= (~&reg247[(1'h1):(1'h0)]);
                  reg306 <= (&wire226[(3'h7):(3'h7)]);
                  reg307 <= (reg244[(1'h1):(1'h0)] - wire228);
                  reg308 <= (~&{(&reg265[(4'hc):(3'h7)]), reg249});
                end
              for (forvar309 = (1'h0); (forvar309 < (2'h3)); forvar309 = (forvar309 + (1'h1)))
                begin
                  reg310 = reg297[(4'h9):(3'h6)];
                end
              for (forvar311 = (1'h0); (forvar311 < (3'h5)); forvar311 = (forvar311 + (1'h1)))
                begin
                  reg312 <= reg243;
                  reg313 <= (8'h9e);
                  reg314 <= (8'hb2);
                  reg315 <= reg305[(2'h2):(2'h2)];
                  reg316 = (~^(($signed((forvar286 & reg289)) ?
                      {$unsigned((8'hb5)),
                          reg295[(3'h6):(3'h4)]} : "E2qxWa") << reg234));
                  reg317 = $unsigned($unsigned(((+"h") && {reg235[(1'h0):(1'h0)]})));
                end
            end
        end
      if ($unsigned((8'hbe)))
        begin
          reg318 <= $unsigned(forvar296[(4'he):(1'h1)]);
          reg319 <= (reg315[(3'h5):(1'h0)] ?
              ({reg259} == reg305[(3'h4):(2'h3)]) : {{($unsigned(reg280) >>> $unsigned(wire268))}});
          for (forvar320 = (1'h0); (forvar320 < (1'h1)); forvar320 = (forvar320 + (1'h1)))
            begin
              for (forvar321 = (1'h0); (forvar321 < (2'h2)); forvar321 = (forvar321 + (1'h1)))
                begin
                  reg322 <= $signed("");
                  reg323 = $unsigned((|$unsigned(($signed(reg254) ^ $unsigned((8'hb5))))));
                  reg324 <= ("dDvHV9zASW" + (!(~|$unsigned($signed(reg253)))));
                end
              reg325 <= forvar252;
            end
          reg326 <= (~^(+$unsigned((8'ha9))));
        end
      else
        begin
          reg318 = ($signed(($signed((&reg262)) <<< $signed({reg281}))) ?
              (^(&($unsigned(reg255) && (!forvar238)))) : ((!("iQ1qUfl2rEGL" ?
                  "x5" : $unsigned(reg255))) == (reg245 ?
                  ({reg284} ?
                      reg276[(4'hc):(3'h4)] : "ebiO7klZ") : ((reg305 >= reg273) ^ "4TahYmSEJ2ognhnMTX"))));
          reg319 <= forvar321[(3'h4):(1'h1)];
          reg320 <= reg236;
          reg321 <= (forvar299[(2'h2):(1'h0)] ^~ forvar252[(5'h13):(1'h1)]);
          reg322 = ("bRCy9n2DP57pGXHK" ?
              $unsigned(($signed($signed((8'h9e))) ?
                  reg313[(4'ha):(1'h0)] : reg251)) : reg316[(3'h5):(3'h4)]);
          for (forvar323 = (1'h0); (forvar323 < (1'h0)); forvar323 = (forvar323 + (1'h1)))
            begin
              reg324 <= reg318;
              for (forvar325 = (1'h0); (forvar325 < (3'h4)); forvar325 = (forvar325 + (1'h1)))
                begin
                  reg326 <= $signed(($signed(((|reg249) ^~ $signed(reg323))) - ($unsigned(wire226[(1'h1):(1'h1)]) ^~ $unsigned(reg274[(2'h3):(2'h3)]))));
                  reg327 <= $signed($unsigned((~^reg250[(5'h11):(4'he)])));
                end
              reg328 = $unsigned($signed({(8'hbf)}));
              reg329 = ((~|"1QAQuaAVFXiDVtJO4PFol3") << reg323[(5'h10):(4'hb)]);
              reg330 <= ("oGnLB9CZPyqqAWQD0" ?
                  ("h4R6EiWpG" >> (8'hb7)) : $unsigned((8'ha5)));
              reg331 <= "";
            end
        end
    end
  assign wire332 = {$signed(reg229)};
  always
    @(posedge clk) begin
      reg333 <= (+(-(|{{reg290}, reg315[(4'ha):(3'h5)]})));
      reg334 <= (-forvar296);
      for (forvar335 = (1'h0); (forvar335 < (1'h1)); forvar335 = (forvar335 + (1'h1)))
        begin
          for (forvar336 = (1'h0); (forvar336 < (2'h2)); forvar336 = (forvar336 + (1'h1)))
            begin
              if (reg229[(1'h0):(1'h0)])
                begin
                  reg337 = $unsigned($signed(wire226));
                end
              else
                begin
                  reg337 <= reg244[(3'h5):(1'h0)];
                  reg338 <= $signed({"P6AitT",
                      (($unsigned(forvar238) + $signed(wire332)) ?
                          "CDao75pOpe3D" : ("0c2InmifAOyI" ?
                              (reg295 ~^ (8'ha4)) : "i47C7RSALBs71xIsDN7XVIyP"))});
                end
              for (forvar339 = (1'h0); (forvar339 < (1'h1)); forvar339 = (forvar339 + (1'h1)))
                begin
                  reg340 <= $unsigned((+$unsigned(forvar323)));
                  reg341 = $unsigned(("oH0IldvPxC" ?
                      $unsigned((|((8'hbf) ?
                          forvar285 : reg287))) : (((~&(8'ha5)) ?
                              (forvar311 ? reg261 : forvar320) : (~reg282)) ?
                          "Cc5gHoY5NSWCb04vIRdQ1T7F2" : reg230[(2'h3):(1'h0)])));
                  reg342 = "yCwpSAbdcUFJM1pkbJ";
                  reg343 <= {$unsigned($signed((forvar252[(5'h15):(3'h5)] ?
                          $unsigned(reg331) : $unsigned(reg246))))};
                  reg344 <= $unsigned($unsigned($unsigned(((reg277 != forvar321) ?
                      "OO2gWvgtaNAppa" : "omDECyswl7aZGLs4t0"))));
                  reg345 <= {$signed(reg290)};
                end
            end
          reg346 <= (reg318[(1'h1):(1'h0)] ?
              ("0CBDq6rkMXWyf21ys" * "cS") : $signed(($signed((^~reg300)) ?
                  $signed($unsigned(reg229)) : $signed("JPQIoAGJibs618pt2R3QVaXt"))));
          reg347 <= $unsigned(reg274);
          reg348 = $unsigned({(^~(^(reg343 ? reg277 : forvar325)))});
          reg349 <= reg318[(4'ha):(1'h0)];
        end
      reg350 <= (~reg349);
      for (forvar351 = (1'h0); (forvar351 < (2'h2)); forvar351 = (forvar351 + (1'h1)))
        begin
          reg352 <= reg320;
          reg353 = (^$unsigned(wire332[(4'ha):(3'h6)]));
          for (forvar354 = (1'h0); (forvar354 < (2'h2)); forvar354 = (forvar354 + (1'h1)))
            begin
              reg355 <= $signed((&(+$unsigned("he"))));
              reg356 = $unsigned((reg279[(2'h3):(2'h2)] + $unsigned({(~^(8'ha2))})));
            end
          reg357 <= $signed($unsigned(reg295[(4'h8):(3'h5)]));
        end
      reg358 <= $unsigned((^wire264));
    end
  always
    @(posedge clk) begin
      reg359 = ("nlxJz7dgh8evb2dEs1ka0RZzJ" - reg342);
      for (forvar360 = (1'h0); (forvar360 < (1'h1)); forvar360 = (forvar360 + (1'h1)))
        begin
          reg361 <= reg263;
          reg362 <= reg251[(3'h4):(1'h0)];
        end
    end
  assign wire363 = reg266[(4'h8):(3'h6)];
  always
    @(posedge clk) begin
      reg364 <= (&(~&{($unsigned(reg347) == (^~forvar311))}));
      reg365 <= "4bVOAZ";
    end
  always
    @(posedge clk) begin
      reg366 <= (~reg331);
      reg367 = (((~&(~^$unsigned(forvar260))) ^ (7'h47)) ?
          (reg245[(1'h1):(1'h0)] ?
              ($signed(reg362) ?
                  (reg231[(5'h10):(3'h4)] ?
                      reg236[(4'hb):(3'h6)] : {(7'h4d)}) : (8'ha2)) : reg346) : $signed("lS6plGtqNmp7IdR"));
      reg368 <= $signed(((|wire332[(1'h0):(1'h0)]) ?
          "kxlgO2cLektzkprRyk0YPDpBs" : (~&$signed(reg308))));
      for (forvar369 = (1'h0); (forvar369 < (3'h5)); forvar369 = (forvar369 + (1'h1)))
        begin
          reg370 = $unsigned((reg326[(1'h0):(1'h0)] + reg318[(4'h8):(4'h8)]));
          reg371 <= (|($unsigned((!(reg244 ? reg324 : (7'h4c)))) >> reg356));
          reg372 <= $unsigned((+(reg233[(2'h3):(2'h3)] & ("SmwHdNWYdoDAfKKaguxFM" != $signed(forvar325)))));
          for (forvar373 = (1'h0); (forvar373 < (3'h4)); forvar373 = (forvar373 + (1'h1)))
            begin
              for (forvar374 = (1'h0); (forvar374 < (2'h3)); forvar374 = (forvar374 + (1'h1)))
                begin
                  reg375 = "rPzbV";
                  reg376 <= (7'h45);
                  reg377 <= ((reg300 ?
                      ("XpQxIGqeQi" ?
                          (((8'hb7) ? reg361 : (8'ha4)) ?
                              reg371[(2'h2):(1'h1)] : reg275) : "sweMJAEg7iX2Yi43HsXp") : (8'hb4)) * ($unsigned("") ^~ reg258));
                  reg378 <= $signed((-reg320[(4'hc):(2'h3)]));
                  reg379 <= $unsigned((|$signed((~&(reg287 ?
                      forvar232 : reg370)))));
                  reg380 <= reg284[(4'hb):(4'h8)];
                end
              reg381 = (reg347 << (~^reg247));
              reg382 <= "tJPLQfaV";
              reg383 <= ("LitWh2D4iCn5Eq" > reg322);
              reg384 = ($signed((8'hb1)) >> $signed(((&(~|reg356)) <= {(forvar301 >= forvar237)})));
              reg385 <= $signed(("dmJ3gPpP8x3eM5Ypa" ?
                  reg355[(4'h9):(3'h4)] : {((reg283 ? forvar354 : forvar351) ?
                          "FZ0qzWyCBF" : $signed((8'haa)))}));
            end
        end
      reg386 <= {({forvar325[(4'hb):(3'h6)],
              ("eNvHSha2T7Fa2l6Mdd9U3WCUE" < (forvar323 > (7'h48)))} && {"BRMoQlmGuoeDwE6eZQ9KeXDa"}),
          "aBnw9wbKJcQCbJ78M9A"};
    end
  always
    @(posedge clk) begin
      reg387 <= $unsigned(("PR0hW6cbUShrd" & "FO6F845PbaHKzcH0466ncOBFc"));
    end
  always
    @(posedge clk) begin
      if ((|(reg283[(4'h9):(4'h9)] ?
          $unsigned(reg331[(1'h1):(1'h1)]) : {reg343,
              (wire226 != (reg310 >>> (8'hbf)))})))
        begin
          reg388 <= (((!{(forvar339 - reg254), $unsigned(reg287)}) ?
                  (+(reg297 ~^ (^~reg256))) : "uSeSawFLHeh") ?
              (8'hb5) : reg319[(1'h1):(1'h0)]);
          reg389 <= $unsigned(reg340);
          reg390 <= "VrT87nFsgEwxSp";
          for (forvar391 = (1'h0); (forvar391 < (1'h1)); forvar391 = (forvar391 + (1'h1)))
            begin
              reg392 <= (^(+reg280));
              reg393 <= $unsigned($unsigned($signed((^~$signed(reg387)))));
            end
          reg394 <= (^~forvar270);
        end
      else
        begin
          reg388 = "Z18NcwtmVlmQzu4JAeuLsaMS";
          reg389 <= (~|({$signed((forvar354 ? reg315 : reg308))} ?
              $signed(reg329) : reg255[(3'h7):(2'h3)]));
          reg390 = wire363;
          reg391 <= $unsigned((!$unsigned((reg297 < (8'hbd)))));
          reg392 <= forvar335;
          reg393 <= $signed($signed((-{(8'hbe)})));
        end
    end
  assign wire395 = forvar301;
  assign wire396 = reg381[(3'h6):(1'h0)];
  assign wire397 = (((~($unsigned(reg386) ? reg276 : reg259[(4'hc):(4'hb)])) ?
                           ({reg330} ?
                               (reg362 ?
                                   (wire267 >= (8'hac)) : reg337[(1'h1):(1'h1)]) : (forvar309[(2'h3):(2'h2)] && forvar252[(1'h0):(1'h0)])) : $unsigned("IxJZ")) ?
                       "CbU" : reg266);
  always
    @(posedge clk) begin
      reg398 <= (!$signed(reg312));
      reg399 <= $signed($unsigned($signed(($signed(reg393) < $signed(reg257)))));
      reg400 <= reg355;
      reg401 = ($signed(reg393[(3'h5):(3'h5)]) ?
          forvar301[(2'h2):(2'h2)] : (reg245 ?
              $unsigned(($unsigned(reg350) << forvar272)) : reg308[(4'h8):(1'h1)]));
      reg402 <= (reg257[(4'he):(3'h5)] + {$signed((7'h4b)),
          ({((7'h4a) || reg283), $signed(reg375)} << ("WB6TF9KOwKV9PMgS2iqxc" ?
              "9duSR0UeDRm" : "lqlemn0glHoIPuNQPIZPA2FL"))});
      reg403 <= reg393[(3'h4):(1'h0)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1753  (y, clk, wire1757, wire1756, wire1755, wire1754);
  output wire [(32'h9e7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h18):(1'h0)] wire1757;
  input wire [(4'h8):(1'h0)] wire1756;
  input wire signed [(5'h10):(1'h0)] wire1755;
  input wire [(4'h8):(1'h0)] wire1754;
  wire signed [(4'hc):(1'h0)] wire1931;
  reg signed [(2'h3):(1'h0)] reg1930 = (1'h0);
  wire [(5'h13):(1'h0)] wire1929;
  wire signed [(4'hc):(1'h0)] wire1928;
  wire signed [(5'h18):(1'h0)] wire1927;
  reg [(5'h14):(1'h0)] reg1926 = (1'h0);
  reg [(5'h11):(1'h0)] reg1925 = (1'h0);
  reg [(3'h4):(1'h0)] reg1922 = (1'h0);
  reg [(4'he):(1'h0)] forvar1920 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1915 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1914 = (1'h0);
  reg [(3'h6):(1'h0)] reg1924 = (1'h0);
  reg [(2'h3):(1'h0)] reg1923 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1922 = (1'h0);
  reg [(5'h14):(1'h0)] reg1921 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1920 = (1'h0);
  reg [(2'h2):(1'h0)] reg1919 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1918 = (1'h0);
  reg [(5'h17):(1'h0)] reg1917 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1916 = (1'h0);
  reg [(5'h17):(1'h0)] reg1915 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1914 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1913 = (1'h0);
  reg [(4'he):(1'h0)] reg1912 = (1'h0);
  reg [(5'h10):(1'h0)] reg1911 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1910 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1909 = (1'h0);
  reg [(4'he):(1'h0)] reg1908 = (1'h0);
  reg [(5'h15):(1'h0)] reg1907 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1906 = (1'h0);
  reg [(4'ha):(1'h0)] reg1905 = (1'h0);
  reg [(4'hf):(1'h0)] reg1904 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1903 = (1'h0);
  reg [(3'h7):(1'h0)] reg1902 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1901 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1900 = (1'h0);
  reg [(5'h16):(1'h0)] reg1899 = (1'h0);
  reg [(5'h15):(1'h0)] reg1898 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1897 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1896 = (1'h0);
  reg [(5'h13):(1'h0)] reg1895 = (1'h0);
  reg [(3'h7):(1'h0)] reg1894 = (1'h0);
  reg [(4'h9):(1'h0)] reg1893 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1892 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1891 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1890 = (1'h0);
  reg [(5'h10):(1'h0)] reg1889 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1888 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1887 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1886 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1885 = (1'h0);
  reg [(3'h7):(1'h0)] reg1884 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1883 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1882 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1881 = (1'h0);
  reg [(4'hd):(1'h0)] reg1880 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1879 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1878 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1877 = (1'h0);
  reg [(5'h19):(1'h0)] reg1876 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1875 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1874 = (1'h0);
  reg [(4'he):(1'h0)] forvar1873 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1872 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1871 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1870 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1869 = (1'h0);
  reg [(5'h17):(1'h0)] reg1868 = (1'h0);
  reg [(5'h14):(1'h0)] reg1867 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1866 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1865 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1864 = (1'h0);
  reg [(2'h3):(1'h0)] reg1863 = (1'h0);
  reg [(5'h19):(1'h0)] reg1862 = (1'h0);
  reg [(5'h18):(1'h0)] reg1861 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1860 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1859 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1858 = (1'h0);
  reg [(5'h12):(1'h0)] reg1857 = (1'h0);
  reg [(4'hd):(1'h0)] reg1856 = (1'h0);
  reg [(5'h13):(1'h0)] reg1855 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1854 = (1'h0);
  reg [(5'h11):(1'h0)] reg1853 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1852 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1851 = (1'h0);
  reg [(5'h16):(1'h0)] reg1850 = (1'h0);
  reg [(4'hf):(1'h0)] reg1849 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1848 = (1'h0);
  reg [(5'h15):(1'h0)] reg1847 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1846 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1845 = (1'h0);
  wire [(5'h16):(1'h0)] wire1844;
  reg [(5'h18):(1'h0)] reg1843 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1842 = (1'h0);
  reg [(3'h7):(1'h0)] reg1841 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1840 = (1'h0);
  reg [(4'hc):(1'h0)] reg1839 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1838 = (1'h0);
  reg [(5'h16):(1'h0)] reg1837 = (1'h0);
  reg [(4'hf):(1'h0)] reg1836 = (1'h0);
  reg [(4'hc):(1'h0)] reg1835 = (1'h0);
  reg [(3'h7):(1'h0)] reg1834 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1833 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1832 = (1'h0);
  reg [(4'hf):(1'h0)] reg1831 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1830 = (1'h0);
  reg [(5'h11):(1'h0)] reg1829 = (1'h0);
  reg [(3'h6):(1'h0)] reg1828 = (1'h0);
  reg [(4'ha):(1'h0)] reg1827 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1826 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1825 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1824 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1823 = (1'h0);
  reg [(4'hf):(1'h0)] reg1822 = (1'h0);
  reg [(4'hd):(1'h0)] reg1821 = (1'h0);
  reg [(4'hf):(1'h0)] reg1820 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1819 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1818 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1817 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1816 = (1'h0);
  reg [(4'he):(1'h0)] forvar1815 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1814 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1813 = (1'h0);
  reg [(3'h7):(1'h0)] reg1812 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1811 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1810 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1809 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1808 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1807 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1806 = (1'h0);
  reg [(5'h11):(1'h0)] reg1805 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1804 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1803 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1802 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1801 = (1'h0);
  reg [(2'h3):(1'h0)] reg1800 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1799 = (1'h0);
  reg [(5'h15):(1'h0)] reg1798 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire1797;
  reg signed [(2'h2):(1'h0)] reg1796 = (1'h0);
  reg [(3'h6):(1'h0)] reg1795 = (1'h0);
  reg [(5'h19):(1'h0)] reg1794 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1793 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1792 = (1'h0);
  reg [(5'h19):(1'h0)] reg1791 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1790 = (1'h0);
  reg [(3'h4):(1'h0)] reg1789 = (1'h0);
  reg [(3'h6):(1'h0)] reg1788 = (1'h0);
  reg [(4'h8):(1'h0)] reg1787 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire1786;
  reg [(4'h8):(1'h0)] reg1785 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1784 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1783 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1782 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1781 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1780 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1779 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1778 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1777 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1776 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1775 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1774 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1773 = (1'h0);
  reg [(5'h11):(1'h0)] reg1772 = (1'h0);
  reg [(5'h18):(1'h0)] reg1771 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1770 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1769 = (1'h0);
  reg [(5'h15):(1'h0)] reg1768 = (1'h0);
  reg [(4'ha):(1'h0)] reg1767 = (1'h0);
  reg [(3'h4):(1'h0)] reg1766 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1765 = (1'h0);
  reg [(5'h17):(1'h0)] reg1764 = (1'h0);
  reg [(3'h6):(1'h0)] reg1763 = (1'h0);
  reg [(5'h16):(1'h0)] reg1762 = (1'h0);
  reg [(2'h3):(1'h0)] reg1761 = (1'h0);
  reg [(3'h4):(1'h0)] reg1760 = (1'h0);
  reg [(3'h6):(1'h0)] reg1759 = (1'h0);
  reg [(4'hc):(1'h0)] reg1758 = (1'h0);
  assign y = {wire1931,
                 reg1930,
                 wire1929,
                 wire1928,
                 wire1927,
                 reg1926,
                 reg1925,
                 reg1922,
                 forvar1920,
                 forvar1915,
                 reg1914,
                 reg1924,
                 reg1923,
                 forvar1922,
                 reg1921,
                 reg1920,
                 reg1919,
                 reg1918,
                 reg1917,
                 reg1916,
                 reg1915,
                 forvar1914,
                 reg1913,
                 reg1912,
                 reg1911,
                 reg1910,
                 forvar1909,
                 reg1908,
                 reg1907,
                 reg1906,
                 reg1905,
                 reg1904,
                 reg1903,
                 reg1902,
                 reg1901,
                 forvar1900,
                 reg1899,
                 reg1898,
                 reg1897,
                 reg1896,
                 reg1895,
                 reg1894,
                 reg1893,
                 reg1892,
                 forvar1891,
                 forvar1890,
                 reg1889,
                 reg1888,
                 forvar1887,
                 forvar1886,
                 reg1885,
                 reg1884,
                 reg1883,
                 reg1882,
                 reg1881,
                 reg1880,
                 forvar1879,
                 forvar1878,
                 reg1877,
                 reg1876,
                 reg1875,
                 reg1874,
                 forvar1873,
                 reg1872,
                 forvar1871,
                 forvar1870,
                 reg1869,
                 reg1868,
                 reg1867,
                 reg1866,
                 reg1865,
                 reg1864,
                 reg1863,
                 reg1862,
                 reg1861,
                 forvar1860,
                 reg1859,
                 reg1858,
                 reg1857,
                 reg1856,
                 reg1855,
                 reg1854,
                 reg1853,
                 reg1852,
                 forvar1851,
                 reg1850,
                 reg1849,
                 forvar1848,
                 reg1847,
                 reg1846,
                 reg1845,
                 wire1844,
                 reg1843,
                 reg1842,
                 reg1841,
                 reg1840,
                 reg1839,
                 reg1838,
                 reg1837,
                 reg1836,
                 reg1835,
                 reg1834,
                 reg1833,
                 reg1832,
                 reg1831,
                 reg1830,
                 reg1829,
                 reg1828,
                 reg1827,
                 forvar1826,
                 forvar1825,
                 reg1824,
                 reg1823,
                 reg1822,
                 reg1821,
                 reg1820,
                 reg1819,
                 reg1818,
                 reg1817,
                 reg1816,
                 forvar1815,
                 forvar1814,
                 reg1813,
                 reg1812,
                 reg1811,
                 reg1810,
                 reg1809,
                 reg1808,
                 forvar1807,
                 reg1806,
                 reg1805,
                 forvar1804,
                 reg1803,
                 forvar1802,
                 forvar1801,
                 reg1800,
                 reg1799,
                 reg1798,
                 wire1797,
                 reg1796,
                 reg1795,
                 reg1794,
                 reg1793,
                 reg1792,
                 reg1791,
                 reg1790,
                 reg1789,
                 reg1788,
                 reg1787,
                 wire1786,
                 reg1785,
                 reg1784,
                 reg1783,
                 reg1782,
                 reg1781,
                 reg1780,
                 reg1779,
                 reg1778,
                 reg1777,
                 reg1776,
                 reg1775,
                 forvar1774,
                 reg1773,
                 reg1772,
                 reg1771,
                 reg1770,
                 reg1769,
                 reg1768,
                 reg1767,
                 reg1766,
                 forvar1765,
                 reg1764,
                 reg1763,
                 reg1762,
                 reg1761,
                 reg1760,
                 reg1759,
                 reg1758,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1758 = wire1756;
      reg1759 <= wire1756[(4'h8):(2'h2)];
      reg1760 <= reg1758[(2'h3):(2'h2)];
      reg1761 <= ("xkM5pSDEAk7anEIWkyPCO5sD" <<< (^(^(!"SXr8NBi0J"))));
      reg1762 <= wire1755[(4'hd):(3'h6)];
    end
  always
    @(posedge clk) begin
      reg1763 <= ({$unsigned("p36FMqsk")} ? "BheL6gNXBbVB3" : "xiaW");
    end
  always
    @(posedge clk) begin
      reg1764 <= (~$unsigned((~&reg1763)));
      for (forvar1765 = (1'h0); (forvar1765 < (3'h5)); forvar1765 = (forvar1765 + (1'h1)))
        begin
          reg1766 = $unsigned("8EstBZUNga");
        end
      reg1767 <= $unsigned($unsigned({(reg1762[(5'h10):(4'ha)] ?
              $unsigned(reg1761) : "ntaCdEoUZTRcBDzmP3h"),
          $unsigned((-wire1757))}));
      reg1768 = "MHevPr7HX2pRNMN9TwoAD6A5f";
      reg1769 <= $unsigned(reg1764[(5'h16):(5'h16)]);
    end
  always
    @(posedge clk) begin
      reg1770 <= "A9Ev8cYOrQ3xtvD";
      reg1771 <= $unsigned(((({reg1760, reg1761} > reg1766) == (reg1759 ?
              forvar1765 : {(8'haa), reg1768})) ?
          (~&reg1763[(1'h0):(1'h0)]) : ($unsigned(reg1764) >>> $signed(reg1759[(2'h2):(1'h1)]))));
      reg1772 <= (&$signed($signed($signed($unsigned(reg1771)))));
      reg1773 = "muRDx";
    end
  always
    @(posedge clk) begin
      for (forvar1774 = (1'h0); (forvar1774 < (3'h5)); forvar1774 = (forvar1774 + (1'h1)))
        begin
          reg1775 <= $unsigned(forvar1774[(5'h15):(3'h6)]);
          reg1776 <= {$signed(($signed((~wire1755)) + $unsigned($signed(wire1754))))};
          reg1777 <= "gCwiYwfHVaJDP50Jlw";
          reg1778 <= (((!((reg1770 ?
                  (8'hbf) : reg1775) ^ $unsigned((8'hab)))) >>> "TXs3qqRA76GHQZDJ") ?
              ("LBJS4Am2RYAXuSfXb" ?
                  (("RhpVdGE3p1fmBZ" && "ayPFNcerZFmYhGO") ?
                      (forvar1774[(5'h16):(4'ha)] ?
                          (wire1756 + reg1766) : "EVgskB35aoFESo") : reg1775) : {forvar1774[(2'h3):(1'h1)]}) : (7'h4d));
        end
      reg1779 <= wire1756[(3'h7):(3'h4)];
    end
  always
    @(posedge clk) begin
      reg1780 <= wire1756;
      reg1781 <= $unsigned((((^~wire1756[(2'h3):(1'h0)]) <<< ($signed(wire1754) ?
              reg1764[(3'h4):(1'h0)] : "1Chw9L9a")) ?
          $signed("rgEJ") : (reg1772[(4'he):(3'h7)] ?
              reg1763[(3'h4):(2'h2)] : $signed($unsigned(reg1771)))));
      reg1782 = "FLdqS7XBPtNf132D0";
    end
  always
    @(posedge clk) begin
      reg1783 <= forvar1774;
      reg1784 <= reg1780[(3'h4):(3'h4)];
      reg1785 = "es7xtRqx4";
    end
  assign wire1786 = (|$unsigned((~&(|reg1785))));
  always
    @(posedge clk) begin
      reg1787 <= (("w" ?
              {{$signed(reg1781), wire1757},
                  reg1769[(4'hb):(3'h7)]} : "Vnr3M7eStZ8CU") ?
          {(+($unsigned((8'hab)) >>> $signed(reg1778)))} : "aF");
      reg1788 <= ("L2vXOVwv" ?
          reg1772[(4'hf):(4'hd)] : (reg1767[(2'h3):(2'h3)] ?
              reg1778 : $signed(($signed(reg1770) ? (&(8'ha5)) : reg1772))));
      reg1789 <= "IIUOqE4eE4eNG6BURuT";
      reg1790 = "2dDeMSZaIJKT";
    end
  always
    @(posedge clk) begin
      reg1791 = $unsigned((($unsigned(((8'hbd) || reg1762)) | "n5Xk0KRYlvR2eP") || (reg1782 - ($signed(reg1784) ?
          (reg1769 ? reg1773 : (7'h4e)) : "MWP0yipSiLzqJkBafUhMVa"))));
      reg1792 <= $signed(reg1791);
      reg1793 = reg1761;
      reg1794 <= forvar1774[(2'h2):(2'h2)];
      reg1795 <= ((8'hb1) ?
          $signed("OfcLGthoX9OzmB78OAsbYR") : (forvar1765 + {((reg1792 ?
                      reg1788 : reg1773) ?
                  (8'haa) : {(8'ha9), reg1763})}));
      reg1796 <= "JR";
    end
  assign wire1797 = (-{reg1781[(5'h15):(4'hd)],
                        ($signed("d0pVAT") && ($unsigned(reg1767) ?
                            (reg1792 ^ reg1788) : (+wire1755)))});
  always
    @(posedge clk) begin
      reg1798 <= {""};
      reg1799 <= "N7D";
    end
  always
    @(posedge clk) begin
      reg1800 <= reg1780[(3'h4):(3'h4)];
    end
  always
    @(posedge clk) begin
      for (forvar1801 = (1'h0); (forvar1801 < (3'h5)); forvar1801 = (forvar1801 + (1'h1)))
        begin
          for (forvar1802 = (1'h0); (forvar1802 < (3'h4)); forvar1802 = (forvar1802 + (1'h1)))
            begin
              reg1803 <= (reg1761[(2'h3):(1'h0)] | reg1785[(4'h8):(2'h3)]);
            end
          for (forvar1804 = (1'h0); (forvar1804 < (2'h3)); forvar1804 = (forvar1804 + (1'h1)))
            begin
              reg1805 <= ("mCnUMLEBd6DE40Id" & reg1768[(3'h6):(3'h4)]);
              reg1806 <= "yrw";
              for (forvar1807 = (1'h0); (forvar1807 < (3'h5)); forvar1807 = (forvar1807 + (1'h1)))
                begin
                  reg1808 <= ((reg1795[(2'h3):(1'h0)] | (~&($signed(reg1806) ?
                      $unsigned(reg1777) : $signed(forvar1765)))) >= reg1761);
                  reg1809 = reg1796;
                  reg1810 <= $unsigned($unsigned(($signed("wphTmgC1CQiHfMMlI") == $signed(reg1808))));
                  reg1811 <= ($signed((!($signed(reg1808) >>> forvar1802[(3'h4):(3'h4)]))) ?
                      (reg1810[(4'hc):(1'h1)] ?
                          $signed($signed("fk3")) : "pYrImNb0IFCcFmobSDD") : (^""));
                  reg1812 <= reg1768[(1'h0):(1'h0)];
                  reg1813 <= {$unsigned($unsigned($unsigned($unsigned(forvar1765))))};
                end
            end
          for (forvar1814 = (1'h0); (forvar1814 < (2'h2)); forvar1814 = (forvar1814 + (1'h1)))
            begin
              for (forvar1815 = (1'h0); (forvar1815 < (3'h5)); forvar1815 = (forvar1815 + (1'h1)))
                begin
                  reg1816 <= ((reg1785 ?
                          (~{forvar1774, reg1776}) : (($unsigned(reg1806) ?
                                  (reg1787 ?
                                      (8'ha5) : (8'hb6)) : (reg1779 ^ reg1781)) ?
                              "SU" : wire1756[(4'h8):(4'h8)])) ?
                      wire1757 : reg1794[(1'h0):(1'h0)]);
                  reg1817 <= ($signed(($signed(reg1799[(2'h3):(2'h2)]) ?
                          reg1803[(5'h13):(2'h2)] : (~(reg1799 ?
                              reg1760 : (8'ha4))))) ?
                      wire1786[(2'h3):(2'h2)] : (-reg1764[(5'h17):(5'h13)]));
                  reg1818 = wire1754[(1'h1):(1'h1)];
                  reg1819 = forvar1807[(4'hb):(3'h6)];
                  reg1820 = ($signed(reg1781) >= $signed("u"));
                end
            end
          reg1821 <= $signed("pNiGnO");
          reg1822 <= (~&(|reg1760[(2'h3):(2'h3)]));
        end
      reg1823 <= $signed(forvar1814);
      reg1824 = reg1761;
      for (forvar1825 = (1'h0); (forvar1825 < (2'h3)); forvar1825 = (forvar1825 + (1'h1)))
        begin
          for (forvar1826 = (1'h0); (forvar1826 < (1'h0)); forvar1826 = (forvar1826 + (1'h1)))
            begin
              reg1827 = reg1770;
              reg1828 = ((((^(reg1788 ? forvar1814 : reg1821)) ?
                      {reg1803[(5'h12):(4'hc)]} : ("NukaDJwIJkQCLfe7LzeoJ" == (reg1764 >>> (7'h41)))) ?
                  (&reg1775[(5'h16):(3'h5)]) : "kVTNqM") >= (~($signed(reg1806[(3'h5):(3'h5)]) != "HGGfA1uUzWayMAbU3g7x1H90o")));
              reg1829 <= reg1778[(3'h5):(1'h0)];
              reg1830 <= (7'h4c);
            end
          if (reg1806[(1'h0):(1'h0)])
            begin
              reg1831 = ("4zguNaiCsBxaw4tf32I3tNZ" < reg1760[(3'h4):(2'h2)]);
              reg1832 <= ($signed((wire1757 ?
                      ((forvar1774 >> reg1794) >> $signed(reg1775)) : ("akInz" ?
                          reg1828[(3'h4):(2'h2)] : reg1823[(5'h10):(4'he)]))) ?
                  ((+reg1778[(1'h0):(1'h0)]) ?
                      {$signed($signed(reg1823)),
                          wire1755} : (^forvar1801[(3'h5):(3'h4)])) : $signed($unsigned(reg1805)));
              reg1833 <= "yPJGOT";
              reg1834 = (-reg1813[(3'h4):(3'h4)]);
              reg1835 <= "9DJFW2";
            end
          else
            begin
              reg1831 = (^"aI8");
              reg1832 <= $unsigned((^(((reg1819 >= reg1792) ?
                      {forvar1801, forvar1765} : "bSBH2") ?
                  $unsigned("NbU3vHSWqd2nK4Pd") : ((!(8'hbb)) ?
                      forvar1807[(5'h11):(4'h8)] : (reg1817 + reg1775)))));
              reg1833 <= $unsigned(forvar1807[(1'h1):(1'h0)]);
              reg1834 = ((|reg1789) & (+"bROvPZm3vs"));
            end
          if (($unsigned({wire1786}) ?
              "kR5LUsCie4BLcKiP8G3kFDDH" : (({(^~reg1812)} ^~ $signed($signed(reg1766))) ?
                  reg1760 : $signed((reg1803 ?
                      reg1779 : $unsigned(forvar1807))))))
            begin
              reg1836 <= $unsigned(($signed($unsigned("0lY9LTvoXrlZhnCIJVkeW0f")) << reg1818[(1'h1):(1'h0)]));
              reg1837 <= $signed((+reg1767[(3'h6):(1'h0)]));
            end
          else
            begin
              reg1836 <= (!reg1773);
              reg1837 <= reg1791;
              reg1838 <= $unsigned($unsigned($signed("nhIi2A337VcsE2gc4J")));
              reg1839 <= $signed((reg1792 ?
                  {($unsigned((8'ha3)) ? reg1827[(4'ha):(3'h5)] : reg1776),
                      $unsigned($signed(reg1758))} : reg1784));
              reg1840 <= forvar1815[(2'h2):(1'h0)];
            end
          reg1841 <= (~&reg1771);
          reg1842 <= ((reg1772[(1'h0):(1'h0)] ?
                  ($unsigned(reg1790) + "VYS0y5") : forvar1774) ?
              ((((reg1772 ? reg1823 : reg1818) ? (~^reg1837) : {reg1827}) ?
                  ((reg1787 ^ reg1784) ?
                      (8'ha4) : "gz") : {reg1829[(3'h4):(3'h4)],
                      "RB9kvaiRAA7R"}) << reg1798[(3'h4):(1'h1)]) : "eCp2ZHlbdIXrYkup4");
          reg1843 <= $signed(reg1830);
        end
    end
  assign wire1844 = $signed(((+($unsigned(reg1817) ~^ reg1835)) ?
                        $signed("12n05x76JMW8J9nMmIS6") : (($unsigned(reg1788) ~^ (reg1823 ?
                                reg1776 : forvar1774)) ?
                            ((reg1781 ?
                                reg1792 : reg1796) >>> $unsigned(reg1780)) : (&$signed((8'ha9))))));
  always
    @(posedge clk) begin
      reg1845 <= $unsigned(("paTQqZq" | $signed(reg1770[(4'h8):(1'h0)])));
      reg1846 <= $signed($unsigned({"eHR55", (^~forvar1814[(4'he):(4'hd)])}));
      reg1847 <= $unsigned($signed(($signed(reg1763) && $signed((8'h9c)))));
      for (forvar1848 = (1'h0); (forvar1848 < (2'h2)); forvar1848 = (forvar1848 + (1'h1)))
        begin
          reg1849 <= "f8htsiVM";
          reg1850 <= $signed($signed((reg1837[(5'h11):(4'he)] ?
              "aBFbZByYLHXpe" : $signed({reg1782, reg1779}))));
          for (forvar1851 = (1'h0); (forvar1851 < (1'h0)); forvar1851 = (forvar1851 + (1'h1)))
            begin
              reg1852 <= (reg1812[(3'h4):(1'h1)] ?
                  "b0Xst4H67" : {"BZXG8omBfZ8r",
                      {((+wire1797) ? (wire1844 ? (8'hbb) : reg1782) : reg1805),
                          reg1794}});
              reg1853 <= $unsigned(((!(reg1800[(2'h3):(1'h0)] ?
                  "aKOn3DPcCgf" : (reg1758 ? reg1852 : reg1758))) ~^ reg1841));
              reg1854 <= $signed($signed(reg1796[(1'h0):(1'h0)]));
              reg1855 <= {{reg1821}};
              reg1856 <= {(reg1760[(1'h1):(1'h0)] <<< $signed($unsigned(reg1817)))};
              reg1857 = ({"lJx9iL7wSAcVFiCu4Uqx", reg1839[(4'h9):(2'h2)]} ?
                  reg1798 : {{$unsigned(reg1762),
                          {(reg1769 ? reg1821 : forvar1807)}}});
            end
          reg1858 <= (reg1791 && $unsigned(("xKuIA7F6LL9" >> $signed((reg1798 | reg1796)))));
          reg1859 <= $unsigned($unsigned(($unsigned("zsG3") + reg1798[(4'he):(4'h9)])));
          for (forvar1860 = (1'h0); (forvar1860 < (1'h1)); forvar1860 = (forvar1860 + (1'h1)))
            begin
              reg1861 <= $signed($unsigned(reg1835[(3'h4):(2'h2)]));
              reg1862 = (~"ofPnLfDbaPO5");
              reg1863 <= "i";
              reg1864 <= $signed(({(8'hb7), $signed((reg1822 >= (8'ha2)))} ?
                  ((^~(~&forvar1814)) < ($signed(reg1792) ?
                      (reg1763 ?
                          reg1779 : forvar1765) : "vNqpV")) : ("NYfNXzUlPwkA2FDBw2" ?
                      reg1782 : "VBC")));
            end
        end
      reg1865 <= "9Ooq0pGffRaBAUaR81wRqd9";
    end
  always
    @(posedge clk) begin
      reg1866 <= reg1770[(4'h8):(3'h5)];
      reg1867 = reg1782;
      reg1868 <= {$unsigned(reg1817), {(&(+reg1819[(1'h0):(1'h0)]))}};
      reg1869 <= reg1780;
      for (forvar1870 = (1'h0); (forvar1870 < (2'h3)); forvar1870 = (forvar1870 + (1'h1)))
        begin
          for (forvar1871 = (1'h0); (forvar1871 < (2'h2)); forvar1871 = (forvar1871 + (1'h1)))
            begin
              reg1872 = $signed(reg1853[(5'h10):(4'hc)]);
              for (forvar1873 = (1'h0); (forvar1873 < (2'h3)); forvar1873 = (forvar1873 + (1'h1)))
                begin
                  reg1874 <= reg1800[(2'h3):(2'h2)];
                  reg1875 <= "Xzm9w2cn9";
                  reg1876 <= forvar1765;
                  reg1877 <= (reg1781[(5'h10):(4'ha)] ?
                      $signed(({{reg1770}, reg1847[(5'h10):(1'h1)]} ?
                          reg1810[(5'h17):(1'h1)] : $signed(reg1769))) : reg1853[(3'h6):(3'h4)]);
                end
            end
          for (forvar1878 = (1'h0); (forvar1878 < (3'h4)); forvar1878 = (forvar1878 + (1'h1)))
            begin
              for (forvar1879 = (1'h0); (forvar1879 < (1'h1)); forvar1879 = (forvar1879 + (1'h1)))
                begin
                  reg1880 <= "MhWS9TFVZUks6";
                  reg1881 <= $unsigned(reg1855[(3'h6):(2'h3)]);
                  reg1882 = $unsigned($unsigned((($signed(forvar1804) >>> (forvar1879 << reg1821)) >>> ("Wk61y3slgyJFQ2NEvUYn" ?
                      wire1844[(1'h1):(1'h1)] : {reg1794, reg1880}))));
                  reg1883 <= $signed(((~{forvar1815}) ?
                      {reg1852[(1'h1):(1'h1)]} : $signed($unsigned($signed(forvar1774)))));
                end
            end
          reg1884 <= (+(!forvar1871[(1'h1):(1'h0)]));
          reg1885 <= (~&(reg1834[(2'h3):(1'h0)] ?
              wire1756 : ($signed(reg1767[(4'h8):(4'h8)]) ?
                  reg1812 : (~(forvar1801 ? reg1810 : reg1872)))));
        end
      for (forvar1886 = (1'h0); (forvar1886 < (3'h5)); forvar1886 = (forvar1886 + (1'h1)))
        begin
          for (forvar1887 = (1'h0); (forvar1887 < (2'h2)); forvar1887 = (forvar1887 + (1'h1)))
            begin
              reg1888 <= (!"");
            end
          reg1889 <= ($signed({{reg1845[(3'h6):(2'h3)]}}) ?
              $unsigned(reg1872[(4'h9):(3'h4)]) : "dI7hHg");
          for (forvar1890 = (1'h0); (forvar1890 < (1'h1)); forvar1890 = (forvar1890 + (1'h1)))
            begin
              for (forvar1891 = (1'h0); (forvar1891 < (2'h2)); forvar1891 = (forvar1891 + (1'h1)))
                begin
                  reg1892 <= {forvar1807};
                  reg1893 <= forvar1890;
                  reg1894 = reg1841;
                  reg1895 <= reg1767[(3'h6):(3'h5)];
                end
              reg1896 <= (reg1824 ~^ (|(("b3hLrsyde6S1RPgn8zg" + "TxAKMM3Rkzx1XpL") == (reg1767 ?
                  "59fV1tMYmuzewxAbHNPai" : $signed(forvar1802)))));
              reg1897 <= $unsigned("XlhwczRY1WXN");
            end
          reg1898 <= $unsigned((reg1824 ?
              (reg1884[(3'h7):(3'h6)] ^ (reg1779[(1'h0):(1'h0)] ^~ "PWm3G")) : $unsigned($unsigned("aP8MckohesWWvcHJLuLK9"))));
          reg1899 <= (|$unsigned((|$signed({reg1829}))));
          for (forvar1900 = (1'h0); (forvar1900 < (1'h0)); forvar1900 = (forvar1900 + (1'h1)))
            begin
              reg1901 <= $signed((("I5ShadyS7r2oEaDGsOAo0hfN" - (8'ha2)) ?
                  ((!$signed((7'h40))) - (7'h43)) : $signed(((forvar1774 ?
                      reg1829 : reg1770) <= {reg1865}))));
              reg1902 <= $unsigned(reg1758);
              reg1903 <= reg1800[(2'h3):(2'h3)];
              reg1904 <= reg1777;
              reg1905 <= (+(|({(reg1827 != (7'h4d)),
                      "bqlae7nnz9ZXbwzRZyZc0Mc6"} ?
                  $signed((reg1828 || reg1764)) : (~&reg1813))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg1906 <= {"U"};
      reg1907 <= reg1874;
      reg1908 <= $signed(("qLrDYFHKgedz0mmMKot" ?
          $signed($unsigned(((8'hb0) && reg1781))) : forvar1804));
      for (forvar1909 = (1'h0); (forvar1909 < (1'h1)); forvar1909 = (forvar1909 + (1'h1)))
        begin
          reg1910 = "tIR0Gcrtf";
          reg1911 <= $signed((("GHoDxLREvzwERlLc" << reg1761) ?
              ($unsigned(reg1865[(5'h16):(2'h2)]) ?
                  (+$signed(reg1763)) : $signed((reg1828 ?
                      reg1853 : reg1872))) : "3"));
          reg1912 <= (^$signed(reg1880));
          if (($unsigned($signed(forvar1891[(3'h5):(1'h0)])) ?
              (reg1810[(4'hc):(3'h5)] ?
                  (^~{$signed(reg1859)}) : {"84sOzczzVqN"}) : (~$unsigned((reg1845 >= $unsigned(reg1877))))))
            begin
              reg1913 = $signed(reg1911[(3'h7):(3'h4)]);
              for (forvar1914 = (1'h0); (forvar1914 < (1'h0)); forvar1914 = (forvar1914 + (1'h1)))
                begin
                  reg1915 = $unsigned($signed(forvar1804[(4'h9):(3'h5)]));
                  reg1916 = (|reg1762);
                  reg1917 <= "8nIVpmwJpe2J4uE43tg";
                  reg1918 <= (^~(reg1868[(5'h16):(4'hc)] ^~ $unsigned(reg1770[(4'ha):(2'h3)])));
                  reg1919 = $signed({(+(~&(forvar1886 ? (8'ha8) : reg1837))),
                      ((-$signed((7'h43))) ~^ ($unsigned(reg1762) ^~ {(8'hbb),
                          reg1889}))});
                  reg1920 = forvar1870;
                end
              reg1921 <= $signed($unsigned($unsigned((~^$signed((8'ha7))))));
              for (forvar1922 = (1'h0); (forvar1922 < (2'h3)); forvar1922 = (forvar1922 + (1'h1)))
                begin
                  reg1923 = reg1884;
                end
              reg1924 <= reg1863[(1'h1):(1'h0)];
            end
          else
            begin
              reg1913 = $unsigned({$unsigned((!$signed(reg1766)))});
              reg1914 = (("x5slExVs" > (((forvar1860 ? reg1769 : reg1812) ?
                      $signed(reg1808) : (reg1896 || reg1782)) ?
                  $signed($signed(reg1829)) : ($signed((7'h47)) ?
                      {reg1917} : (reg1862 >> reg1772)))) == "3puumeBgCAlaK");
              for (forvar1915 = (1'h0); (forvar1915 < (3'h4)); forvar1915 = (forvar1915 + (1'h1)))
                begin
                  reg1916 <= ($signed(reg1817) != reg1812);
                  reg1917 <= $signed(reg1912);
                  reg1918 <= ((reg1867 >= $signed($unsigned($unsigned(reg1916)))) ?
                      reg1915 : reg1881[(2'h2):(2'h2)]);
                  reg1919 <= reg1903[(3'h5):(1'h0)];
                end
              for (forvar1920 = (1'h0); (forvar1920 < (3'h5)); forvar1920 = (forvar1920 + (1'h1)))
                begin
                  reg1921 <= (^(!reg1805[(4'h8):(3'h6)]));
                  reg1922 <= reg1798;
                end
              reg1923 <= $unsigned("OrM");
            end
        end
      reg1925 = reg1792;
      reg1926 <= (-$signed((~^reg1855[(5'h11):(3'h7)])));
    end
  assign wire1927 = ((reg1841 != forvar1801) < {forvar1765,
                        (-$unsigned((^~reg1766)))});
  assign wire1928 = "hI9BxDbIJdNeeA7";
  assign wire1929 = $unsigned(((("1LPG" - (wire1755 ? reg1914 : reg1859)) ?
                            ((reg1872 ? reg1921 : reg1858) ?
                                reg1867[(3'h4):(2'h3)] : $unsigned(reg1857)) : forvar1774[(4'h8):(3'h4)]) ?
                        (reg1771 & reg1831[(3'h6):(1'h1)]) : reg1846[(3'h7):(3'h5)]));
  always
    @(posedge clk) begin
      reg1930 = reg1913[(1'h0):(1'h0)];
    end
  assign wire1931 = (({($signed(reg1822) != wire1929)} >= reg1806[(3'h4):(1'h1)]) ?
                        {$signed(("A97z6HAaJAkglz43lds20RMm" * (reg1915 >> forvar1815))),
                            $signed((~|reg1913))} : reg1824);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1554
#( parameter param1662 = ({(~&(((8'hba) || (7'h45)) ? ((7'h49) << (7'h47)) : ((8'hb4) == (8'hb3)))), (({(8'h9e), (8'ha3)} || ((8'hbe) <= (7'h43))) & (7'h48))} != (({(&(8'ha8)), {(8'hba), (7'h4d)}} ? (((8'ha4) <= (8'hb8)) ? ((8'haa) ? (8'hac) : (8'hb3)) : (+(7'h45))) : ((&(8'hb5)) ? {(8'h9d)} : (^~(7'h49)))) && {{((7'h47) ? (8'hbc) : (8'ha7))}}))
, parameter param1663 = (~^param1662) )
(y, clk, wire1559, wire1558, wire1557, wire1556, wire1555);
  output wire [(32'h5a6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire1559;
  input wire signed [(3'h7):(1'h0)] wire1558;
  input wire [(4'ha):(1'h0)] wire1557;
  input wire [(4'he):(1'h0)] wire1556;
  input wire signed [(5'h15):(1'h0)] wire1555;
  reg [(5'h16):(1'h0)] reg1661 = (1'h0);
  reg [(4'h8):(1'h0)] reg1660 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1659 = (1'h0);
  reg [(4'he):(1'h0)] reg1658 = (1'h0);
  reg [(5'h17):(1'h0)] reg1657 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1656 = (1'h0);
  reg [(5'h17):(1'h0)] reg1655 = (1'h0);
  reg [(2'h3):(1'h0)] reg1654 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1653 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1652 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1651 = (1'h0);
  reg [(4'he):(1'h0)] reg1650 = (1'h0);
  reg [(5'h18):(1'h0)] reg1643 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1649 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1648 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1647 = (1'h0);
  reg [(5'h16):(1'h0)] reg1646 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1645 = (1'h0);
  reg [(3'h5):(1'h0)] reg1644 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1643 = (1'h0);
  reg [(4'h8):(1'h0)] reg1642 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1641 = (1'h0);
  reg [(2'h2):(1'h0)] reg1640 = (1'h0);
  reg [(4'hd):(1'h0)] reg1639 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1638 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1637 = (1'h0);
  reg [(4'hd):(1'h0)] reg1636 = (1'h0);
  reg [(4'hd):(1'h0)] reg1635 = (1'h0);
  reg [(3'h6):(1'h0)] reg1634 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1633 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1632 = (1'h0);
  reg [(5'h12):(1'h0)] reg1631 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1630 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire1629;
  reg [(3'h6):(1'h0)] reg1628 = (1'h0);
  reg [(5'h12):(1'h0)] reg1627 = (1'h0);
  wire signed [(4'he):(1'h0)] wire1626;
  reg signed [(5'h11):(1'h0)] reg1625 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1624 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1623 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1622 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1621 = (1'h0);
  reg [(2'h2):(1'h0)] reg1620 = (1'h0);
  reg [(4'he):(1'h0)] reg1619 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1618 = (1'h0);
  reg [(5'h12):(1'h0)] reg1617 = (1'h0);
  reg [(5'h11):(1'h0)] reg1616 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1615 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1614 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1613 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1612 = (1'h0);
  reg [(5'h10):(1'h0)] reg1611 = (1'h0);
  reg [(4'h8):(1'h0)] reg1610 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1609 = (1'h0);
  reg [(4'ha):(1'h0)] reg1608 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1607 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1606 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1605 = (1'h0);
  reg [(4'hb):(1'h0)] reg1604 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1603 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1602 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1601 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1600 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1599 = (1'h0);
  reg [(4'hf):(1'h0)] reg1598 = (1'h0);
  reg [(5'h16):(1'h0)] reg1597 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1596 = (1'h0);
  reg [(5'h19):(1'h0)] reg1595 = (1'h0);
  reg [(5'h13):(1'h0)] reg1594 = (1'h0);
  reg [(5'h19):(1'h0)] reg1593 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1592 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1591 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1590 = (1'h0);
  reg [(3'h5):(1'h0)] reg1589 = (1'h0);
  reg [(4'hc):(1'h0)] reg1588 = (1'h0);
  reg [(5'h12):(1'h0)] reg1587 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1586 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1585 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1584 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1583 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1582 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1581 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1580 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1579 = (1'h0);
  reg [(2'h3):(1'h0)] reg1578 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1577 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1576 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1575 = (1'h0);
  reg [(5'h14):(1'h0)] reg1574 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1573 = (1'h0);
  reg [(5'h18):(1'h0)] reg1572 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1571 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1570 = (1'h0);
  reg [(4'hf):(1'h0)] reg1569 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1568 = (1'h0);
  reg [(4'hf):(1'h0)] reg1567 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1566 = (1'h0);
  reg [(3'h4):(1'h0)] reg1565 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1564 = (1'h0);
  wire [(5'h12):(1'h0)] wire1563;
  wire [(3'h7):(1'h0)] wire1562;
  wire signed [(5'h17):(1'h0)] wire1561;
  reg signed [(5'h16):(1'h0)] reg1560 = (1'h0);
  assign y = {reg1661,
                 reg1660,
                 reg1659,
                 reg1658,
                 reg1657,
                 reg1656,
                 reg1655,
                 reg1654,
                 forvar1653,
                 forvar1652,
                 reg1651,
                 reg1650,
                 reg1643,
                 reg1649,
                 reg1648,
                 reg1647,
                 reg1646,
                 reg1645,
                 reg1644,
                 forvar1643,
                 reg1642,
                 reg1641,
                 reg1640,
                 reg1639,
                 reg1638,
                 reg1637,
                 reg1636,
                 reg1635,
                 reg1634,
                 forvar1633,
                 reg1632,
                 reg1631,
                 forvar1630,
                 wire1629,
                 reg1628,
                 reg1627,
                 wire1626,
                 reg1625,
                 reg1624,
                 reg1623,
                 reg1622,
                 reg1621,
                 reg1620,
                 reg1619,
                 reg1618,
                 reg1617,
                 reg1616,
                 forvar1615,
                 reg1614,
                 reg1613,
                 reg1612,
                 reg1611,
                 reg1610,
                 reg1609,
                 reg1608,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1604,
                 reg1603,
                 reg1602,
                 forvar1601,
                 reg1600,
                 reg1599,
                 reg1598,
                 reg1597,
                 forvar1596,
                 reg1595,
                 reg1594,
                 reg1593,
                 reg1592,
                 forvar1591,
                 reg1590,
                 reg1589,
                 reg1588,
                 reg1587,
                 reg1586,
                 forvar1585,
                 forvar1584,
                 reg1583,
                 reg1582,
                 reg1581,
                 reg1580,
                 reg1579,
                 reg1578,
                 forvar1577,
                 forvar1576,
                 reg1575,
                 reg1574,
                 reg1573,
                 reg1572,
                 forvar1571,
                 reg1570,
                 reg1569,
                 reg1568,
                 reg1567,
                 reg1566,
                 reg1565,
                 reg1564,
                 wire1563,
                 wire1562,
                 wire1561,
                 reg1560,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1560 <= wire1558[(3'h4):(1'h0)];
    end
  assign wire1561 = $signed(wire1559[(3'h7):(3'h6)]);
  assign wire1562 = ("7uS1gaAc6q9TrMO4lG54fvI" ?
                        ($unsigned(wire1555[(5'h14):(4'h9)]) ~^ "5") : (reg1560[(4'h8):(4'h8)] ?
                            (!wire1556) : ($signed(wire1557[(4'h9):(4'h9)]) ?
                                $unsigned((+reg1560)) : "vd4anQ0g")));
  assign wire1563 = $unsigned($signed(wire1557[(2'h3):(2'h2)]));
  always
    @(posedge clk) begin
      reg1564 <= wire1558;
      reg1565 <= $signed(($unsigned("NNCnmqb3Om") ?
          wire1555 : $signed((wire1558[(3'h4):(3'h4)] == (wire1558 ?
              reg1560 : wire1561)))));
      reg1566 <= wire1557;
    end
  always
    @(posedge clk) begin
      reg1567 <= reg1564;
      reg1568 <= reg1565[(2'h2):(2'h2)];
      reg1569 <= wire1558[(2'h3):(1'h0)];
      reg1570 = wire1557[(3'h5):(2'h3)];
    end
  always
    @(posedge clk) begin
      for (forvar1571 = (1'h0); (forvar1571 < (3'h4)); forvar1571 = (forvar1571 + (1'h1)))
        begin
          reg1572 <= (8'ha6);
          reg1573 <= {($unsigned($unsigned({wire1555,
                  (8'h9c)})) >= (!(-"SdPdxR"))),
              $unsigned(reg1566)};
          reg1574 <= (!$signed($unsigned(({wire1561} <<< wire1557))));
          reg1575 <= reg1572;
        end
      for (forvar1576 = (1'h0); (forvar1576 < (3'h4)); forvar1576 = (forvar1576 + (1'h1)))
        begin
          for (forvar1577 = (1'h0); (forvar1577 < (2'h3)); forvar1577 = (forvar1577 + (1'h1)))
            begin
              reg1578 <= ($unsigned(reg1565) >> (~$signed($signed(wire1562[(2'h3):(1'h1)]))));
              reg1579 <= reg1564[(4'h8):(2'h2)];
              reg1580 <= wire1563[(4'hc):(4'h8)];
              reg1581 <= reg1567[(4'h9):(3'h4)];
            end
          reg1582 = $unsigned({($signed({forvar1571}) ?
                  wire1557[(4'ha):(2'h3)] : {reg1569, $signed(wire1561)}),
              (&"0qikC4")});
          reg1583 = wire1555[(3'h7):(1'h1)];
          for (forvar1584 = (1'h0); (forvar1584 < (2'h3)); forvar1584 = (forvar1584 + (1'h1)))
            begin
              for (forvar1585 = (1'h0); (forvar1585 < (1'h1)); forvar1585 = (forvar1585 + (1'h1)))
                begin
                  reg1586 = ({"6h8ZzDLLoVz", reg1574[(1'h1):(1'h1)]} ?
                      $signed(($signed({reg1582}) <= ($unsigned(forvar1571) ?
                          reg1570 : reg1569[(4'ha):(2'h3)]))) : forvar1584);
                  reg1587 <= reg1566;
                  reg1588 <= reg1586[(3'h5):(1'h0)];
                end
              reg1589 <= {({((wire1562 ?
                              wire1556 : (8'h9c)) + $unsigned((8'hb1))),
                          $signed({reg1564})} ?
                      (8'hb5) : (8'ha9)),
                  reg1568[(1'h1):(1'h0)]};
              reg1590 = $signed($signed($signed("ND")));
              for (forvar1591 = (1'h0); (forvar1591 < (1'h1)); forvar1591 = (forvar1591 + (1'h1)))
                begin
                  reg1592 <= "mxA";
                end
            end
          reg1593 <= $signed("AcVf02gwVJP");
          reg1594 <= $unsigned(forvar1571);
        end
      reg1595 <= $signed(((reg1583[(3'h5):(3'h5)] ?
          {$signed(wire1561)} : (!wire1557[(3'h6):(3'h4)])) - (~^$signed({(8'h9f)}))));
      for (forvar1596 = (1'h0); (forvar1596 < (2'h2)); forvar1596 = (forvar1596 + (1'h1)))
        begin
          reg1597 <= $signed("WWeC8Wsb3W6");
          reg1598 <= ($signed((!(8'hb1))) ^ "niUlfftRIpFRwWqWAbBltVXa");
          reg1599 <= $unsigned("bX8bmZ4");
          reg1600 <= (8'ha8);
        end
    end
  always
    @(posedge clk) begin
      for (forvar1601 = (1'h0); (forvar1601 < (1'h0)); forvar1601 = (forvar1601 + (1'h1)))
        begin
          reg1602 <= ($unsigned(("MxQUnhsqRv" >> (-(wire1561 ?
                  wire1555 : (8'had))))) ?
              $unsigned({forvar1576[(1'h0):(1'h0)]}) : reg1594[(4'ha):(2'h2)]);
          reg1603 <= {reg1600[(4'hb):(2'h2)],
              $unsigned(($signed({(8'ha0), reg1586}) ?
                  (8'ha3) : $signed(reg1589)))};
          reg1604 <= reg1564[(2'h3):(2'h2)];
          reg1605 = "";
          reg1606 <= (~^("bHZgNDgypBJD5Eu" == $signed($unsigned((8'hbc)))));
          reg1607 = ((8'hbd) ?
              (((~&(reg1595 ? reg1600 : forvar1601)) ?
                  (8'ha4) : {"LfM0cVJbi7k"}) << $unsigned((!$unsigned(reg1582)))) : "UdA2f2qiCmILKkThPRah0R1EZ");
        end
      reg1608 <= "fiswqH9uqCxMeDtkzkx";
      reg1609 = (|"lIzqMIx3T07BIu");
      reg1610 <= reg1574;
    end
  always
    @(posedge clk) begin
      reg1611 <= ("ZsCIlhEi1B9" << reg1595[(1'h0):(1'h0)]);
      reg1612 = reg1599;
      reg1613 <= ($signed((reg1583 ^~ $signed((reg1606 ?
              forvar1576 : (8'ha0))))) ?
          reg1609[(4'ha):(3'h4)] : (8'hb0));
      reg1614 <= "h1BrFKaH2z1YsvIg";
      for (forvar1615 = (1'h0); (forvar1615 < (2'h2)); forvar1615 = (forvar1615 + (1'h1)))
        begin
          reg1616 <= reg1589[(3'h4):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      reg1617 <= (reg1588[(4'h8):(3'h7)] ?
          $signed(($signed("f3NcB1DtQZ53V95") ?
              reg1578[(2'h3):(2'h2)] : $signed({reg1581}))) : (^~(8'hb7)));
    end
  always
    @(posedge clk) begin
      reg1618 <= $signed((((|(reg1592 * (8'ha2))) ?
              ($signed(reg1594) ?
                  (reg1603 ? (8'ha0) : reg1573) : (&forvar1577)) : reg1612) ?
          (reg1578 ? reg1580 : reg1603[(4'hc):(3'h5)]) : ($signed({reg1575}) ?
              reg1592 : reg1566)));
      reg1619 <= {forvar1591};
      reg1620 <= (-(8'hb5));
      reg1621 <= (~|{(reg1589 ?
              (~{wire1559, (8'hbc)}) : $unsigned($unsigned(forvar1577)))});
    end
  always
    @(posedge clk) begin
      reg1622 <= (wire1558[(3'h6):(3'h4)] - (~|(reg1567[(4'he):(4'ha)] << {(wire1557 ^ reg1574)})));
      reg1623 <= "Va";
      reg1624 <= (+($unsigned(("hQWu7R01sgE" + "6PYAvOaWK1mzbyMbE")) ?
          reg1560 : {wire1559}));
      reg1625 <= (-(forvar1577[(1'h0):(1'h0)] || reg1608));
    end
  assign wire1626 = (~&(&reg1619[(4'h8):(1'h1)]));
  always
    @(posedge clk) begin
      reg1627 <= {($unsigned(($signed(reg1580) >= reg1608)) << $signed((reg1599 - (reg1593 ?
              forvar1615 : reg1624)))),
          $signed(($unsigned((reg1568 ? reg1604 : reg1572)) * ((forvar1576 ?
              (7'h42) : reg1579) ^~ (forvar1577 ? reg1614 : wire1555))))};
      reg1628 <= reg1578[(2'h3):(2'h3)];
    end
  assign wire1629 = (-$signed(("Dh5hCtdQbP" >> $unsigned(reg1628[(2'h2):(1'h1)]))));
  always
    @(posedge clk) begin
      for (forvar1630 = (1'h0); (forvar1630 < (2'h2)); forvar1630 = (forvar1630 + (1'h1)))
        begin
          reg1631 = reg1606;
        end
      reg1632 <= $signed((~^(^~$signed($signed(reg1606)))));
      for (forvar1633 = (1'h0); (forvar1633 < (3'h5)); forvar1633 = (forvar1633 + (1'h1)))
        begin
          reg1634 <= reg1606[(4'h8):(1'h0)];
          reg1635 <= (&(("yrrbzo7EwRmBgEGCm" >= "6kwgw5") ?
              (-(forvar1615[(5'h10):(4'hf)] ?
                  (forvar1630 && reg1627) : "l9ltrUVz")) : ($unsigned(forvar1633) ?
                  reg1597[(5'h12):(5'h10)] : "")));
          reg1636 <= $signed(reg1564);
          reg1637 <= $unsigned((~|reg1610));
          reg1638 <= (reg1624 * $signed({reg1632[(4'hf):(4'hb)]}));
          if (($unsigned((&wire1626)) ?
              (~&$unsigned({$signed(reg1617),
                  $unsigned((7'h41))})) : (reg1568 || ($unsigned(reg1567) ~^ $unsigned((8'hb5))))))
            begin
              reg1639 <= "vDshSa4EYWQ";
              reg1640 <= (reg1589[(3'h5):(3'h4)] ^ (~^(~(~|$signed(reg1589)))));
              reg1641 <= $unsigned(reg1594);
              reg1642 <= reg1578;
              for (forvar1643 = (1'h0); (forvar1643 < (3'h4)); forvar1643 = (forvar1643 + (1'h1)))
                begin
                  reg1644 = (((~("tsWtJ" * forvar1585)) ?
                      (((forvar1596 - reg1617) + forvar1643) ?
                          (^~(wire1629 ?
                              (8'hbc) : reg1607)) : $unsigned((reg1611 * reg1631))) : "WgEnZrQ3xe8hd1KVvwSqS0wu3") == (reg1640[(2'h2):(1'h0)] ?
                      {$signed($signed((8'h9d)))} : $unsigned(($unsigned(reg1569) ?
                          {reg1565, reg1583} : (reg1593 ?
                              reg1610 : reg1565)))));
                  reg1645 <= (^~"Cc0R0KSMh");
                  reg1646 <= $unsigned(({reg1588[(4'h8):(3'h4)]} <= (reg1638 <= ((reg1623 ?
                      forvar1576 : reg1631) <= (wire1558 ?
                      reg1565 : reg1638)))));
                  reg1647 <= (~$unsigned((wire1558 ?
                      $unsigned((~|reg1619)) : (|reg1639))));
                  reg1648 <= wire1555;
                end
              reg1649 <= reg1600[(4'he):(4'ha)];
            end
          else
            begin
              reg1639 <= wire1629[(4'ha):(2'h2)];
              reg1640 <= $unsigned($unsigned((~^$signed(reg1564[(3'h7):(3'h5)]))));
              reg1641 <= $unsigned("HtQqOUfMsUW3md9o1XE1mhUp5");
              reg1642 <= ({reg1574, {{"a1"}}} ? forvar1585 : (~"X2iKkdGCE"));
              reg1643 <= reg1578;
            end
        end
      reg1650 <= ("6i" ?
          "kFQODhtUUH9p" : {(~({wire1555, (8'hae)} ?
                  reg1611 : reg1647[(4'h9):(4'h9)]))});
    end
  always
    @(posedge clk) begin
      reg1651 <= $unsigned(reg1560);
    end
  always
    @(posedge clk) begin
      for (forvar1652 = (1'h0); (forvar1652 < (2'h2)); forvar1652 = (forvar1652 + (1'h1)))
        begin
          for (forvar1653 = (1'h0); (forvar1653 < (1'h1)); forvar1653 = (forvar1653 + (1'h1)))
            begin
              reg1654 <= reg1570;
              reg1655 <= forvar1596[(4'hf):(3'h6)];
              reg1656 <= (8'ha4);
              reg1657 = {reg1603,
                  $unsigned($signed(((wire1563 >> reg1651) * $signed((7'h48)))))};
            end
          reg1658 <= "Ss74sEoGFrEwIlng0rWcogQ";
        end
      reg1659 <= (+(^("JKx2nykwaQ8EJEVT46qeob" ?
          (~|reg1649[(4'h8):(3'h5)]) : ((~forvar1576) ?
              $signed(reg1640) : reg1654))));
      reg1660 <= (!"a1h");
      reg1661 <= $unsigned("zDNPxcAV6X7");
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1446
#( parameter param1548 = (+(^(({(8'ha5), (8'ha4)} ? ((8'h9f) + (8'ha9)) : ((8'ha7) * (8'ha9))) ? {{(8'ha4)}} : ({(8'hb0)} + ((8'hba) ^ (8'h9c))))))
, parameter param1549 = {param1548} )
(y, clk, wire1450, wire1449, wire1448, wire1447);
  output wire [(32'h58a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire1450;
  input wire [(5'h13):(1'h0)] wire1449;
  input wire signed [(5'h1a):(1'h0)] wire1448;
  input wire [(5'h15):(1'h0)] wire1447;
  reg signed [(5'h14):(1'h0)] reg1547 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1546 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1545 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1544 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1543 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire1542;
  wire signed [(4'h8):(1'h0)] wire1541;
  reg signed [(4'hc):(1'h0)] reg1540 = (1'h0);
  reg [(4'ha):(1'h0)] reg1539 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1538 = (1'h0);
  reg [(5'h15):(1'h0)] reg1537 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1536 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1535 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1531 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1532 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1530 = (1'h0);
  reg [(4'hd):(1'h0)] reg1534 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1533 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1532 = (1'h0);
  reg [(5'h11):(1'h0)] reg1531 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1530 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1529 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1528 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1527 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1526 = (1'h0);
  reg [(5'h17):(1'h0)] reg1525 = (1'h0);
  reg [(2'h2):(1'h0)] reg1524 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1523 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1522 = (1'h0);
  reg [(5'h13):(1'h0)] reg1521 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1520 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1519 = (1'h0);
  reg [(3'h7):(1'h0)] reg1518 = (1'h0);
  reg [(5'h12):(1'h0)] reg1517 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1516 = (1'h0);
  reg [(2'h3):(1'h0)] reg1515 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1514 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1513 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1512 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1511 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1510 = (1'h0);
  reg [(5'h18):(1'h0)] reg1509 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1508 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1507 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1506 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1505 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire1504;
  wire signed [(4'he):(1'h0)] wire1503;
  reg signed [(4'he):(1'h0)] reg1502 = (1'h0);
  reg [(5'h14):(1'h0)] reg1501 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1500 = (1'h0);
  reg [(4'he):(1'h0)] reg1499 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1498 = (1'h0);
  reg [(5'h12):(1'h0)] reg1497 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1496 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1495 = (1'h0);
  reg [(3'h4):(1'h0)] reg1494 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1493 = (1'h0);
  reg [(3'h7):(1'h0)] reg1492 = (1'h0);
  reg [(3'h4):(1'h0)] reg1491 = (1'h0);
  reg [(5'h17):(1'h0)] reg1490 = (1'h0);
  reg [(4'hd):(1'h0)] reg1489 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1488 = (1'h0);
  wire [(4'ha):(1'h0)] wire1487;
  reg signed [(3'h6):(1'h0)] reg1486 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1485 = (1'h0);
  reg [(4'he):(1'h0)] reg1484 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1483 = (1'h0);
  reg [(4'h8):(1'h0)] reg1482 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1481 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1480 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1479 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1478 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1477 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1476 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1475 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1474 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1473 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1472 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1471 = (1'h0);
  reg [(4'hd):(1'h0)] reg1470 = (1'h0);
  reg [(5'h16):(1'h0)] reg1469 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1468 = (1'h0);
  reg [(3'h4):(1'h0)] reg1467 = (1'h0);
  reg [(5'h16):(1'h0)] reg1466 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1465 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1464 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire1463;
  wire signed [(2'h2):(1'h0)] wire1462;
  reg signed [(5'h10):(1'h0)] reg1461 = (1'h0);
  reg [(4'hb):(1'h0)] reg1460 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire1459;
  reg [(4'hf):(1'h0)] reg1458 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1457 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1456 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1455 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1454 = (1'h0);
  reg [(4'he):(1'h0)] reg1453 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1452 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1451 = (1'h0);
  assign y = {reg1547,
                 reg1546,
                 reg1545,
                 reg1544,
                 reg1543,
                 wire1542,
                 wire1541,
                 reg1540,
                 reg1539,
                 reg1538,
                 reg1537,
                 reg1536,
                 forvar1535,
                 forvar1531,
                 reg1532,
                 reg1530,
                 reg1534,
                 reg1533,
                 forvar1532,
                 reg1531,
                 forvar1530,
                 reg1529,
                 reg1528,
                 reg1527,
                 forvar1526,
                 reg1525,
                 reg1524,
                 reg1523,
                 reg1522,
                 reg1521,
                 reg1520,
                 reg1519,
                 reg1518,
                 reg1517,
                 reg1516,
                 reg1515,
                 forvar1514,
                 reg1513,
                 reg1512,
                 reg1511,
                 reg1510,
                 reg1509,
                 forvar1508,
                 reg1507,
                 reg1506,
                 forvar1505,
                 wire1504,
                 wire1503,
                 reg1502,
                 reg1501,
                 reg1500,
                 reg1499,
                 forvar1498,
                 reg1497,
                 reg1496,
                 reg1495,
                 reg1494,
                 forvar1493,
                 reg1492,
                 reg1491,
                 reg1490,
                 reg1489,
                 forvar1488,
                 wire1487,
                 reg1486,
                 reg1485,
                 reg1484,
                 reg1483,
                 reg1482,
                 reg1481,
                 reg1480,
                 reg1479,
                 reg1478,
                 reg1477,
                 reg1476,
                 reg1475,
                 reg1474,
                 reg1473,
                 reg1472,
                 forvar1471,
                 reg1470,
                 reg1469,
                 reg1468,
                 reg1467,
                 reg1466,
                 reg1465,
                 forvar1464,
                 wire1463,
                 wire1462,
                 reg1461,
                 reg1460,
                 wire1459,
                 reg1458,
                 forvar1457,
                 reg1456,
                 reg1455,
                 reg1454,
                 reg1453,
                 reg1452,
                 reg1451,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1451 <= wire1449[(3'h5):(3'h4)];
      reg1452 = ("0dgJEiRSVvLcTySq0GfcGW6KG" >>> ($signed((((8'ha8) >> wire1450) ?
              reg1451[(2'h3):(2'h3)] : $signed((8'ha7)))) ?
          $signed(reg1451) : (8'hac)));
      reg1453 <= $signed((wire1449[(5'h12):(1'h0)] ?
          ("FatG1uRzZ9eCIEBUq0ly67" || ((+(8'hb9)) && {reg1452,
              wire1447})) : (~^reg1451[(2'h3):(1'h0)])));
      reg1454 <= (($unsigned("z") < $signed($signed($unsigned(wire1447)))) ?
          (wire1450[(1'h0):(1'h0)] | "Vmea4wUXVds5JnoeprTBB") : "AnhGxcotY");
      reg1455 <= wire1447;
      reg1456 <= reg1453[(2'h3):(2'h3)];
    end
  always
    @(posedge clk) begin
      for (forvar1457 = (1'h0); (forvar1457 < (3'h5)); forvar1457 = (forvar1457 + (1'h1)))
        begin
          reg1458 <= reg1455;
        end
    end
  assign wire1459 = ((+(reg1454[(4'hc):(4'h8)] ?
                            (reg1455 | (reg1452 ^ reg1453)) : ((wire1449 > reg1458) ?
                                reg1455[(3'h4):(1'h1)] : (wire1449 <<< wire1450)))) ?
                        ($unsigned(wire1449[(4'h8):(3'h7)]) < wire1447) : (($unsigned($signed(reg1456)) ?
                            reg1454[(1'h0):(1'h0)] : (reg1451 ?
                                reg1451[(4'h9):(2'h3)] : (wire1450 << wire1447))) ^ $unsigned(reg1455)));
  always
    @(posedge clk) begin
      reg1460 <= $unsigned("1Koy56mirZ5v1QbIGYYk0v");
      reg1461 = {$unsigned((-wire1447))};
    end
  assign wire1462 = ({("m0hp1nix" ?
                            $unsigned((forvar1457 >= reg1461)) : (~reg1458))} < wire1459[(1'h0):(1'h0)]);
  assign wire1463 = reg1452;
  always
    @(posedge clk) begin
      for (forvar1464 = (1'h0); (forvar1464 < (1'h0)); forvar1464 = (forvar1464 + (1'h1)))
        begin
          reg1465 <= (~^$signed(reg1451[(3'h5):(3'h5)]));
          reg1466 <= (reg1455 ?
              reg1454 : ((-(((8'hb7) | wire1459) >> ((8'hb9) | (7'h42)))) ?
                  reg1452 : $unsigned("AAZTr4")));
          reg1467 <= (&reg1456[(1'h1):(1'h1)]);
          reg1468 <= (-(~|$unsigned(("LHoHr9" << (wire1449 != wire1463)))));
          reg1469 = reg1454;
          reg1470 <= ({reg1453} | $unsigned((^~$unsigned((reg1469 == (8'hab))))));
        end
      for (forvar1471 = (1'h0); (forvar1471 < (1'h0)); forvar1471 = (forvar1471 + (1'h1)))
        begin
          reg1472 <= {($unsigned(wire1462) > (~^reg1455[(2'h2):(1'h1)])),
              (|(((reg1469 | reg1467) <<< $signed(wire1463)) != {$signed(wire1463)}))};
        end
      reg1473 = reg1465[(3'h5):(1'h1)];
      reg1474 <= ("G7kZ0FlaMrf" * reg1453[(3'h6):(3'h4)]);
      reg1475 <= {wire1448};
    end
  always
    @(posedge clk) begin
      reg1476 <= ({(8'ha9)} ?
          (reg1474[(1'h0):(1'h0)] ~^ ("dADQW3PzIXWBDL3O9lYWZa" - wire1462)) : forvar1457);
      reg1477 = "LEHu8ff";
      reg1478 <= $unsigned(reg1466);
      reg1479 <= $unsigned($signed(wire1462));
    end
  always
    @(posedge clk) begin
      reg1480 <= (~|wire1459);
      reg1481 = ($unsigned((((reg1456 << wire1459) ?
              $signed(reg1469) : $unsigned((7'h4d))) != $unsigned((~&forvar1464)))) ?
          reg1461 : "cSdsdTAx");
    end
  always
    @(posedge clk) begin
      reg1482 <= {$unsigned((reg1476[(3'h4):(1'h0)] + $unsigned((+wire1449))))};
      reg1483 <= ("MIgUaLFxf" >> ({{(forvar1457 * reg1451),
              $unsigned(reg1451)}} << (((reg1458 * reg1482) <= reg1481[(3'h5):(1'h1)]) ^~ (&$unsigned(reg1454)))));
      reg1484 <= (~^wire1462);
      reg1485 = (&(wire1463[(4'h8):(3'h7)] ~^ reg1481));
      reg1486 <= (|{reg1483[(2'h3):(1'h1)],
          ($signed(wire1449[(5'h13):(3'h6)]) ~^ (reg1477 ?
              reg1460 : ((8'hb2) ? reg1451 : reg1461)))});
    end
  assign wire1487 = $unsigned((!wire1449));
  always
    @(posedge clk) begin
      for (forvar1488 = (1'h0); (forvar1488 < (1'h0)); forvar1488 = (forvar1488 + (1'h1)))
        begin
          reg1489 = (+$signed((~^$signed((+reg1482)))));
          reg1490 = $signed($unsigned($signed($unsigned(reg1478))));
          reg1491 = (wire1487[(3'h5):(3'h4)] ?
              $signed((!forvar1471[(1'h1):(1'h1)])) : (+("lu5OFHFisfICWw0" && $signed("emS60Xhe"))));
          reg1492 = $signed($signed(({reg1472[(3'h6):(1'h1)]} + ($signed(reg1482) != (reg1479 | reg1454)))));
          for (forvar1493 = (1'h0); (forvar1493 < (1'h0)); forvar1493 = (forvar1493 + (1'h1)))
            begin
              reg1494 = $unsigned($signed((8'haf)));
              reg1495 <= $signed(reg1476[(1'h0):(1'h0)]);
            end
          reg1496 <= "6";
        end
      reg1497 <= $unsigned(((^wire1487) ~^ $unsigned("KOUM5V7rgbMaffi")));
      for (forvar1498 = (1'h0); (forvar1498 < (1'h0)); forvar1498 = (forvar1498 + (1'h1)))
        begin
          reg1499 <= "VbUk";
          reg1500 = forvar1457[(2'h2):(1'h0)];
          reg1501 = reg1477[(3'h5):(1'h1)];
          reg1502 <= "ibXIS0hy";
        end
    end
  assign wire1503 = reg1458;
  assign wire1504 = "t7MPGQhZ2Nbo5";
  always
    @(posedge clk) begin
      for (forvar1505 = (1'h0); (forvar1505 < (2'h3)); forvar1505 = (forvar1505 + (1'h1)))
        begin
          reg1506 <= "tSv6Y4JGQRhQQ";
          reg1507 <= (+(wire1462 * $signed(reg1467[(1'h1):(1'h0)])));
          for (forvar1508 = (1'h0); (forvar1508 < (1'h1)); forvar1508 = (forvar1508 + (1'h1)))
            begin
              reg1509 <= (8'h9e);
              reg1510 <= reg1455;
            end
          reg1511 <= "uf";
        end
      reg1512 <= ((~&("CJtM48Yvi" ?
          (((8'hab) ? reg1458 : wire1448) ?
              (8'hbd) : $signed(reg1474)) : "mcu4ncW4nWLAB")) >>> $unsigned(("4dU2ufPYAogf" ?
          $unsigned("HYMrmoXc0rYQXz") : reg1470[(2'h2):(1'h0)])));
      reg1513 <= (&$unsigned($signed($signed((wire1462 != reg1512)))));
      for (forvar1514 = (1'h0); (forvar1514 < (1'h1)); forvar1514 = (forvar1514 + (1'h1)))
        begin
          reg1515 <= reg1480;
          reg1516 <= reg1506[(3'h6):(2'h3)];
          reg1517 <= $unsigned(reg1490[(4'ha):(4'h9)]);
        end
    end
  always
    @(posedge clk) begin
      reg1518 = (^"8WmcV");
      reg1519 <= reg1495[(3'h4):(2'h3)];
      if ($unsigned(reg1483))
        begin
          reg1520 <= "K";
          reg1521 = ((~&("A69oprHb9tizFUxn90P61P" ?
              ($unsigned((7'h4e)) ?
                  $unsigned((7'h43)) : {forvar1493,
                      reg1456}) : $unsigned($signed(reg1502)))) ^ (8'hb4));
          reg1522 = (reg1480 >>> ((^~(^$signed(wire1504))) == reg1452[(4'he):(4'he)]));
          reg1523 = (8'ha5);
          reg1524 <= (8'hb1);
        end
      else
        begin
          reg1520 = (8'hb8);
          reg1521 <= reg1452;
        end
      reg1525 <= ((&(8'hbf)) & reg1500);
    end
  always
    @(posedge clk) begin
      for (forvar1526 = (1'h0); (forvar1526 < (1'h0)); forvar1526 = (forvar1526 + (1'h1)))
        begin
          reg1527 <= (~$signed("5hTNH"));
          reg1528 <= reg1472;
        end
      if (("qQIT4YXu0bYZntx4iZtLUNce" ?
          $signed({$unsigned((!reg1520))}) : wire1447))
        begin
          reg1529 <= $unsigned(reg1470[(4'hb):(1'h1)]);
          for (forvar1530 = (1'h0); (forvar1530 < (2'h2)); forvar1530 = (forvar1530 + (1'h1)))
            begin
              reg1531 <= reg1456[(3'h4):(2'h2)];
              for (forvar1532 = (1'h0); (forvar1532 < (3'h5)); forvar1532 = (forvar1532 + (1'h1)))
                begin
                  reg1533 = "PaTiBRXqry4doywcE";
                end
            end
          reg1534 = reg1454;
        end
      else
        begin
          reg1529 <= ((((^~reg1460[(4'ha):(1'h0)]) ? "Nk" : (^(!reg1482))) ?
                  $signed({$signed(reg1520),
                      $signed(reg1524)}) : ($unsigned({wire1503}) ~^ (((8'ha0) ?
                          reg1474 : reg1451) ?
                      (~^wire1503) : (reg1515 ? (8'ha4) : reg1522)))) ?
              "AMG" : "M");
          reg1530 <= ({"Osldqt00hqwRNW15a2B0zf"} ?
              reg1494[(2'h2):(1'h0)] : $unsigned(reg1534));
          if ($signed($unsigned(($unsigned((&reg1520)) * $signed((!reg1481))))))
            begin
              reg1531 <= (|"Qtus5");
              reg1532 = "UEL";
              reg1533 <= (^~("hhEEPKF" ?
                  $unsigned(($unsigned(forvar1514) ?
                      reg1472 : {reg1494})) : reg1525[(3'h4):(3'h4)]));
            end
          else
            begin
              for (forvar1531 = (1'h0); (forvar1531 < (3'h4)); forvar1531 = (forvar1531 + (1'h1)))
                begin
                  reg1532 <= (|reg1511[(3'h4):(1'h0)]);
                end
              reg1533 <= reg1525[(5'h13):(4'hf)];
              reg1534 <= (((((reg1476 || reg1473) >>> wire1450[(3'h4):(1'h1)]) ?
                  "h6SYPFAhNmyf" : (forvar1464 ~^ (7'h4b))) * $signed("70MhpOm")) != ((~|($unsigned(reg1484) ?
                      ((7'h4b) != reg1452) : $signed(reg1502))) ?
                  reg1510 : (^((reg1484 != forvar1532) ?
                      $unsigned(reg1482) : "95any9"))));
              for (forvar1535 = (1'h0); (forvar1535 < (3'h5)); forvar1535 = (forvar1535 + (1'h1)))
                begin
                  reg1536 = $signed((~&$signed(reg1490[(5'h17):(4'hf)])));
                end
            end
          reg1537 = $signed("XwJBSrOlzen");
          reg1538 <= ($signed(reg1491[(3'h4):(1'h1)]) ^~ ((((reg1486 ?
              (8'hb9) : reg1461) ^~ (-reg1482)) == $unsigned(reg1472[(3'h7):(2'h2)])) | reg1515));
        end
      reg1539 <= $unsigned(((($unsigned(reg1453) >>> $signed((8'h9f))) && "cbDkmPnOQlirC3") ^ "9"));
      reg1540 <= ((~^"6pNZO7ehRPqehldV2GzeBRK") & (+$signed("N5YDR2au3AXUoLZ2n")));
    end
  assign wire1541 = $unsigned("HSQHe58E5KfHYTdbIaqMbiBI");
  assign wire1542 = $signed("NPrbQo8yQPHZS");
  always
    @(posedge clk) begin
      reg1543 <= $unsigned($unsigned(reg1477[(4'h8):(2'h3)]));
      reg1544 <= "JuTLoV";
      reg1545 <= $unsigned(reg1486[(3'h5):(2'h3)]);
      reg1546 = "LPAqahrKqxiXFi4JZbt4IY";
      reg1547 <= "uNi5pCt2pkXH5aSB";
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1383
#( parameter param1441 = {(~(({(7'h41), (8'hb9)} ? ((7'h41) ? (7'h4d) : (8'hab)) : {(7'h41), (8'h9c)}) & ((~&(8'ha6)) ? ((8'hb7) >>> (7'h4d)) : (~&(8'ha5)))))}
, parameter param1442 = (~|(~|param1441)) )
(y, clk, wire1387, wire1386, wire1385, wire1384);
  output wire [(32'h23f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire1387;
  input wire [(4'ha):(1'h0)] wire1386;
  input wire signed [(5'h17):(1'h0)] wire1385;
  input wire signed [(5'h12):(1'h0)] wire1384;
  reg [(2'h3):(1'h0)] reg1440 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1439 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1438 = (1'h0);
  reg [(3'h4):(1'h0)] reg1437 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1436 = (1'h0);
  reg [(4'h9):(1'h0)] reg1435 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1434 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1433 = (1'h0);
  reg [(3'h4):(1'h0)] reg1432 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1431 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1430 = (1'h0);
  reg [(5'h16):(1'h0)] reg1429 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1428 = (1'h0);
  reg [(5'h16):(1'h0)] reg1427 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1426 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1425 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1424 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1423 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1422 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1421 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1420 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1419 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1418 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1417 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1416 = (1'h0);
  reg [(2'h2):(1'h0)] reg1415 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1414 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1413 = (1'h0);
  reg [(4'hb):(1'h0)] reg1412 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1411 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1410 = (1'h0);
  reg [(4'h9):(1'h0)] reg1409 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1408 = (1'h0);
  reg [(3'h7):(1'h0)] reg1407 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1406 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1405 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1404 = (1'h0);
  reg [(5'h11):(1'h0)] reg1403 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1402 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1401 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1400 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1399 = (1'h0);
  reg [(5'h10):(1'h0)] reg1398 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1397 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1396 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1395 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire1394;
  reg [(2'h2):(1'h0)] reg1393 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1392 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1391 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1390 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1389 = (1'h0);
  reg [(4'hf):(1'h0)] reg1388 = (1'h0);
  assign y = {reg1440,
                 reg1439,
                 forvar1438,
                 reg1437,
                 reg1436,
                 reg1435,
                 reg1434,
                 reg1433,
                 reg1432,
                 forvar1431,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1427,
                 reg1426,
                 forvar1425,
                 forvar1424,
                 reg1423,
                 reg1422,
                 reg1421,
                 forvar1420,
                 forvar1419,
                 reg1418,
                 reg1417,
                 reg1416,
                 reg1415,
                 reg1414,
                 reg1413,
                 reg1412,
                 reg1411,
                 reg1410,
                 reg1409,
                 reg1408,
                 reg1407,
                 forvar1406,
                 forvar1405,
                 reg1404,
                 reg1403,
                 forvar1402,
                 reg1401,
                 reg1400,
                 forvar1399,
                 reg1398,
                 reg1397,
                 reg1396,
                 forvar1395,
                 wire1394,
                 reg1393,
                 reg1392,
                 reg1391,
                 reg1390,
                 reg1389,
                 reg1388,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1388 <= (7'h4c);
      reg1389 <= $signed($unsigned("COV0z4lH7UhG"));
      reg1390 <= $unsigned({"rl0RzTZwfUVviK", $signed(reg1389)});
      reg1391 <= {(wire1384 ?
              (reg1389[(3'h6):(2'h2)] << (((8'hb0) == reg1390) ^~ $unsigned(wire1386))) : wire1386[(2'h3):(2'h3)])};
      reg1392 <= $unsigned($signed(wire1384[(4'hc):(3'h7)]));
      reg1393 <= $signed(reg1390);
    end
  assign wire1394 = ($unsigned("") < ($unsigned((reg1392[(3'h4):(2'h3)] ?
                        reg1393 : (reg1388 ? reg1393 : reg1392))) >> reg1393));
  always
    @(posedge clk) begin
      for (forvar1395 = (1'h0); (forvar1395 < (1'h1)); forvar1395 = (forvar1395 + (1'h1)))
        begin
          reg1396 = "KcGtyi";
          reg1397 <= (~|$unsigned(reg1389));
          reg1398 = $unsigned("Y6SFZt");
        end
      for (forvar1399 = (1'h0); (forvar1399 < (1'h1)); forvar1399 = (forvar1399 + (1'h1)))
        begin
          reg1400 <= ($signed(($signed(forvar1395) ?
                  reg1398 : $signed((reg1392 ? reg1398 : forvar1395)))) ?
              reg1392 : (reg1390 ?
                  (^$unsigned((|reg1396))) : reg1390[(4'hc):(4'hc)]));
          reg1401 <= reg1389;
        end
    end
  always
    @(posedge clk) begin
      for (forvar1402 = (1'h0); (forvar1402 < (2'h3)); forvar1402 = (forvar1402 + (1'h1)))
        begin
          reg1403 <= "TVzRyz9";
          reg1404 <= {"5X5y63HZfB"};
          for (forvar1405 = (1'h0); (forvar1405 < (1'h1)); forvar1405 = (forvar1405 + (1'h1)))
            begin
              for (forvar1406 = (1'h0); (forvar1406 < (2'h2)); forvar1406 = (forvar1406 + (1'h1)))
                begin
                  reg1407 = "9yDDRZBsr0l";
                  reg1408 <= $unsigned(($unsigned($unsigned((~|wire1386))) ?
                      (wire1385[(4'hf):(3'h6)] ?
                          $signed(forvar1406[(3'h7):(1'h1)]) : $signed((reg1403 ?
                              reg1391 : reg1397))) : "S6O1Mg"));
                  reg1409 <= wire1387;
                  reg1410 = ($signed(reg1400[(2'h2):(1'h1)]) ~^ (8'hb9));
                end
            end
          reg1411 <= "pCw7VUGLZwAKwi0EKUo1Uf";
        end
      reg1412 <= reg1409[(4'h8):(3'h6)];
      reg1413 <= wire1387[(4'h8):(2'h3)];
      reg1414 <= $signed((^~($unsigned((forvar1395 - (8'hb0))) ?
          "WDEZZs3iCJd1nnK" : ("WFCYe24nDiB7lIygTbxpefGQ" << (reg1391 ?
              reg1412 : reg1392)))));
      reg1415 <= $signed(reg1412);
      reg1416 <= (&((reg1410 & reg1388[(1'h1):(1'h0)]) + reg1403));
    end
  always
    @(posedge clk) begin
      reg1417 <= ($signed(reg1411[(2'h2):(1'h1)]) ?
          $signed(((-reg1410) ?
              $signed(((8'h9e) ?
                  (8'hb3) : reg1390)) : ({reg1400} <= (reg1404 <= reg1398)))) : ({("g7GB2BK1R79M" ?
                      wire1385 : "2mSmrt5Ulr00y")} ?
              ("REskuo1L9mq" ?
                  ((8'hbf) ?
                      "8fA3VZyHFTfbLOpOqeUi3m" : reg1393) : forvar1406) : "6QL45GnI5l87f"));
      reg1418 = forvar1402;
    end
  always
    @(posedge clk) begin
      for (forvar1419 = (1'h0); (forvar1419 < (1'h1)); forvar1419 = (forvar1419 + (1'h1)))
        begin
          for (forvar1420 = (1'h0); (forvar1420 < (1'h1)); forvar1420 = (forvar1420 + (1'h1)))
            begin
              reg1421 = (~^$signed($unsigned((~|reg1389))));
              reg1422 <= ({"eYgd"} ^~ ((reg1412 ?
                      (reg1400[(1'h0):(1'h0)] ^ reg1414) : (~^reg1415)) ?
                  reg1391 : (reg1408[(2'h3):(2'h2)] ?
                      $signed("z9o74ykU5uFh1ysJIskG") : ($unsigned(forvar1406) * forvar1420[(1'h0):(1'h0)]))));
              reg1423 = $signed("4Mu");
            end
          for (forvar1424 = (1'h0); (forvar1424 < (1'h1)); forvar1424 = (forvar1424 + (1'h1)))
            begin
              for (forvar1425 = (1'h0); (forvar1425 < (3'h5)); forvar1425 = (forvar1425 + (1'h1)))
                begin
                  reg1426 <= reg1415;
                  reg1427 <= $unsigned({($unsigned("CasLgmyGP1wOctMSi5vr7gEB") || forvar1419),
                      $signed($unsigned($signed(wire1387)))});
                  reg1428 <= $signed((7'h47));
                  reg1429 <= "7n30wbVDbHkfnB5TFy";
                  reg1430 <= {$signed("YQuzXo"), reg1398};
                end
              for (forvar1431 = (1'h0); (forvar1431 < (3'h5)); forvar1431 = (forvar1431 + (1'h1)))
                begin
                  reg1432 <= (~&({$signed((+reg1408)),
                      $unsigned((~|reg1415))} ^ reg1417));
                end
              reg1433 <= ((({(~|reg1421)} < {reg1432[(2'h3):(1'h1)]}) >= $unsigned($signed((!reg1422)))) << "f");
              reg1434 <= reg1412;
              reg1435 <= "zhAM592Sgvxa";
            end
          reg1436 = $signed((^(~|{(&reg1414)})));
          reg1437 <= (wire1384 ? "KmNMFubF1" : reg1432[(1'h1):(1'h1)]);
          for (forvar1438 = (1'h0); (forvar1438 < (1'h1)); forvar1438 = (forvar1438 + (1'h1)))
            begin
              reg1439 <= (-forvar1402[(1'h0):(1'h0)]);
              reg1440 <= $unsigned($signed(forvar1424));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1146
#( parameter param1371 = ((~((((8'h9d) != (7'h43)) >= ((8'had) << (8'hbe))) * (((8'hac) ? (8'haa) : (7'h46)) ? ((7'h48) ? (8'had) : (7'h44)) : ((8'hbb) ? (8'hb0) : (8'ha2))))) ? {({((8'hba) ? (8'ha1) : (8'hb2))} <<< ({(8'hb8), (8'hab)} ? ((7'h44) ? (8'ha6) : (8'ha0)) : ((7'h45) ? (8'hb2) : (7'h4c))))} : ((&(~^((8'ha5) >>> (8'hb6)))) ? (~^((&(8'ha4)) != ((8'ha4) > (8'ha6)))) : ({((8'hba) == (8'ha5))} == {{(8'hab)}, (~|(8'hae))}))) )
(y, clk, wire1151, wire1150, wire1149, wire1148, wire1147);
  output wire [(32'hc1d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h19):(1'h0)] wire1151;
  input wire signed [(4'h8):(1'h0)] wire1150;
  input wire [(5'h14):(1'h0)] wire1149;
  input wire [(5'h17):(1'h0)] wire1148;
  input wire [(2'h3):(1'h0)] wire1147;
  reg signed [(5'h12):(1'h0)] reg1370 = (1'h0);
  reg [(5'h17):(1'h0)] reg1369 = (1'h0);
  reg [(5'h11):(1'h0)] reg1368 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1367 = (1'h0);
  reg [(4'hd):(1'h0)] reg1366 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1365 = (1'h0);
  reg [(2'h3):(1'h0)] reg1364 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1363 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar1362 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1361 = (1'h0);
  reg [(4'h9):(1'h0)] reg1360 = (1'h0);
  reg [(4'hd):(1'h0)] reg1359 = (1'h0);
  reg [(2'h2):(1'h0)] reg1358 = (1'h0);
  reg [(5'h13):(1'h0)] reg1357 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar1356 = (1'h0);
  reg [(3'h5):(1'h0)] reg1355 = (1'h0);
  reg [(5'h17):(1'h0)] reg1354 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1353 = (1'h0);
  reg [(4'h8):(1'h0)] reg1352 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1351 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1350 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1349 = (1'h0);
  reg [(5'h14):(1'h0)] reg1348 = (1'h0);
  reg [(4'he):(1'h0)] reg1347 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1346 = (1'h0);
  reg [(2'h2):(1'h0)] reg1345 = (1'h0);
  reg [(3'h6):(1'h0)] reg1344 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1343 = (1'h0);
  reg [(4'hc):(1'h0)] reg1342 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1341 = (1'h0);
  reg [(2'h3):(1'h0)] reg1340 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1339 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1338 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1337 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1336 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1335 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1334 = (1'h0);
  reg [(5'h12):(1'h0)] reg1333 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1332 = (1'h0);
  reg [(4'ha):(1'h0)] reg1331 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1330 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1329 = (1'h0);
  reg [(2'h2):(1'h0)] reg1328 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1327 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1326 = (1'h0);
  reg [(3'h5):(1'h0)] reg1325 = (1'h0);
  reg [(5'h17):(1'h0)] reg1324 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1323 = (1'h0);
  reg [(4'hf):(1'h0)] reg1322 = (1'h0);
  reg [(5'h12):(1'h0)] reg1321 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1320 = (1'h0);
  reg [(5'h13):(1'h0)] reg1319 = (1'h0);
  reg [(3'h5):(1'h0)] reg1318 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1317 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1316 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1315 = (1'h0);
  reg [(4'hb):(1'h0)] reg1314 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1313 = (1'h0);
  reg [(4'hd):(1'h0)] reg1312 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1311 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1310 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1309 = (1'h0);
  reg [(5'h18):(1'h0)] reg1308 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1307 = (1'h0);
  reg [(5'h14):(1'h0)] reg1306 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1305 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1304 = (1'h0);
  reg [(3'h5):(1'h0)] reg1303 = (1'h0);
  reg [(4'hd):(1'h0)] reg1302 = (1'h0);
  reg [(3'h6):(1'h0)] reg1301 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1300 = (1'h0);
  reg [(5'h11):(1'h0)] reg1299 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1298 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1297 = (1'h0);
  reg [(4'hf):(1'h0)] reg1296 = (1'h0);
  reg [(5'h11):(1'h0)] reg1295 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1294 = (1'h0);
  reg [(4'ha):(1'h0)] reg1293 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1292 = (1'h0);
  reg [(2'h2):(1'h0)] reg1291 = (1'h0);
  reg [(3'h4):(1'h0)] reg1290 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1289 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1288 = (1'h0);
  reg [(3'h6):(1'h0)] reg1287 = (1'h0);
  reg [(4'ha):(1'h0)] reg1286 = (1'h0);
  reg [(4'hf):(1'h0)] reg1285 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1284 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1283 = (1'h0);
  reg [(5'h14):(1'h0)] reg1282 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1281 = (1'h0);
  reg [(4'hc):(1'h0)] reg1280 = (1'h0);
  reg [(5'h13):(1'h0)] reg1279 = (1'h0);
  reg [(3'h5):(1'h0)] reg1278 = (1'h0);
  reg [(5'h11):(1'h0)] reg1277 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1276 = (1'h0);
  wire [(3'h4):(1'h0)] wire1275;
  reg [(5'h12):(1'h0)] reg1274 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1273 = (1'h0);
  reg [(3'h7):(1'h0)] reg1272 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1271 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1270 = (1'h0);
  reg [(3'h4):(1'h0)] reg1269 = (1'h0);
  reg [(5'h12):(1'h0)] reg1268 = (1'h0);
  reg [(2'h2):(1'h0)] reg1267 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1266 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1265 = (1'h0);
  reg [(2'h3):(1'h0)] reg1264 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1263 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1262 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1261 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1260 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1259 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1258 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1257 = (1'h0);
  reg [(3'h7):(1'h0)] reg1256 = (1'h0);
  reg [(4'h8):(1'h0)] reg1255 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1254 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1253 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1252 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1251 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1250 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1249 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1248 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1247 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1246 = (1'h0);
  reg [(3'h6):(1'h0)] reg1245 = (1'h0);
  reg [(4'hf):(1'h0)] reg1244 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1243 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1242 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1241 = (1'h0);
  reg [(4'he):(1'h0)] reg1240 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1239 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1238 = (1'h0);
  reg [(4'hf):(1'h0)] reg1237 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1236 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1235 = (1'h0);
  reg [(4'h9):(1'h0)] reg1234 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1233 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1232 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1231 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire1230;
  reg [(4'hb):(1'h0)] reg1229 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1228 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1227 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1226;
  reg signed [(4'hc):(1'h0)] reg1225 = (1'h0);
  wire signed [(5'h18):(1'h0)] wire1224;
  reg signed [(5'h18):(1'h0)] reg1223 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1222 = (1'h0);
  reg [(2'h2):(1'h0)] reg1221 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1220 = (1'h0);
  reg [(4'hf):(1'h0)] reg1219 = (1'h0);
  reg [(4'hb):(1'h0)] reg1218 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1217 = (1'h0);
  reg [(5'h16):(1'h0)] reg1216 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1215 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1214 = (1'h0);
  reg [(4'hf):(1'h0)] reg1213 = (1'h0);
  reg [(4'he):(1'h0)] reg1212 = (1'h0);
  reg [(5'h19):(1'h0)] reg1211 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1210 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1209 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1208 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1207 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1206 = (1'h0);
  reg [(4'ha):(1'h0)] reg1205 = (1'h0);
  reg [(3'h6):(1'h0)] reg1204 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1203 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1202 = (1'h0);
  reg [(3'h4):(1'h0)] reg1201 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1200 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1199 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1198 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1197 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1196 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1195 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1194 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1193 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1192 = (1'h0);
  reg [(5'h13):(1'h0)] reg1191 = (1'h0);
  reg [(4'ha):(1'h0)] reg1190 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1189 = (1'h0);
  reg [(5'h12):(1'h0)] reg1188 = (1'h0);
  reg [(4'h9):(1'h0)] reg1187 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1186 = (1'h0);
  reg [(5'h13):(1'h0)] reg1185 = (1'h0);
  reg [(5'h19):(1'h0)] reg1184 = (1'h0);
  reg [(5'h15):(1'h0)] reg1183 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire1182;
  reg [(4'h8):(1'h0)] reg1181 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1180 = (1'h0);
  reg [(4'hb):(1'h0)] reg1179 = (1'h0);
  reg [(5'h13):(1'h0)] reg1178 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1177 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1176 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1175 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1174 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1173 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1172 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1171 = (1'h0);
  reg [(5'h15):(1'h0)] reg1170 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1169 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1168 = (1'h0);
  reg [(5'h18):(1'h0)] reg1167 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1166 = (1'h0);
  reg [(5'h15):(1'h0)] reg1165 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1164 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1163 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1162 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1161 = (1'h0);
  reg [(4'h9):(1'h0)] reg1160 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1159 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1158 = (1'h0);
  reg [(2'h2):(1'h0)] reg1157 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1156 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1155 = (1'h0);
  reg [(5'h13):(1'h0)] reg1154 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1153 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire1152;
  assign y = {reg1370,
                 reg1369,
                 reg1368,
                 reg1367,
                 reg1366,
                 reg1365,
                 reg1364,
                 reg1363,
                 forvar1362,
                 reg1361,
                 reg1360,
                 reg1359,
                 reg1358,
                 reg1357,
                 forvar1356,
                 reg1355,
                 reg1354,
                 forvar1353,
                 reg1352,
                 reg1351,
                 reg1350,
                 reg1349,
                 reg1348,
                 reg1347,
                 forvar1346,
                 reg1345,
                 reg1344,
                 reg1343,
                 reg1342,
                 forvar1341,
                 reg1340,
                 reg1339,
                 reg1338,
                 reg1337,
                 reg1336,
                 reg1335,
                 reg1334,
                 reg1333,
                 reg1332,
                 reg1331,
                 forvar1330,
                 forvar1329,
                 reg1328,
                 reg1327,
                 forvar1326,
                 reg1325,
                 reg1324,
                 reg1323,
                 reg1322,
                 reg1321,
                 reg1320,
                 reg1319,
                 reg1318,
                 forvar1317,
                 reg1316,
                 reg1315,
                 reg1314,
                 reg1313,
                 reg1312,
                 reg1311,
                 forvar1310,
                 forvar1309,
                 reg1308,
                 reg1307,
                 reg1306,
                 reg1305,
                 reg1304,
                 reg1303,
                 reg1302,
                 reg1301,
                 reg1300,
                 reg1299,
                 reg1298,
                 forvar1297,
                 reg1296,
                 reg1295,
                 reg1294,
                 reg1293,
                 forvar1292,
                 reg1291,
                 reg1290,
                 reg1289,
                 reg1288,
                 reg1287,
                 reg1286,
                 reg1285,
                 forvar1284,
                 reg1283,
                 reg1282,
                 forvar1281,
                 reg1280,
                 reg1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 wire1275,
                 reg1274,
                 reg1273,
                 reg1272,
                 reg1271,
                 forvar1270,
                 reg1269,
                 reg1268,
                 reg1267,
                 reg1266,
                 forvar1265,
                 reg1264,
                 reg1263,
                 reg1262,
                 reg1261,
                 reg1260,
                 reg1259,
                 reg1258,
                 reg1257,
                 reg1256,
                 reg1255,
                 reg1254,
                 forvar1253,
                 reg1252,
                 forvar1251,
                 reg1250,
                 reg1249,
                 reg1248,
                 reg1247,
                 reg1246,
                 reg1245,
                 reg1244,
                 reg1243,
                 reg1242,
                 reg1241,
                 reg1240,
                 forvar1239,
                 reg1238,
                 reg1237,
                 reg1236,
                 reg1235,
                 reg1234,
                 forvar1233,
                 forvar1232,
                 reg1231,
                 wire1230,
                 reg1229,
                 reg1228,
                 reg1227,
                 wire1226,
                 reg1225,
                 wire1224,
                 reg1223,
                 reg1222,
                 reg1221,
                 forvar1220,
                 reg1219,
                 reg1218,
                 reg1217,
                 reg1216,
                 reg1215,
                 reg1214,
                 reg1213,
                 reg1212,
                 reg1211,
                 reg1210,
                 reg1209,
                 reg1208,
                 reg1207,
                 reg1206,
                 reg1205,
                 reg1204,
                 reg1203,
                 reg1202,
                 reg1201,
                 reg1200,
                 reg1199,
                 reg1198,
                 forvar1197,
                 reg1196,
                 forvar1195,
                 reg1194,
                 forvar1193,
                 reg1192,
                 reg1191,
                 reg1190,
                 reg1189,
                 reg1188,
                 reg1187,
                 forvar1186,
                 reg1185,
                 reg1184,
                 reg1183,
                 wire1182,
                 reg1181,
                 reg1180,
                 reg1179,
                 reg1178,
                 forvar1177,
                 forvar1176,
                 reg1175,
                 reg1174,
                 reg1173,
                 reg1172,
                 reg1171,
                 reg1170,
                 forvar1169,
                 reg1168,
                 reg1167,
                 reg1166,
                 reg1165,
                 reg1164,
                 reg1163,
                 reg1162,
                 reg1161,
                 reg1160,
                 forvar1159,
                 reg1158,
                 reg1157,
                 forvar1156,
                 reg1155,
                 reg1154,
                 forvar1153,
                 wire1152,
                 (1'h0)};
  assign wire1152 = wire1148[(5'h15):(5'h13)];
  always
    @(posedge clk) begin
      for (forvar1153 = (1'h0); (forvar1153 < (1'h0)); forvar1153 = (forvar1153 + (1'h1)))
        begin
          reg1154 = ($unsigned(wire1151[(3'h7):(3'h4)]) & wire1150[(3'h6):(2'h2)]);
          reg1155 <= (^~$unsigned(((((8'ha7) ?
              forvar1153 : wire1147) * (wire1148 < forvar1153)) >= "")));
          for (forvar1156 = (1'h0); (forvar1156 < (1'h0)); forvar1156 = (forvar1156 + (1'h1)))
            begin
              reg1157 <= {reg1155, wire1150};
              reg1158 <= $unsigned($unsigned(wire1150));
              for (forvar1159 = (1'h0); (forvar1159 < (3'h4)); forvar1159 = (forvar1159 + (1'h1)))
                begin
                  reg1160 <= wire1149[(1'h1):(1'h1)];
                  reg1161 = "phUMEwZ1";
                  reg1162 <= wire1150[(3'h5):(2'h3)];
                end
              reg1163 <= (((reg1160[(2'h2):(2'h2)] * ("mkxY4hS" ^~ (reg1162 != wire1147))) && (wire1152 & ((reg1160 >>> reg1154) >> (8'ha5)))) >>> (forvar1159[(3'h7):(3'h6)] ?
                  ($unsigned((~&(8'hb0))) != (reg1155 - $signed(wire1150))) : forvar1153));
              if ((|forvar1159[(4'h8):(1'h1)]))
                begin
                  reg1164 <= "wrIcbfQOWA4";
                end
              else
                begin
                  reg1164 <= "DcRM1GO6MDsC2yeQMmT5x";
                  reg1165 <= (|(-{$unsigned((wire1150 & wire1149)),
                      "WRSlIyeXwTlvf5fGTQvW6"}));
                  reg1166 <= ("ZQvwKmp9ngOQAdHFDSs" ^ (&(reg1154[(4'hd):(4'ha)] ?
                      $unsigned($signed(wire1147)) : $unsigned(wire1151))));
                  reg1167 = (+("DShU9RaOe5DRZVqx" ?
                      reg1154[(4'h8):(2'h3)] : ($unsigned({(7'h42)}) ?
                          $unsigned($signed(reg1154)) : reg1163)));
                  reg1168 <= (8'hbc);
                end
              for (forvar1169 = (1'h0); (forvar1169 < (2'h2)); forvar1169 = (forvar1169 + (1'h1)))
                begin
                  reg1170 <= reg1163;
                  reg1171 <= "Y8kJaM2MztpDJ3UiWB";
                  reg1172 = $unsigned(reg1154);
                end
            end
        end
      reg1173 = (($unsigned((~&{reg1167})) ^ $signed(wire1150)) ?
          $signed((reg1171 ?
              $signed((!(8'h9c))) : $unsigned((reg1166 ?
                  reg1166 : (8'haf))))) : (~&wire1148[(4'ha):(2'h3)]));
      reg1174 <= (8'ha8);
      reg1175 <= (reg1166[(1'h0):(1'h0)] ?
          $unsigned("HKU96T637") : ($unsigned({(reg1171 ?
                      forvar1153 : wire1148),
                  (8'h9c)}) ?
              $unsigned(reg1174) : $signed($unsigned((reg1167 <<< forvar1156)))));
      for (forvar1176 = (1'h0); (forvar1176 < (3'h5)); forvar1176 = (forvar1176 + (1'h1)))
        begin
          for (forvar1177 = (1'h0); (forvar1177 < (2'h2)); forvar1177 = (forvar1177 + (1'h1)))
            begin
              reg1178 <= (reg1167[(4'h8):(1'h1)] ?
                  (-$signed({(~&wire1150)})) : reg1165);
            end
          reg1179 = ($unsigned($unsigned(wire1151[(5'h16):(4'h8)])) * "kP4mCSl5Lrw");
          reg1180 <= $signed(wire1149);
          reg1181 = reg1155[(1'h0):(1'h0)];
        end
    end
  assign wire1182 = (reg1172[(3'h7):(3'h7)] ?
                        $signed("8FmHJiaM8n") : ($signed((|wire1149[(2'h2):(2'h2)])) ?
                            reg1161 : reg1167));
  always
    @(posedge clk) begin
      if ("25NfNLQxk")
        begin
          reg1183 = ($unsigned((~&{$signed(reg1160)})) >> (~&(|$unsigned($signed(reg1180)))));
          reg1184 <= reg1155;
          reg1185 <= $unsigned(("bT" | (~^($signed(reg1158) ?
              ((8'ha9) ? reg1168 : reg1175) : "r2ZBnTriRV"))));
        end
      else
        begin
          reg1183 <= ((|$signed((!{(8'hac), reg1179}))) ?
              $unsigned((-(forvar1153 > (reg1167 ?
                  reg1154 : reg1180)))) : {(^(+$signed((8'ha3))))});
          reg1184 = reg1183;
          reg1185 <= forvar1156;
          for (forvar1186 = (1'h0); (forvar1186 < (3'h5)); forvar1186 = (forvar1186 + (1'h1)))
            begin
              reg1187 <= ($signed(reg1168) ?
                  $unsigned((wire1151[(4'hb):(3'h5)] >>> ($signed(reg1157) << {reg1172}))) : $unsigned(("c2z1avLyK3yw" + $unsigned(forvar1176[(3'h6):(1'h0)]))));
              reg1188 = "9EEa7NOQyt5";
            end
          reg1189 <= {"Cb2n2RD6a65XktFXkGxzB"};
        end
      reg1190 <= ("yWRWq9kZypT" ?
          reg1164 : ($signed((~|((7'h45) & reg1155))) ?
              "kMTYuUPcRZ" : wire1152[(4'h8):(2'h3)]));
      reg1191 = "vA0T";
      reg1192 <= reg1175;
      for (forvar1193 = (1'h0); (forvar1193 < (1'h0)); forvar1193 = (forvar1193 + (1'h1)))
        begin
          reg1194 = wire1182[(2'h3):(1'h1)];
          for (forvar1195 = (1'h0); (forvar1195 < (2'h2)); forvar1195 = (forvar1195 + (1'h1)))
            begin
              reg1196 <= reg1191[(4'he):(2'h2)];
              for (forvar1197 = (1'h0); (forvar1197 < (2'h3)); forvar1197 = (forvar1197 + (1'h1)))
                begin
                  reg1198 <= reg1167;
                  reg1199 = (7'h40);
                  reg1200 = "cdf6XwB2JM3";
                  reg1201 <= (|{$unsigned("W8Y23dLrGRkofhkx83rk2SpKy"),
                      (&{reg1184, $signed(reg1166)})});
                  reg1202 <= (reg1155 > reg1165[(3'h4):(3'h4)]);
                end
              reg1203 <= (reg1170[(1'h1):(1'h0)] << reg1157[(1'h1):(1'h0)]);
              reg1204 = (-"NwI5C7Zy5");
              reg1205 <= (+$signed($unsigned(reg1196[(4'h9):(3'h5)])));
            end
          reg1206 <= reg1173[(1'h0):(1'h0)];
          reg1207 <= "YgOPYnLRG88sfXdXkAe4";
          reg1208 <= reg1187;
          reg1209 <= "";
        end
    end
  always
    @(posedge clk) begin
      reg1210 = ({(wire1150[(3'h5):(2'h3)] | reg1172[(1'h1):(1'h1)])} > $unsigned({wire1182[(4'hc):(4'hc)]}));
    end
  always
    @(posedge clk) begin
      reg1211 <= reg1165[(5'h13):(3'h5)];
    end
  always
    @(posedge clk) begin
      reg1212 = $signed(reg1194);
      reg1213 <= {{$signed({"hEFUryIhkHM0sVUw", ((7'h49) * wire1149)})}};
      reg1214 <= reg1174;
      reg1215 <= (((!($signed(forvar1186) ^~ $unsigned((8'h9f)))) ?
              {reg1190} : forvar1193[(2'h3):(2'h3)]) ?
          (reg1199[(4'ha):(2'h3)] ?
              "2dpxqi2PMp3pXVxxzyeNTh" : reg1188[(3'h7):(3'h5)]) : (~^(^~((~|reg1178) ?
              wire1151 : $signed(reg1166)))));
    end
  always
    @(posedge clk) begin
      reg1216 <= "pTIhfxyhHIntkKHJnJ7GybDUE";
      reg1217 <= "";
      reg1218 <= reg1212[(4'hc):(1'h1)];
      reg1219 <= ($signed((|$signed((forvar1186 * forvar1177)))) ~^ {$signed($unsigned(((8'hb6) ?
              reg1217 : wire1150)))});
      for (forvar1220 = (1'h0); (forvar1220 < (3'h5)); forvar1220 = (forvar1220 + (1'h1)))
        begin
          reg1221 <= {($unsigned(reg1180[(1'h0):(1'h0)]) ^~ "W"),
              $signed({(((8'had) ? reg1214 : reg1191) ?
                      $signed(reg1163) : (&reg1172))})};
        end
      reg1222 <= "zBxpeg";
    end
  always
    @(posedge clk) begin
      reg1223 = $unsigned(({($unsigned(reg1168) ^~ $signed(reg1173)),
              $unsigned($signed(reg1162))} ?
          reg1167 : ($unsigned(reg1155) - (~reg1194[(4'hd):(4'h8)]))));
    end
  assign wire1224 = (~$unsigned(forvar1156[(1'h1):(1'h0)]));
  always
    @(posedge clk) begin
      reg1225 <= "5NanlXI1Us6aDYFB45O";
    end
  assign wire1226 = "PsLPKEyOp9qT4p4326H7oCGft";
  always
    @(posedge clk) begin
      reg1227 <= $signed((reg1206 >= $signed({forvar1153[(4'h9):(3'h7)]})));
      reg1228 <= $signed(({($signed(reg1178) ? "Phd94Srk7qeD4El7" : (+reg1181)),
              ($signed((8'hb5)) || $signed(reg1222))} ?
          (reg1157 != reg1211) : $signed($unsigned({reg1206, forvar1159}))));
      reg1229 <= forvar1186[(1'h1):(1'h1)];
    end
  assign wire1230 = ((((reg1198 <<< reg1188[(1'h0):(1'h0)]) ?
                        reg1225[(1'h1):(1'h0)] : wire1149) == $signed((-(^reg1201)))) << {"nD8aUtHe73Vo",
                        reg1210});
  always
    @(posedge clk) begin
      reg1231 <= (8'ha2);
      for (forvar1232 = (1'h0); (forvar1232 < (1'h1)); forvar1232 = (forvar1232 + (1'h1)))
        begin
          for (forvar1233 = (1'h0); (forvar1233 < (3'h4)); forvar1233 = (forvar1233 + (1'h1)))
            begin
              reg1234 = ((^$signed((~&$signed((8'haa))))) * "Lo7xl58BQPx");
              reg1235 <= wire1230;
              reg1236 = (^{{((~&(7'h4e)) ? (forvar1197 + wire1147) : reg1158)},
                  reg1202[(2'h2):(1'h1)]});
              reg1237 <= (|wire1152[(4'ha):(4'ha)]);
              reg1238 <= ({reg1207} ?
                  $signed(reg1210[(5'h15):(3'h6)]) : ((reg1172 <= "5CINcNuJXaTcZieneIGC5EiT") ?
                      $signed(reg1203) : (8'hac)));
              for (forvar1239 = (1'h0); (forvar1239 < (3'h4)); forvar1239 = (forvar1239 + (1'h1)))
                begin
                  reg1240 <= "l3ZOmGeV0VPya057LcAB";
                  reg1241 = $signed(reg1200);
                  reg1242 <= reg1227[(3'h7):(1'h0)];
                  reg1243 <= (!"hpFsKGaC8o");
                  reg1244 <= (^"LtJH2Ixm8fO8dgVw9wsiW");
                end
            end
          reg1245 <= (^~"aEmOu");
          reg1246 <= $unsigned({{$signed((reg1196 ~^ reg1237)),
                  (!"HCEp71EZvUYy6dJfd5lZvX2")},
              $unsigned(reg1174[(2'h2):(2'h2)])});
        end
    end
  always
    @(posedge clk) begin
      reg1247 <= reg1196[(3'h7):(2'h3)];
      reg1248 <= forvar1186;
      reg1249 <= (reg1154 ? reg1246 : $signed($signed(reg1168[(4'he):(4'hc)])));
      reg1250 = "wtU1bPAlGMzT4TIB4kxJeCD";
    end
  always
    @(posedge clk) begin
      for (forvar1251 = (1'h0); (forvar1251 < (2'h2)); forvar1251 = (forvar1251 + (1'h1)))
        begin
          reg1252 <= $signed({reg1183[(1'h1):(1'h0)]});
          for (forvar1253 = (1'h0); (forvar1253 < (2'h3)); forvar1253 = (forvar1253 + (1'h1)))
            begin
              reg1254 <= (~"N7tOSLT");
              reg1255 <= {"9vnZk"};
              reg1256 = forvar1156;
              reg1257 <= (8'ha6);
              reg1258 = $unsigned("6gPV");
              reg1259 = ("wHftCrCX4uw08" ~^ reg1198);
            end
          reg1260 = "";
        end
    end
  always
    @(posedge clk) begin
      reg1261 <= ("2kiZsIOSK10JmXMhzvLztZ1p" <= (forvar1233 ^~ $unsigned((8'hb0))));
      reg1262 <= forvar1153[(4'h8):(1'h0)];
      reg1263 = reg1255[(4'h8):(2'h2)];
      reg1264 = reg1258[(2'h3):(1'h0)];
      for (forvar1265 = (1'h0); (forvar1265 < (1'h0)); forvar1265 = (forvar1265 + (1'h1)))
        begin
          reg1266 = {(($signed(reg1191[(4'ha):(3'h4)]) ?
                      {$unsigned(forvar1186),
                          forvar1265[(3'h5):(2'h3)]} : reg1191[(5'h10):(2'h2)]) ?
                  (~|(~|reg1178)) : (({forvar1220, wire1182} ?
                      reg1235[(4'h9):(3'h4)] : "kNSfqSJANLqNAQk8wi8ex8Y") <= (~&"0")))};
          reg1267 <= ((^("Cgq" | "WhrpiKGBW8nrd3mbdd5Zn4")) >> (~($unsigned(reg1260) ?
              (~^forvar1232) : (-(reg1260 >= reg1216)))));
          reg1268 = ((|$signed($unsigned("XueHricuS6K"))) < $unsigned((({reg1211} || {reg1164}) & $unsigned(forvar1153))));
          reg1269 <= ((^wire1226) ?
              reg1154 : ($unsigned(({(7'h4d), reg1222} ?
                      $signed(reg1163) : "kpKdOEqNhWx9ZmCO4wpKDwze")) ?
                  reg1231[(5'h11):(5'h10)] : (((8'hbd) ?
                      (reg1267 >= reg1189) : $signed(reg1240)) * (~|$unsigned(reg1178)))));
          for (forvar1270 = (1'h0); (forvar1270 < (3'h4)); forvar1270 = (forvar1270 + (1'h1)))
            begin
              reg1271 <= (-reg1249[(3'h5):(3'h5)]);
              reg1272 <= $signed(reg1264);
              reg1273 <= ((($signed((reg1188 + forvar1239)) ?
                      (8'ha8) : (&reg1250)) ?
                  ((+(!reg1223)) >= "ACSV") : reg1206[(5'h12):(4'hf)]) ^ reg1162);
            end
        end
      reg1274 = (8'ha7);
    end
  assign wire1275 = "Op6RHNpC50ntFlRIg";
  always
    @(posedge clk) begin
      reg1276 = ($unsigned($unsigned($signed((reg1249 | (8'hae))))) != "aoFqzRbwW8ypxlPYp");
      reg1277 <= forvar1253[(1'h0):(1'h0)];
      reg1278 <= $signed($signed(($unsigned(reg1269[(2'h2):(1'h0)]) ?
          {$signed(reg1262), reg1252} : reg1213[(3'h4):(1'h0)])));
      reg1279 <= reg1210[(3'h4):(2'h3)];
      reg1280 <= $unsigned($signed((8'hb6)));
      for (forvar1281 = (1'h0); (forvar1281 < (1'h1)); forvar1281 = (forvar1281 + (1'h1)))
        begin
          reg1282 <= (-($unsigned(($signed(reg1261) <= (~|reg1198))) ?
              reg1267 : (&((!(7'h49)) << reg1208[(1'h0):(1'h0)]))));
          reg1283 = reg1200;
          for (forvar1284 = (1'h0); (forvar1284 < (3'h5)); forvar1284 = (forvar1284 + (1'h1)))
            begin
              reg1285 <= $signed((&$unsigned(reg1157)));
            end
          reg1286 <= ((("IP6meHVT7g3nsfpa" << reg1162[(5'h11):(4'h9)]) ?
              $signed("v1dvFWMMSGWZYs") : $signed(reg1268[(3'h6):(2'h2)])) || ($signed((^(+(7'h4b)))) ^~ reg1205[(4'h8):(1'h0)]));
          reg1287 <= $unsigned((|"u2KSC9FawUNis18KOhZKaet"));
        end
    end
  always
    @(posedge clk) begin
      reg1288 = $unsigned(((8'hbb) ? "M0840OxzufgPL9xeQz" : (7'h42)));
      reg1289 <= forvar1159[(4'h9):(3'h4)];
      reg1290 <= $unsigned((~$signed(((reg1243 & reg1231) << wire1150))));
      reg1291 <= {$unsigned(reg1158)};
      for (forvar1292 = (1'h0); (forvar1292 < (2'h3)); forvar1292 = (forvar1292 + (1'h1)))
        begin
          reg1293 <= (~|{"S8"});
          reg1294 <= (reg1240 >= ((^((forvar1176 ? reg1180 : forvar1193) ?
              reg1221[(1'h0):(1'h0)] : (reg1238 ?
                  reg1194 : reg1250))) + $unsigned(wire1226[(1'h1):(1'h1)])));
          reg1295 <= (!reg1277[(4'hd):(2'h2)]);
        end
      reg1296 <= "JOy4ET9VAmQoou1X23HilfN";
    end
  always
    @(posedge clk) begin
      for (forvar1297 = (1'h0); (forvar1297 < (3'h5)); forvar1297 = (forvar1297 + (1'h1)))
        begin
          reg1298 = ($unsigned(reg1164[(3'h6):(3'h4)]) * (^~({(reg1285 ?
                      reg1221 : reg1266),
                  reg1269} ?
              ($signed(forvar1251) ?
                  $signed(forvar1220) : (reg1185 ?
                      forvar1153 : reg1243)) : reg1267[(2'h2):(2'h2)])));
        end
      reg1299 <= $signed($signed(($signed("Yd5VUTTgX") ^ $signed(reg1269[(1'h0):(1'h0)]))));
      reg1300 <= ("VAaUQzwgv1p" && reg1279[(3'h6):(2'h2)]);
      reg1301 = reg1207;
      reg1302 <= reg1269;
      reg1303 <= $signed(($unsigned(reg1194[(3'h4):(1'h0)]) ?
          (((reg1276 ^~ reg1287) ?
              $signed(reg1212) : (wire1182 + reg1295)) | ((reg1234 ?
              wire1275 : forvar1197) > (reg1240 ~^ reg1215))) : reg1208[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg1304 <= "o";
      reg1305 = reg1264[(1'h1):(1'h0)];
      reg1306 = (reg1210[(5'h10):(4'hb)] || "CiZ4ZzU");
      reg1307 <= (|($signed(forvar1159) ?
          reg1154[(5'h13):(2'h3)] : (reg1179 >> (~^reg1296[(3'h4):(3'h4)]))));
      reg1308 <= (reg1241 != ((~(wire1151 ^ (forvar1265 ?
          reg1264 : reg1302))) && (reg1234 | forvar1233)));
    end
  always
    @(posedge clk) begin
      for (forvar1309 = (1'h0); (forvar1309 < (1'h0)); forvar1309 = (forvar1309 + (1'h1)))
        begin
          for (forvar1310 = (1'h0); (forvar1310 < (1'h1)); forvar1310 = (forvar1310 + (1'h1)))
            begin
              reg1311 = "";
              if ($signed($signed("aREd5tHzkeFiKLsNDYc")))
                begin
                  reg1312 = {(!reg1180[(4'h8):(3'h6)])};
                  reg1313 <= (reg1185[(4'hf):(4'ha)] ?
                      reg1223[(3'h6):(1'h0)] : (reg1199[(3'h6):(2'h2)] << $unsigned((^(-reg1308)))));
                end
              else
                begin
                  reg1312 <= (~&(reg1301[(2'h2):(2'h2)] || "E1"));
                  reg1313 <= ($signed(("Y2" ?
                          (^reg1264) : ("S" ?
                              ((8'hb0) ?
                                  reg1305 : (8'ha8)) : $unsigned(reg1269)))) ?
                      "NP0bAscu07K4JgXiaSCvuN" : "U");
                  reg1314 <= reg1234[(3'h7):(1'h1)];
                  reg1315 <= {$unsigned($signed(reg1272)), {"iS02"}};
                  reg1316 = {(^(-(~|"VE4pefUHC4AaMYizpzwe")))};
                end
            end
          for (forvar1317 = (1'h0); (forvar1317 < (3'h4)); forvar1317 = (forvar1317 + (1'h1)))
            begin
              reg1318 <= $unsigned({{{(reg1261 ? reg1158 : (8'hb4)),
                          "JWs7ff7xpcOAnTrfpc"},
                      (~&(~&(8'hbc)))},
                  "A"});
              reg1319 <= reg1173;
              reg1320 = $unsigned(reg1312[(3'h7):(2'h3)]);
              reg1321 = forvar1251[(1'h1):(1'h0)];
            end
          reg1322 = $unsigned((reg1271 ?
              (&$signed(((7'h4a) ?
                  reg1206 : reg1315))) : reg1307[(4'hc):(4'h8)]));
          reg1323 <= (7'h45);
          reg1324 = (reg1305 <= ($signed({forvar1197}) >>> "4MuYU"));
          reg1325 <= (7'h42);
        end
    end
  always
    @(posedge clk) begin
      for (forvar1326 = (1'h0); (forvar1326 < (3'h5)); forvar1326 = (forvar1326 + (1'h1)))
        begin
          reg1327 <= "H1yu51";
        end
      reg1328 = (((-$signed(reg1240[(4'hc):(4'hb)])) ?
              "YdC3pVoskEHJYM" : "Jc0DHE8b2eOS") ?
          reg1237[(3'h6):(2'h3)] : (7'h4b));
      for (forvar1329 = (1'h0); (forvar1329 < (1'h0)); forvar1329 = (forvar1329 + (1'h1)))
        begin
          for (forvar1330 = (1'h0); (forvar1330 < (3'h4)); forvar1330 = (forvar1330 + (1'h1)))
            begin
              reg1331 <= ($unsigned(reg1249) << ({((reg1299 ?
                          reg1174 : wire1275) ?
                      $unsigned(reg1302) : (+reg1208))} | $unsigned("dagvVgpKuI3U68RnPlT")));
              if (($unsigned((^{(reg1215 ? (7'h49) : reg1252),
                      {reg1257, reg1168}})) ?
                  $unsigned({"b52zDcbMCqSkJC",
                      $signed(((8'hb2) ?
                          reg1218 : reg1321))}) : ((&($unsigned(reg1166) == $unsigned(reg1258))) ?
                      reg1207[(5'h17):(1'h1)] : $unsigned(reg1194[(4'hd):(1'h0)]))))
                begin
                  reg1332 <= ($unsigned((~reg1264[(1'h0):(1'h0)])) != "PDVV2hCBdbsBzsnVEqkIkpdQX");
                  reg1333 <= ($signed(reg1246[(3'h5):(1'h1)]) ?
                      reg1183 : forvar1239);
                  reg1334 <= (~^forvar1292);
                  reg1335 <= reg1266[(2'h2):(2'h2)];
                  reg1336 = wire1150[(3'h5):(2'h2)];
                end
              else
                begin
                  reg1332 <= (!wire1226);
                  reg1333 <= $signed((("nOA6ggIhvWhAa8qSDhozWt" == ((wire1182 == reg1274) ?
                          reg1234[(2'h2):(2'h2)] : reg1321[(4'he):(2'h3)])) ?
                      $signed($unsigned($unsigned(reg1166))) : $signed($signed((+reg1313)))));
                  reg1334 <= ((^~$unsigned((reg1231[(5'h11):(5'h10)] ?
                      ((7'h46) ?
                          forvar1239 : wire1275) : (~&reg1242)))) >= reg1268);
                end
              reg1337 <= reg1321;
              reg1338 <= $unsigned("ybownOW");
            end
          reg1339 <= {reg1181};
        end
      reg1340 <= reg1331[(2'h3):(2'h2)];
      for (forvar1341 = (1'h0); (forvar1341 < (1'h1)); forvar1341 = (forvar1341 + (1'h1)))
        begin
          reg1342 <= (!"LtATcimPB5QlCzqSz");
          reg1343 = $unsigned(reg1274);
          reg1344 = $unsigned((8'ha9));
          reg1345 <= (reg1268 ?
              forvar1329 : (("uVvMnFiux" ?
                      reg1225[(4'hb):(1'h1)] : (~&(reg1207 < wire1148))) ?
                  $unsigned(((reg1245 ? reg1282 : wire1150) ?
                      "EYGtM1vF09" : reg1171)) : $unsigned((&$signed(reg1227)))));
          for (forvar1346 = (1'h0); (forvar1346 < (3'h5)); forvar1346 = (forvar1346 + (1'h1)))
            begin
              reg1347 <= reg1248;
              reg1348 <= "Ch";
              reg1349 <= {$unsigned(reg1287)};
              reg1350 <= reg1261[(3'h7):(2'h3)];
              reg1351 <= wire1150[(1'h0):(1'h0)];
              reg1352 <= (~^({reg1184[(4'he):(4'he)],
                  {(reg1351 ?
                          (8'hae) : reg1165)}} ^~ $signed((reg1318[(2'h3):(2'h2)] >> (reg1320 ?
                  wire1230 : reg1262)))));
            end
          for (forvar1353 = (1'h0); (forvar1353 < (3'h5)); forvar1353 = (forvar1353 + (1'h1)))
            begin
              reg1354 <= ($unsigned(reg1168[(2'h3):(2'h3)]) ?
                  $unsigned((((reg1321 ? reg1335 : reg1335) - "2at") ?
                      $signed(reg1170[(4'hd):(4'h8)]) : ("JNlmFkJf8YdyE3IVm7" ~^ reg1301[(3'h4):(2'h3)]))) : (7'h4c));
              reg1355 = (($signed((reg1345 ^~ (reg1189 ~^ reg1305))) | wire1224[(3'h7):(1'h1)]) ?
                  reg1332 : (&reg1305[(1'h1):(1'h1)]));
              for (forvar1356 = (1'h0); (forvar1356 < (1'h0)); forvar1356 = (forvar1356 + (1'h1)))
                begin
                  reg1357 <= ($unsigned($unsigned((~&$signed(reg1271)))) ?
                      wire1149 : $unsigned((7'h44)));
                  reg1358 <= (forvar1186 ?
                      (+"4hYfKBSQ04iZ") : (($unsigned({forvar1317}) ?
                          $signed("QIY55ECLKYP") : (reg1274 ?
                              (~reg1179) : $signed(reg1319))) + (reg1237[(4'hb):(3'h5)] ?
                          {$signed(forvar1281)} : $unsigned($signed(reg1298)))));
                  reg1359 <= "";
                  reg1360 <= $signed(reg1168);
                  reg1361 <= "r8scqfsH7";
                end
              for (forvar1362 = (1'h0); (forvar1362 < (2'h2)); forvar1362 = (forvar1362 + (1'h1)))
                begin
                  reg1363 <= reg1299;
                  reg1364 <= (({forvar1232[(1'h1):(1'h1)],
                              (-(reg1173 ? reg1168 : (7'h46)))} ?
                          ("EasGrZDOJWAh0OsW0ZoBd2w" ?
                              reg1293[(3'h7):(3'h4)] : "X1kLvvL") : ({(reg1198 ?
                                      reg1335 : reg1255),
                                  reg1254[(5'h13):(4'hd)]} ?
                              {reg1248[(4'h8):(2'h3)],
                                  (reg1332 < reg1296)} : reg1215[(2'h3):(1'h0)])) ?
                      "" : {(!$signed((reg1228 ? forvar1239 : reg1223))),
                          {forvar1310[(4'hf):(4'he)]}});
                  reg1365 = $unsigned((($unsigned($signed(wire1147)) ?
                      ((~^reg1219) + $signed(reg1347)) : reg1243[(3'h4):(2'h3)]) > reg1242));
                  reg1366 = (-(reg1334 ~^ {$unsigned(reg1217),
                      $unsigned("m2cnpnqUQUsL8")}));
                  reg1367 <= reg1191[(4'hf):(4'hb)];
                end
              reg1368 <= $signed(reg1339);
              reg1369 = (reg1190 > $signed((!(reg1300 == reg1218))));
            end
        end
      reg1370 = (((&$signed((reg1228 ?
          forvar1362 : reg1171))) != reg1178) - reg1179[(4'h8):(3'h5)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module957
#( parameter param1142 = {(!((~^(-(8'ha1))) ? (((7'h42) ? (7'h48) : (7'h4d)) ? (~^(8'haf)) : ((8'hbd) ? (8'ha2) : (8'hb3))) : (((8'haa) >>> (8'ha3)) | (+(8'haa)))))}
, parameter param1143 = ((~((!(param1142 ? (8'ha9) : param1142)) && param1142)) ? param1142 : (+(+param1142))) )
(y, clk, wire962, wire961, wire960, wire959, wire958);
  output wire [(32'h936):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire962;
  input wire signed [(5'h14):(1'h0)] wire961;
  input wire signed [(5'h14):(1'h0)] wire960;
  input wire [(4'hd):(1'h0)] wire959;
  input wire [(4'h8):(1'h0)] wire958;
  reg [(4'ha):(1'h0)] reg1141 = (1'h0);
  reg [(4'h9):(1'h0)] reg1140 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1139 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1138 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1137 = (1'h0);
  reg [(4'hf):(1'h0)] reg1136 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire1135;
  reg [(4'hc):(1'h0)] reg1134 = (1'h0);
  reg [(5'h10):(1'h0)] reg1133 = (1'h0);
  reg [(4'hf):(1'h0)] reg1132 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1131 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire1130;
  wire [(5'h16):(1'h0)] wire1129;
  wire [(5'h11):(1'h0)] wire1128;
  reg signed [(3'h5):(1'h0)] reg1127 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1126 = (1'h0);
  reg [(4'hd):(1'h0)] reg1125 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1124 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1123 = (1'h0);
  reg [(5'h16):(1'h0)] reg1122 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1121 = (1'h0);
  reg [(3'h6):(1'h0)] reg1120 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1119 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1118 = (1'h0);
  reg [(3'h4):(1'h0)] reg1117 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1116 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1115 = (1'h0);
  reg [(5'h19):(1'h0)] reg1114 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1113 = (1'h0);
  reg [(4'hf):(1'h0)] reg1112 = (1'h0);
  reg [(4'hf):(1'h0)] reg1111 = (1'h0);
  reg [(5'h11):(1'h0)] reg1110 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1109 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1108 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1107 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1106 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1105 = (1'h0);
  reg [(4'he):(1'h0)] reg1104 = (1'h0);
  reg [(5'h11):(1'h0)] reg1103 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1102 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1101 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1100 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1099 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1098 = (1'h0);
  reg [(5'h12):(1'h0)] reg1097 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1096 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1095 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1094 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1093 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1092 = (1'h0);
  reg [(5'h18):(1'h0)] reg1091 = (1'h0);
  reg [(5'h17):(1'h0)] reg1090 = (1'h0);
  reg [(4'hf):(1'h0)] reg1089 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1088 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1087 = (1'h0);
  reg [(3'h6):(1'h0)] reg1086 = (1'h0);
  reg [(4'hd):(1'h0)] reg1085 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1084 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1083 = (1'h0);
  reg [(5'h18):(1'h0)] reg1082 = (1'h0);
  reg [(4'hd):(1'h0)] reg1081 = (1'h0);
  wire [(4'ha):(1'h0)] wire1080;
  reg [(2'h3):(1'h0)] reg1079 = (1'h0);
  reg [(2'h2):(1'h0)] reg1078 = (1'h0);
  reg [(3'h6):(1'h0)] reg1077 = (1'h0);
  reg [(5'h15):(1'h0)] reg1076 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1075 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1074 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1073 = (1'h0);
  reg [(4'h8):(1'h0)] reg1072 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1071 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1070 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1069 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1068 = (1'h0);
  wire [(4'hc):(1'h0)] wire1067;
  reg [(2'h3):(1'h0)] reg1066 = (1'h0);
  reg [(5'h13):(1'h0)] reg1065 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1064 = (1'h0);
  reg [(5'h11):(1'h0)] reg1063 = (1'h0);
  reg [(5'h14):(1'h0)] reg1062 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1061 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1060 = (1'h0);
  reg [(2'h2):(1'h0)] reg1059 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1058 = (1'h0);
  reg [(3'h6):(1'h0)] reg1057 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1056 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1055 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1054 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1053 = (1'h0);
  reg [(5'h16):(1'h0)] reg1052 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1051 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1050 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1049 = (1'h0);
  reg [(3'h7):(1'h0)] reg1048 = (1'h0);
  reg [(4'ha):(1'h0)] reg1047 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1046 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1045 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1044 = (1'h0);
  reg [(5'h16):(1'h0)] reg1043 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1042 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1038 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1041 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1040 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1039 = (1'h0);
  reg [(5'h18):(1'h0)] reg1038 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1037 = (1'h0);
  reg [(4'h8):(1'h0)] reg1036 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1035 = (1'h0);
  reg [(5'h15):(1'h0)] reg1034 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1033 = (1'h0);
  reg [(4'hf):(1'h0)] reg1032 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1031 = (1'h0);
  reg [(3'h7):(1'h0)] reg1030 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1029 = (1'h0);
  reg [(4'he):(1'h0)] reg1028 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1027 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1026 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1025 = (1'h0);
  reg [(5'h11):(1'h0)] reg1024 = (1'h0);
  wire [(5'h13):(1'h0)] wire1023;
  wire [(5'h17):(1'h0)] wire1022;
  reg [(5'h15):(1'h0)] reg1021 = (1'h0);
  reg [(5'h11):(1'h0)] reg1020 = (1'h0);
  reg [(3'h6):(1'h0)] reg1019 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1018 = (1'h0);
  reg [(5'h18):(1'h0)] reg1017 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1016 = (1'h0);
  reg [(4'hc):(1'h0)] reg1015 = (1'h0);
  reg [(5'h11):(1'h0)] reg1014 = (1'h0);
  reg [(4'he):(1'h0)] reg1013 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1012 = (1'h0);
  reg [(4'he):(1'h0)] reg1011 = (1'h0);
  reg [(5'h14):(1'h0)] reg1010 = (1'h0);
  wire [(4'h9):(1'h0)] wire1009;
  reg signed [(4'hf):(1'h0)] reg1008 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1007 = (1'h0);
  reg [(5'h14):(1'h0)] reg1006 = (1'h0);
  reg [(4'hf):(1'h0)] reg1005 = (1'h0);
  reg [(4'hc):(1'h0)] reg1004 = (1'h0);
  reg [(4'hd):(1'h0)] reg1003 = (1'h0);
  reg [(5'h16):(1'h0)] reg1002 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1001 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1000 = (1'h0);
  reg [(5'h16):(1'h0)] reg999 = (1'h0);
  reg [(3'h4):(1'h0)] reg998 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg997 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar996 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg995 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar994 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg993 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg992 = (1'h0);
  reg [(5'h16):(1'h0)] reg991 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg990 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg989 = (1'h0);
  reg [(3'h7):(1'h0)] reg988 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg987 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg986 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar985 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg984 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg983 = (1'h0);
  reg [(4'hd):(1'h0)] reg982 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg981 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg980 = (1'h0);
  reg [(4'h9):(1'h0)] reg979 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg978 = (1'h0);
  reg [(4'hd):(1'h0)] forvar977 = (1'h0);
  reg signed [(4'he):(1'h0)] reg976 = (1'h0);
  reg [(5'h14):(1'h0)] forvar975 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg974 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg973 = (1'h0);
  reg signed [(4'he):(1'h0)] reg972 = (1'h0);
  reg [(3'h4):(1'h0)] forvar971 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar970 = (1'h0);
  reg [(3'h4):(1'h0)] reg969 = (1'h0);
  reg [(5'h1a):(1'h0)] reg968 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg967 = (1'h0);
  reg [(4'hf):(1'h0)] reg966 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg965 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg964 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire963;
  assign y = {reg1141,
                 reg1140,
                 reg1139,
                 reg1138,
                 reg1137,
                 reg1136,
                 wire1135,
                 reg1134,
                 reg1133,
                 reg1132,
                 reg1131,
                 wire1130,
                 wire1129,
                 wire1128,
                 reg1127,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1123,
                 reg1122,
                 forvar1121,
                 reg1120,
                 reg1119,
                 forvar1118,
                 reg1117,
                 reg1116,
                 reg1115,
                 reg1114,
                 reg1113,
                 reg1112,
                 reg1111,
                 reg1110,
                 reg1109,
                 reg1108,
                 forvar1107,
                 reg1106,
                 reg1105,
                 reg1104,
                 reg1103,
                 forvar1102,
                 forvar1101,
                 reg1100,
                 reg1099,
                 reg1098,
                 reg1097,
                 reg1096,
                 reg1095,
                 forvar1094,
                 forvar1093,
                 reg1092,
                 reg1091,
                 reg1090,
                 reg1089,
                 forvar1088,
                 forvar1087,
                 reg1086,
                 reg1085,
                 reg1084,
                 reg1083,
                 reg1082,
                 reg1081,
                 wire1080,
                 reg1079,
                 reg1078,
                 reg1077,
                 reg1076,
                 reg1075,
                 reg1074,
                 reg1073,
                 reg1072,
                 reg1071,
                 forvar1070,
                 reg1069,
                 reg1068,
                 wire1067,
                 reg1066,
                 reg1065,
                 forvar1064,
                 reg1063,
                 reg1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 forvar1058,
                 reg1057,
                 reg1056,
                 reg1055,
                 forvar1054,
                 reg1053,
                 reg1052,
                 reg1051,
                 reg1050,
                 reg1049,
                 reg1048,
                 reg1047,
                 forvar1046,
                 reg1045,
                 reg1044,
                 reg1043,
                 reg1042,
                 forvar1038,
                 reg1041,
                 forvar1040,
                 reg1039,
                 reg1038,
                 reg1037,
                 reg1036,
                 forvar1035,
                 reg1034,
                 forvar1033,
                 reg1032,
                 reg1031,
                 reg1030,
                 reg1029,
                 reg1028,
                 forvar1027,
                 forvar1026,
                 reg1025,
                 reg1024,
                 wire1023,
                 wire1022,
                 reg1021,
                 reg1020,
                 reg1019,
                 reg1018,
                 reg1017,
                 reg1016,
                 reg1015,
                 reg1014,
                 reg1013,
                 forvar1012,
                 reg1011,
                 reg1010,
                 wire1009,
                 reg1008,
                 forvar1007,
                 reg1006,
                 reg1005,
                 reg1004,
                 reg1003,
                 reg1002,
                 reg1001,
                 forvar1000,
                 reg999,
                 reg998,
                 reg997,
                 forvar996,
                 reg995,
                 forvar994,
                 reg993,
                 reg992,
                 reg991,
                 reg990,
                 reg989,
                 reg988,
                 reg987,
                 reg986,
                 forvar985,
                 reg984,
                 reg983,
                 reg982,
                 reg981,
                 reg980,
                 reg979,
                 reg978,
                 forvar977,
                 reg976,
                 forvar975,
                 reg974,
                 reg973,
                 reg972,
                 forvar971,
                 forvar970,
                 reg969,
                 reg968,
                 reg967,
                 reg966,
                 reg965,
                 reg964,
                 wire963,
                 (1'h0)};
  assign wire963 = "X6mr7aqQF";
  always
    @(posedge clk) begin
      reg964 <= $unsigned("65MePCZPW1AdnaqpU9oKbCXYd");
      reg965 <= wire960[(5'h11):(2'h3)];
      reg966 = wire961[(4'hc):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg967 = wire958[(2'h3):(2'h2)];
      reg968 = wire963;
      reg969 = reg965;
      for (forvar970 = (1'h0); (forvar970 < (1'h0)); forvar970 = (forvar970 + (1'h1)))
        begin
          for (forvar971 = (1'h0); (forvar971 < (1'h1)); forvar971 = (forvar971 + (1'h1)))
            begin
              reg972 <= wire960;
              reg973 <= (~|reg966[(4'h8):(1'h1)]);
              reg974 = reg964;
              for (forvar975 = (1'h0); (forvar975 < (2'h3)); forvar975 = (forvar975 + (1'h1)))
                begin
                  reg976 <= forvar975[(2'h3):(2'h2)];
                end
              for (forvar977 = (1'h0); (forvar977 < (2'h3)); forvar977 = (forvar977 + (1'h1)))
                begin
                  reg978 = "DkuDtAYf41Vve";
                  reg979 = $signed((8'ha2));
                  reg980 <= $unsigned($unsigned(forvar971));
                  reg981 <= reg979[(3'h4):(3'h4)];
                  reg982 = ((wire961[(1'h0):(1'h0)] >> {{(reg968 ?
                                  (8'h9e) : wire958)}}) ?
                      {"",
                          ({$unsigned((8'hb7)),
                              $signed((7'h4d))} * {$signed(reg974),
                              "SHnrJPmm4RZMVzZqAA"})} : {{$unsigned(wire958)}});
                  reg983 = ("EuCMDMbhZm" <= $unsigned("1HgHxZ"));
                end
            end
          reg984 <= (($signed(reg980[(1'h0):(1'h0)]) ?
              reg969 : (~&(^$unsigned(wire962)))) * (reg966[(4'h9):(3'h4)] >>> reg983[(1'h0):(1'h0)]));
          for (forvar985 = (1'h0); (forvar985 < (1'h0)); forvar985 = (forvar985 + (1'h1)))
            begin
              reg986 <= (&$unsigned(reg966[(3'h6):(2'h2)]));
              reg987 <= (~forvar977);
              reg988 <= $signed({forvar977[(4'hb):(2'h3)], "8cL4pzzq"});
            end
          reg989 <= (("2G7RAKw4mh0vBIGa6o63fyAS" != $signed({$unsigned(reg969)})) | "FBt2UJ0XygEbiBmrwL6N");
          reg990 <= {(~&(($signed(reg973) <<< $signed(reg986)) + ($unsigned(reg988) * $unsigned(reg979)))),
              (reg989[(1'h0):(1'h0)] ?
                  $unsigned((8'hb4)) : {{"YJfbgBJ13avPaspG3d"}})};
          reg991 <= (($unsigned($unsigned($unsigned(wire963))) ?
                  (($signed(forvar971) || reg976[(3'h5):(2'h3)]) ?
                      ({wire960, reg976} >> (reg987 ?
                          (8'ha5) : (8'hb3))) : $unsigned($unsigned(forvar971))) : "qmO") ?
              (|reg981) : (!"cND"));
        end
    end
  always
    @(posedge clk) begin
      reg992 = $signed(wire959[(1'h0):(1'h0)]);
      reg993 <= ($unsigned($unsigned((+"LRD2WpmyxfW8s40h"))) ?
          (reg968 && (reg976 ?
              reg980[(3'h5):(1'h1)] : (!(reg979 ?
                  forvar970 : reg990)))) : $signed(((-reg992[(5'h19):(5'h18)]) ?
              reg982 : (wire960 || reg973))));
      for (forvar994 = (1'h0); (forvar994 < (3'h4)); forvar994 = (forvar994 + (1'h1)))
        begin
          reg995 <= {"Ng8axqgApOk7c3vv", reg965};
          for (forvar996 = (1'h0); (forvar996 < (1'h1)); forvar996 = (forvar996 + (1'h1)))
            begin
              reg997 = {("SJPTU" ^~ "cxpISbwJyKFiSSlhE"), "U45uJdL3l7a"};
              reg998 <= $signed("qhIk5m");
              reg999 <= (((wire963[(2'h2):(1'h0)] ~^ ($unsigned(reg964) ?
                      (forvar975 ? wire958 : reg989) : (!wire963))) ?
                  {reg974,
                      reg974[(2'h2):(1'h0)]} : {(~|(forvar994 | reg997))}) >= reg978);
              for (forvar1000 = (1'h0); (forvar1000 < (2'h2)); forvar1000 = (forvar1000 + (1'h1)))
                begin
                  reg1001 <= reg983[(3'h4):(1'h1)];
                  reg1002 <= $unsigned(((7'h4d) | (|"esA")));
                end
              reg1003 <= (reg993 == "KFzwuhsoAWRb88DRpwRD");
              reg1004 <= {"7urucCba1neb1AQkL",
                  $signed(("JJZzR4SDRCp" ? ((-reg979) ^ reg966) : wire961))};
            end
        end
      reg1005 <= (reg992[(4'ha):(3'h5)] << (^("YuiteVpe" ?
          $unsigned($signed(reg995)) : (8'h9c))));
      reg1006 <= $unsigned((+("LDGHvPGRQdOD5tbbzdoB" ?
          reg992[(5'h17):(4'hc)] : "K6tBBcK66M0poPacLAKI")));
      for (forvar1007 = (1'h0); (forvar1007 < (1'h0)); forvar1007 = (forvar1007 + (1'h1)))
        begin
          reg1008 <= (8'h9d);
        end
    end
  assign wire1009 = (&reg998);
  always
    @(posedge clk) begin
      reg1010 <= $signed(reg997);
      reg1011 <= reg1005;
      for (forvar1012 = (1'h0); (forvar1012 < (2'h3)); forvar1012 = (forvar1012 + (1'h1)))
        begin
          reg1013 <= (wire959 ^~ {{(forvar996[(4'hf):(3'h6)] || reg964[(4'h8):(4'h8)]),
                  reg983[(3'h7):(2'h2)]},
              ((-"H1TfF71T") ? {reg986} : forvar1012[(3'h4):(2'h2)])});
          reg1014 <= (+reg1010[(4'h8):(1'h1)]);
          reg1015 <= reg978[(4'h8):(3'h5)];
          reg1016 <= ((!$signed("17DfFPFtZGVQt0")) ? "8FtyLZ0tbhq8I" : reg974);
        end
      reg1017 <= (8'hb7);
    end
  always
    @(posedge clk) begin
      reg1018 <= reg1017[(4'h8):(3'h5)];
    end
  always
    @(posedge clk) begin
      reg1019 <= (!(forvar971 ?
          $unsigned(wire961) : "xSUAOB8rHTWUbDBlopNNGhT"));
      reg1020 <= forvar996[(2'h3):(1'h0)];
      reg1021 <= {"",
          ($unsigned(reg988[(3'h5):(1'h0)]) > reg1006[(4'hf):(4'h8)])};
    end
  assign wire1022 = (reg965[(1'h1):(1'h1)] ^ (reg972 <= (wire958 ?
                        {reg969, wire960} : ("R0JHABzQM0urrp" ?
                            (reg1014 - reg1006) : "aUu5P0hr57ph6lQLY2C"))));
  assign wire1023 = ($signed((reg1020[(5'h11):(4'hf)] ?
                            reg997[(1'h1):(1'h1)] : wire960[(4'ha):(3'h6)])) ?
                        (+$signed((((7'h46) & forvar1012) << reg964))) : $unsigned((reg1001[(5'h11):(5'h10)] ?
                            $unsigned($signed(reg978)) : reg1002[(5'h10):(3'h4)])));
  always
    @(posedge clk) begin
      reg1024 <= $unsigned({($signed(wire963) ?
              reg979 : $unsigned((+reg1013)))});
      reg1025 = reg1005;
      for (forvar1026 = (1'h0); (forvar1026 < (1'h0)); forvar1026 = (forvar1026 + (1'h1)))
        begin
          for (forvar1027 = (1'h0); (forvar1027 < (1'h0)); forvar1027 = (forvar1027 + (1'h1)))
            begin
              reg1028 <= $unsigned($unsigned((|"plFxD10phKBR")));
              reg1029 <= reg1016;
              reg1030 <= $unsigned(reg967);
              reg1031 <= reg1019;
              reg1032 <= $unsigned(reg986);
            end
        end
      for (forvar1033 = (1'h0); (forvar1033 < (1'h1)); forvar1033 = (forvar1033 + (1'h1)))
        begin
          reg1034 <= (("XL" && "AnxOB7cAPZY") > {(($unsigned((8'hac)) ?
                      $unsigned(wire963) : (|wire1022)) ?
                  $signed("KFLcKfaQsblJxJngE") : ({wire960, reg991} ?
                      forvar1007[(3'h6):(3'h6)] : $signed(wire1022)))});
        end
      for (forvar1035 = (1'h0); (forvar1035 < (1'h1)); forvar1035 = (forvar1035 + (1'h1)))
        begin
          reg1036 <= "";
        end
    end
  always
    @(posedge clk) begin
      reg1037 <= forvar1033;
      if ((forvar996 ?
          $signed((reg1037 ?
              (reg1013 | (forvar994 + reg999)) : $unsigned((forvar1027 ?
                  reg1037 : reg980)))) : (8'ha7)))
        begin
          reg1038 <= wire961;
          reg1039 <= forvar985[(1'h1):(1'h0)];
          for (forvar1040 = (1'h0); (forvar1040 < (2'h3)); forvar1040 = (forvar1040 + (1'h1)))
            begin
              reg1041 = (~^forvar1012);
            end
        end
      else
        begin
          for (forvar1038 = (1'h0); (forvar1038 < (2'h2)); forvar1038 = (forvar1038 + (1'h1)))
            begin
              reg1039 <= $unsigned(reg980);
              for (forvar1040 = (1'h0); (forvar1040 < (3'h4)); forvar1040 = (forvar1040 + (1'h1)))
                begin
                  reg1041 <= wire960[(4'hc):(4'ha)];
                  reg1042 <= $signed((~|((8'h9f) ?
                      ((!reg1001) ?
                          reg1008[(4'ha):(4'h8)] : $signed(reg980)) : $unsigned($unsigned(reg1006)))));
                  reg1043 <= (-(|$unsigned($unsigned($unsigned(reg1003)))));
                  reg1044 <= "";
                  reg1045 = (+((|$signed(reg1038)) ?
                      (reg1015 ?
                          $unsigned("ytsYN") : reg1036[(3'h7):(3'h7)]) : reg1013));
                end
              for (forvar1046 = (1'h0); (forvar1046 < (1'h0)); forvar1046 = (forvar1046 + (1'h1)))
                begin
                  reg1047 = $signed(($unsigned($signed((reg1015 <= reg1010))) < ("zOBOH" ~^ forvar1046[(4'he):(3'h6)])));
                end
              reg1048 <= reg984[(5'h13):(4'hb)];
              reg1049 = $unsigned("DksYqDx");
              reg1050 = $unsigned("lQMKMBEQCbtcT");
            end
          reg1051 <= (reg1020 <<< reg1024);
          reg1052 <= $unsigned($unsigned({(^((8'hb0) ?
                  forvar1027 : forvar1027))}));
          reg1053 <= "BgROE7";
          for (forvar1054 = (1'h0); (forvar1054 < (1'h0)); forvar1054 = (forvar1054 + (1'h1)))
            begin
              reg1055 <= (~|$signed("yNAxGpQLo83"));
              reg1056 <= $unsigned("4CxfqaCtyGNLT67FOq3");
            end
          reg1057 <= $unsigned((reg989 ~^ "5KQnuW"));
        end
    end
  always
    @(posedge clk) begin
      for (forvar1058 = (1'h0); (forvar1058 < (1'h1)); forvar1058 = (forvar1058 + (1'h1)))
        begin
          reg1059 <= $unsigned((&reg982[(2'h3):(2'h2)]));
          reg1060 <= (({"0ripm8ErOvsJ8TouK"} & (+($unsigned(reg1045) >>> {(8'hb9)}))) - "akK4P328u8rlr4cJ");
          reg1061 = {(reg1011[(3'h5):(3'h4)] >> reg976),
              ((~^reg1051) ?
                  $unsigned($signed(reg1028[(4'he):(1'h0)])) : $unsigned((-reg991)))};
          reg1062 = "CyH9XIX1VgU";
          reg1063 = (reg995[(3'h5):(2'h3)] | (&reg997[(4'h9):(4'h8)]));
        end
      for (forvar1064 = (1'h0); (forvar1064 < (1'h0)); forvar1064 = (forvar1064 + (1'h1)))
        begin
          reg1065 <= "o99IqHRT76Fyifk7";
        end
      reg1066 <= (^~$signed((("XtoevAb" ? (~&reg972) : (reg968 || forvar970)) ?
          ("sLizm8fNKU" < "Y4TiBqT") : $signed($signed(reg1061)))));
    end
  assign wire1067 = $signed((forvar1054 ? reg1057[(1'h0):(1'h0)] : (~&reg972)));
  always
    @(posedge clk) begin
      reg1068 = ($signed(("X77gGk5ulyxZ3" ?
          reg1003[(4'hb):(4'ha)] : "4dp42019B5m9MbnHeZWBsnFGU")) == wire1067);
      reg1069 <= reg1056;
      for (forvar1070 = (1'h0); (forvar1070 < (3'h5)); forvar1070 = (forvar1070 + (1'h1)))
        begin
          reg1071 <= (!reg1013[(4'hb):(1'h1)]);
          reg1072 <= "GeAyqbpREC45We8";
          reg1073 <= (~"CzRSceG7k5xZvCSodHQdMuh7p");
          reg1074 = ("yyZKqxIEByB9LLT6P" & $unsigned(forvar1012));
          reg1075 <= $signed($signed((^(-"kmxJnSTmQ7UP536Lh"))));
          reg1076 <= $unsigned($signed((~|$signed("AUSdo6WcHt9fh7I95kCdC12X"))));
        end
      reg1077 = "ya6O6";
      reg1078 = (-((^$signed($signed(reg1008))) <<< forvar1064[(2'h2):(1'h0)]));
      reg1079 <= $unsigned($unsigned("JbChwFlmAwaHrbqbs"));
    end
  assign wire1080 = (wire963[(2'h2):(2'h2)] ?
                        "2qBm5qVc9a9uy" : $unsigned($signed(reg1016[(3'h6):(2'h3)])));
  always
    @(posedge clk) begin
      reg1081 = reg1076[(3'h5):(2'h2)];
      reg1082 <= (((|reg1029[(3'h5):(3'h4)]) ?
          ($signed((&reg1042)) != (!$signed(reg1030))) : forvar1033) <= $signed("Z"));
      reg1083 <= reg990;
      reg1084 <= (-$unsigned($signed(reg1020[(4'h8):(2'h3)])));
    end
  always
    @(posedge clk) begin
      reg1085 = reg973[(2'h2):(1'h0)];
      reg1086 <= forvar1033[(3'h5):(2'h2)];
      for (forvar1087 = (1'h0); (forvar1087 < (3'h5)); forvar1087 = (forvar1087 + (1'h1)))
        begin
          for (forvar1088 = (1'h0); (forvar1088 < (3'h5)); forvar1088 = (forvar1088 + (1'h1)))
            begin
              reg1089 <= "2Tx8A8CgMblRvJ0k";
              reg1090 <= $signed(forvar1007);
            end
          reg1091 <= reg1017[(4'he):(4'ha)];
          reg1092 <= $signed({$unsigned((~&(~&reg1090))),
              $signed($unsigned(((8'hb0) ? reg969 : reg1044)))});
        end
    end
  always
    @(posedge clk) begin
      for (forvar1093 = (1'h0); (forvar1093 < (1'h1)); forvar1093 = (forvar1093 + (1'h1)))
        begin
          for (forvar1094 = (1'h0); (forvar1094 < (1'h1)); forvar1094 = (forvar1094 + (1'h1)))
            begin
              reg1095 = $unsigned((forvar985 ?
                  reg990[(3'h7):(2'h3)] : $unsigned(((reg978 ?
                          reg1015 : wire1009) ?
                      wire1080[(2'h3):(1'h0)] : $unsigned((8'hb3))))));
              reg1096 <= reg1089;
              reg1097 <= reg1081[(4'hd):(1'h0)];
              reg1098 <= reg989[(2'h3):(1'h0)];
              reg1099 = ("Y" ? wire958 : "4g");
              reg1100 <= (!$unsigned(reg1039));
            end
          for (forvar1101 = (1'h0); (forvar1101 < (3'h5)); forvar1101 = (forvar1101 + (1'h1)))
            begin
              for (forvar1102 = (1'h0); (forvar1102 < (3'h4)); forvar1102 = (forvar1102 + (1'h1)))
                begin
                  reg1103 <= ($unsigned(reg1015) && (reg1011[(4'h9):(1'h1)] ?
                      ($signed(reg1019) >>> (~^(+reg1029))) : ("vye6L6BfqYsONkmlmeQvrpX7k" ?
                          (|((8'h9f) ? reg1079 : reg1021)) : (8'hb8))));
                  reg1104 = ({(|{$signed(forvar1046), $signed(forvar1027)}),
                          reg1049} ?
                      reg1083 : {reg1005});
                  reg1105 = ((($signed("Z5Bm7zYdB1Bn") ?
                              reg1045 : ($unsigned(forvar1038) - forvar1038[(1'h0):(1'h0)])) ?
                          (($unsigned(reg968) ?
                              $signed(reg988) : (^reg1090)) | (forvar971 && $unsigned(forvar996))) : $unsigned(((7'h44) ?
                              reg1029 : $signed((7'h46))))) ?
                      (&{forvar975[(4'hc):(3'h4)]}) : $unsigned(($unsigned({reg1010}) <<< wire962)));
                  reg1106 = (reg997 ^ "x32HTKDdEeBkqcaaOKl2Pdd0r");
                end
              for (forvar1107 = (1'h0); (forvar1107 < (2'h2)); forvar1107 = (forvar1107 + (1'h1)))
                begin
                  reg1108 = forvar1094[(1'h1):(1'h1)];
                  reg1109 <= reg1004[(4'ha):(3'h5)];
                end
            end
          reg1110 <= (-$unsigned({$signed(((8'ha5) * reg1006))}));
          reg1111 <= (&(reg1077[(2'h3):(1'h1)] ?
              $signed({(reg1110 ^ wire1009),
                  $signed(reg1076)}) : ((reg1034 < (+(7'h4b))) - "J5MTTL4Z")));
          reg1112 <= $signed($signed(reg1030[(1'h1):(1'h1)]));
          reg1113 = (!reg1038);
        end
      reg1114 <= "q2CyBbQTxkofI";
      reg1115 = $signed((!(!reg1016)));
      reg1116 <= forvar971[(2'h3):(2'h2)];
      reg1117 = (+($signed((-((8'hbe) < reg1008))) == "5GoxSO7CFgMZm0teaCkRLdW7T"));
      for (forvar1118 = (1'h0); (forvar1118 < (2'h3)); forvar1118 = (forvar1118 + (1'h1)))
        begin
          reg1119 <= {(8'hbc), reg1057};
          reg1120 <= reg1079[(2'h2):(1'h1)];
          for (forvar1121 = (1'h0); (forvar1121 < (3'h4)); forvar1121 = (forvar1121 + (1'h1)))
            begin
              reg1122 <= "vafXcu";
              reg1123 <= forvar985;
              reg1124 <= $unsigned(("FyS8NLpEB7tJTmIW4D" ?
                  reg1025 : (^~$unsigned(reg1025))));
              reg1125 = {(({(reg1113 ? forvar1040 : forvar1027),
                          "8bWpRMr9MAOprhZ"} | (8'hba)) ?
                      {reg1052,
                          (forvar1033[(2'h3):(1'h0)] || reg1104)} : "vMci62XmUuQSnvNKSAp2ody")};
            end
          reg1126 <= ($signed(reg1045) & forvar975);
          reg1127 <= {"eYUT2HAP1eRh7GP7E", reg1028};
        end
    end
  assign wire1128 = (|reg1116[(4'h9):(3'h4)]);
  assign wire1129 = $unsigned($unsigned(reg1055));
  assign wire1130 = (~$signed((^reg981[(4'hf):(3'h4)])));
  always
    @(posedge clk) begin
      reg1131 = ((^(~^forvar1094)) ?
          $signed((reg1125 > $signed({reg972}))) : reg1002[(3'h6):(3'h5)]);
      reg1132 = "RhYAyvGVWOMlfNCww";
      reg1133 = $signed($unsigned($unsigned(($unsigned(wire958) ?
          $signed((7'h47)) : (reg991 <<< reg1119)))));
      reg1134 = "NypMkC8MGdG";
    end
  assign wire1135 = {(~&$signed(({(8'haa), reg1111} * (wire1009 != reg1122))))};
  always
    @(posedge clk) begin
      reg1136 <= $unsigned(wire960);
      reg1137 <= {(-("rw3R" && $unsigned($signed(reg1079)))),
          $signed(((reg998 ?
              (reg1044 & forvar996) : reg1042[(1'h0):(1'h0)]) > "g1yPhWM1Dfb5"))};
      reg1138 = (("UWlXv" && ($signed("75") ?
              "9wCcWCUgovVak2a56MfHhAw" : (^~(8'h9c)))) ?
          (reg983[(4'hb):(3'h7)] & wire961) : ("UCCqwxdyMpIS2mqyC" ~^ $signed((+reg1013[(3'h4):(3'h4)]))));
      reg1139 <= (&reg1011[(1'h1):(1'h1)]);
      reg1140 = reg1103;
      reg1141 = "y";
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module881  (y, clk, wire885, wire884, wire883, wire882);
  output wire [(32'h33f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire885;
  input wire signed [(5'h15):(1'h0)] wire884;
  input wire signed [(5'h13):(1'h0)] wire883;
  input wire [(5'h18):(1'h0)] wire882;
  reg signed [(5'h13):(1'h0)] reg941 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg942 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar941 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg940 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg939 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg938 = (1'h0);
  reg [(3'h5):(1'h0)] forvar937 = (1'h0);
  reg [(3'h4):(1'h0)] reg936 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg935 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar934 = (1'h0);
  reg signed [(4'he):(1'h0)] reg933 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg932 = (1'h0);
  reg [(4'h8):(1'h0)] reg931 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg930 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg929 = (1'h0);
  reg [(3'h6):(1'h0)] reg928 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg927 = (1'h0);
  reg [(4'ha):(1'h0)] reg926 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar925 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar924 = (1'h0);
  wire [(5'h15):(1'h0)] wire923;
  reg [(5'h17):(1'h0)] reg922 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg921 = (1'h0);
  reg [(4'hc):(1'h0)] reg920 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg919 = (1'h0);
  reg [(5'h18):(1'h0)] reg918 = (1'h0);
  reg [(5'h14):(1'h0)] reg917 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg916 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar915 = (1'h0);
  reg [(2'h2):(1'h0)] reg914 = (1'h0);
  reg [(5'h17):(1'h0)] reg913 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg912 = (1'h0);
  reg [(3'h7):(1'h0)] reg911 = (1'h0);
  reg [(5'h10):(1'h0)] reg910 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg909 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg908 = (1'h0);
  reg [(2'h3):(1'h0)] forvar907 = (1'h0);
  reg [(4'h8):(1'h0)] forvar906 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg905 = (1'h0);
  reg [(4'ha):(1'h0)] reg904 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg902 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg901 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar899 = (1'h0);
  reg [(4'h9):(1'h0)] reg898 = (1'h0);
  reg [(5'h14):(1'h0)] reg897 = (1'h0);
  reg [(5'h19):(1'h0)] reg896 = (1'h0);
  reg [(3'h5):(1'h0)] reg895 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg894 = (1'h0);
  reg [(5'h1a):(1'h0)] reg893 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg892 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar891 = (1'h0);
  reg [(4'hc):(1'h0)] forvar890 = (1'h0);
  reg [(5'h12):(1'h0)] forvar889 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg888 = (1'h0);
  reg [(2'h2):(1'h0)] reg887 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg886 = (1'h0);
  assign y = {reg941,
                 reg942,
                 forvar941,
                 reg940,
                 reg939,
                 reg938,
                 forvar937,
                 reg936,
                 reg935,
                 forvar934,
                 reg933,
                 reg932,
                 reg931,
                 reg930,
                 reg929,
                 reg928,
                 reg927,
                 reg926,
                 forvar925,
                 forvar924,
                 wire923,
                 reg922,
                 reg921,
                 reg920,
                 reg919,
                 reg918,
                 reg917,
                 reg916,
                 forvar915,
                 reg914,
                 reg913,
                 reg912,
                 reg911,
                 reg910,
                 reg909,
                 reg908,
                 forvar907,
                 forvar906,
                 reg905,
                 reg904,
                 reg903,
                 reg902,
                 reg901,
                 reg900,
                 forvar899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 reg893,
                 reg892,
                 forvar891,
                 forvar890,
                 forvar889,
                 reg888,
                 reg887,
                 reg886,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg886 <= ((8'hbe) ?
          $unsigned(wire885) : $signed((wire885 || ((7'h44) ?
              {wire882, wire885} : $unsigned(wire882)))));
      reg887 <= wire882[(3'h7):(1'h1)];
      reg888 <= {(~^($signed(reg887) ?
              ("qvYMt9guRT573tN" << wire883) : (|$unsigned(reg887))))};
      for (forvar889 = (1'h0); (forvar889 < (3'h5)); forvar889 = (forvar889 + (1'h1)))
        begin
          for (forvar890 = (1'h0); (forvar890 < (2'h2)); forvar890 = (forvar890 + (1'h1)))
            begin
              for (forvar891 = (1'h0); (forvar891 < (2'h2)); forvar891 = (forvar891 + (1'h1)))
                begin
                  reg892 <= reg886;
                  reg893 = ((reg886 ?
                          $signed($signed($signed(wire885))) : reg888) ?
                      ($signed(forvar890[(2'h3):(2'h2)]) ?
                          ($signed((8'haf)) > (wire882[(3'h7):(3'h4)] ?
                              $unsigned(forvar889) : "RBvgn5Gr1Kx71ywTvme9plQ0")) : (-$unsigned("AsoraGrG2nRRO"))) : {forvar891[(3'h6):(3'h5)]});
                end
            end
          reg894 <= (reg887[(1'h1):(1'h0)] ?
              ($signed("ZJ7lMbNyvtC39tVogBBaL1Mxp") > $unsigned((^$unsigned(wire883)))) : $signed("HXrqERsOA7esg8rH"));
          reg895 <= (~&("IKKXU" >= "Apyik"));
        end
      reg896 <= "XouMXVO2zhTmki7wr7edDYQ";
    end
  always
    @(posedge clk) begin
      reg897 <= wire882[(5'h17):(1'h0)];
      reg898 <= reg893;
      for (forvar899 = (1'h0); (forvar899 < (2'h3)); forvar899 = (forvar899 + (1'h1)))
        begin
          reg900 <= (~^"SXJGp2D51LdnUmHV6lNWOg");
          reg901 <= ("lf6F9ak5gZ47d3PDpV0" ?
              reg900[(5'h11):(3'h4)] : (((+(!reg886)) ?
                  $signed((~reg886)) : (reg898[(2'h3):(2'h3)] ?
                      (|wire883) : reg897[(5'h13):(1'h1)])) <<< ((+{wire882,
                      reg896}) ?
                  reg886[(3'h7):(1'h0)] : reg896)));
          reg902 <= "lrW6HbgZu8";
          reg903 <= "EwecGq9sd0";
        end
      reg904 <= ($unsigned((~&((+reg888) ? (+reg901) : (reg898 ^ reg894)))) ?
          $unsigned($unsigned(($signed(reg898) ?
              $unsigned(reg894) : $signed((8'ha6))))) : (8'hb8));
      reg905 <= reg897[(2'h2):(2'h2)];
      for (forvar906 = (1'h0); (forvar906 < (3'h4)); forvar906 = (forvar906 + (1'h1)))
        begin
          for (forvar907 = (1'h0); (forvar907 < (3'h5)); forvar907 = (forvar907 + (1'h1)))
            begin
              reg908 = $signed("Fu7ufAQ7k0");
              reg909 <= forvar890;
              reg910 <= reg892[(1'h1):(1'h1)];
              reg911 <= $unsigned(((($unsigned(reg901) < (reg886 ?
                  reg909 : reg886)) || ($signed(forvar907) + ((8'hbb) ?
                  reg893 : reg904))) >= (8'h9e)));
            end
          reg912 <= forvar889;
          reg913 <= "xmwFsr";
          reg914 <= ("rD2oIf1zrDKDkhQg6m" >> "Qq");
          for (forvar915 = (1'h0); (forvar915 < (2'h3)); forvar915 = (forvar915 + (1'h1)))
            begin
              reg916 = $signed(($signed((forvar889 != (reg913 || wire882))) && reg914));
              reg917 <= $unsigned((|$signed({reg898})));
              reg918 <= reg888[(2'h2):(1'h1)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg919 <= ($signed($signed($signed({reg912,
          wire883}))) & $unsigned({(~&(+reg914))}));
      reg920 = "u3mlVFpbfJE6z8";
      reg921 <= {("mwFsYibVeAo4QAYBfekNfzr4x" != $signed("cXKCEdAu88Ps")),
          $unsigned(($unsigned((reg908 ^ reg910)) ?
              (^~"9ci3ULDvfnpm3ykSglFLRFw") : $signed((~|reg909))))};
      reg922 <= $unsigned(((wire882[(3'h7):(3'h7)] ?
              reg903[(4'h9):(4'h8)] : {$signed(reg887)}) ?
          {(~&"")} : $signed(reg903[(4'hf):(4'ha)])));
    end
  assign wire923 = $unsigned($unsigned(reg912[(4'hc):(4'ha)]));
  always
    @(posedge clk) begin
      for (forvar924 = (1'h0); (forvar924 < (1'h0)); forvar924 = (forvar924 + (1'h1)))
        begin
          for (forvar925 = (1'h0); (forvar925 < (1'h0)); forvar925 = (forvar925 + (1'h1)))
            begin
              reg926 = $signed((^(8'hbd)));
              reg927 <= reg911;
              reg928 = $unsigned(({($signed((8'hb3)) | reg896), reg919} ?
                  {reg927} : $signed(reg911[(2'h3):(2'h3)])));
            end
        end
      reg929 = reg926;
      reg930 = {$signed("KOELzkE3PO47UFF2zZokZtFyp")};
      reg931 = reg900;
      reg932 <= (|(reg894[(4'hb):(4'h8)] ? (7'h49) : (~&reg921)));
      reg933 <= ($unsigned(reg932) ?
          ($signed(reg892[(5'h12):(3'h4)]) ?
              forvar899 : (reg897[(4'hd):(3'h6)] ?
                  ((reg930 <= reg901) ?
                      $unsigned(reg921) : $signed(reg928)) : "5cKKA")) : {"laze2DhNXcsmK03mLutIL"});
    end
  always
    @(posedge clk) begin
      for (forvar934 = (1'h0); (forvar934 < (2'h3)); forvar934 = (forvar934 + (1'h1)))
        begin
          reg935 <= (^~$unsigned((reg921 >> $unsigned(wire883))));
          reg936 = (~|reg921[(2'h3):(2'h3)]);
        end
      for (forvar937 = (1'h0); (forvar937 < (3'h5)); forvar937 = (forvar937 + (1'h1)))
        begin
          reg938 <= (8'hbe);
          if (((reg903 ?
              {((reg918 ? reg914 : wire884) ?
                      (reg901 ? reg887 : reg936) : (~reg922)),
                  (reg935[(1'h0):(1'h0)] ?
                      $signed(reg933) : reg898)} : (reg909 == ({reg932} <<< ((8'hbc) != reg908)))) | (((~&$unsigned((8'hb6))) <= forvar915) || wire884[(2'h3):(1'h0)])))
            begin
              reg939 <= ($unsigned(forvar906[(1'h1):(1'h0)]) ^ (reg893[(3'h4):(1'h1)] != (^~{"4dEdNaxUxsG"})));
              reg940 <= $signed($unsigned($signed($unsigned(wire923))));
              for (forvar941 = (1'h0); (forvar941 < (3'h4)); forvar941 = (forvar941 + (1'h1)))
                begin
                  reg942 <= reg901[(3'h7):(1'h1)];
                end
            end
          else
            begin
              reg939 = $signed($signed(($unsigned("BcfURQBiau71cRhneg05fw") ?
                  (&(reg932 ?
                      reg921 : reg898)) : $signed((reg916 != reg905)))));
              if ("9rBBm")
                begin
                  reg940 = "9JfXQ9F4SN3vM2ZnbzeEgTukD";
                end
              else
                begin
                  reg940 <= $unsigned(((((~|reg936) * $signed(forvar937)) ?
                          $signed({reg922}) : reg913) ?
                      $unsigned((reg904[(2'h3):(1'h0)] <<< reg921)) : forvar906));
                  reg941 = (~$unsigned(reg895[(2'h2):(1'h0)]));
                  reg942 <= ("ReOyNauNe" ^ ((({reg931} >> forvar899) ?
                      ((reg928 ^~ reg922) * $signed(reg914)) : $unsigned($signed(reg887))) + reg917[(4'hc):(4'h8)]));
                end
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module757
#( parameter param867 = {(((!((7'h4e) ? (7'h47) : (8'ha0))) <<< {((8'hbb) ? (7'h40) : (8'hbc)), ((7'h42) ? (7'h49) : (8'hbf))}) - ((&((8'ha7) + (8'hac))) & (~^((8'hbd) ^~ (8'haf))))), (^~(+(((7'h43) >> (7'h4e)) ? ((8'h9e) != (7'h45)) : {(7'h48), (8'ha5)})))} )
(y, clk, wire761, wire760, wire759, wire758);
  output wire [(32'h5e5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire761;
  input wire signed [(5'h17):(1'h0)] wire760;
  input wire [(5'h13):(1'h0)] wire759;
  input wire signed [(4'he):(1'h0)] wire758;
  reg [(5'h13):(1'h0)] reg866 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg865 = (1'h0);
  reg [(5'h16):(1'h0)] reg864 = (1'h0);
  reg [(4'hd):(1'h0)] reg863 = (1'h0);
  reg [(3'h5):(1'h0)] reg862 = (1'h0);
  reg [(3'h5):(1'h0)] reg861 = (1'h0);
  reg [(4'hc):(1'h0)] reg860 = (1'h0);
  reg [(5'h14):(1'h0)] reg859 = (1'h0);
  reg [(2'h2):(1'h0)] forvar858 = (1'h0);
  reg [(5'h13):(1'h0)] reg857 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar856 = (1'h0);
  reg [(4'hd):(1'h0)] reg855 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg854 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg853 = (1'h0);
  reg [(3'h4):(1'h0)] reg852 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg850 = (1'h0);
  reg [(5'h14):(1'h0)] reg849 = (1'h0);
  reg [(5'h14):(1'h0)] reg848 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg847 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar846 = (1'h0);
  reg [(4'hb):(1'h0)] reg845 = (1'h0);
  reg [(5'h10):(1'h0)] forvar844 = (1'h0);
  reg [(4'hc):(1'h0)] forvar843 = (1'h0);
  reg [(5'h18):(1'h0)] reg842 = (1'h0);
  reg [(3'h6):(1'h0)] reg841 = (1'h0);
  reg [(2'h3):(1'h0)] reg840 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar839 = (1'h0);
  reg [(4'h9):(1'h0)] reg838 = (1'h0);
  reg [(3'h6):(1'h0)] reg837 = (1'h0);
  reg [(5'h19):(1'h0)] reg836 = (1'h0);
  reg [(5'h16):(1'h0)] forvar835 = (1'h0);
  reg [(3'h4):(1'h0)] forvar834 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg833 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar832 = (1'h0);
  reg [(4'hb):(1'h0)] reg831 = (1'h0);
  reg [(4'he):(1'h0)] reg830 = (1'h0);
  reg [(5'h19):(1'h0)] reg829 = (1'h0);
  reg [(5'h19):(1'h0)] reg828 = (1'h0);
  reg [(5'h13):(1'h0)] reg827 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg826 = (1'h0);
  reg [(5'h15):(1'h0)] reg825 = (1'h0);
  reg [(4'ha):(1'h0)] reg824 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg823 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg822 = (1'h0);
  reg [(5'h17):(1'h0)] reg821 = (1'h0);
  reg [(4'hb):(1'h0)] reg820 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg819 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg818 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar817 = (1'h0);
  reg [(3'h6):(1'h0)] reg816 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg815 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg814 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg813 = (1'h0);
  reg [(4'hb):(1'h0)] reg812 = (1'h0);
  reg [(4'hb):(1'h0)] reg811 = (1'h0);
  reg [(5'h15):(1'h0)] forvar810 = (1'h0);
  reg [(3'h5):(1'h0)] reg809 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg808 = (1'h0);
  reg [(3'h7):(1'h0)] reg807 = (1'h0);
  reg [(4'he):(1'h0)] reg806 = (1'h0);
  reg [(5'h19):(1'h0)] reg805 = (1'h0);
  wire [(5'h11):(1'h0)] wire804;
  wire signed [(4'ha):(1'h0)] wire803;
  reg signed [(5'h18):(1'h0)] reg802 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg801 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg800 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg799 = (1'h0);
  reg [(5'h17):(1'h0)] forvar798 = (1'h0);
  reg [(5'h13):(1'h0)] reg797 = (1'h0);
  reg signed [(4'he):(1'h0)] reg796 = (1'h0);
  reg [(5'h14):(1'h0)] reg795 = (1'h0);
  reg [(5'h14):(1'h0)] reg794 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg793 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg792 = (1'h0);
  reg [(5'h1a):(1'h0)] reg791 = (1'h0);
  reg [(5'h13):(1'h0)] reg790 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg789 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire788;
  wire signed [(3'h6):(1'h0)] wire787;
  reg [(3'h6):(1'h0)] reg786 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg785 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg784 = (1'h0);
  reg [(4'h8):(1'h0)] reg783 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar782 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar781 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg780 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg779 = (1'h0);
  reg [(3'h4):(1'h0)] reg778 = (1'h0);
  reg [(5'h15):(1'h0)] reg777 = (1'h0);
  reg [(4'h8):(1'h0)] forvar776 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg775 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg774 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar773 = (1'h0);
  reg [(4'hb):(1'h0)] reg772 = (1'h0);
  reg [(2'h3):(1'h0)] reg771 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar770 = (1'h0);
  reg [(4'h9):(1'h0)] reg769 = (1'h0);
  reg [(4'hc):(1'h0)] reg768 = (1'h0);
  reg [(5'h18):(1'h0)] reg767 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg766 = (1'h0);
  reg [(5'h18):(1'h0)] reg765 = (1'h0);
  reg [(2'h2):(1'h0)] reg764 = (1'h0);
  wire [(5'h1a):(1'h0)] wire763;
  reg [(2'h2):(1'h0)] reg762 = (1'h0);
  assign y = {reg866,
                 reg865,
                 reg864,
                 reg863,
                 reg862,
                 reg861,
                 reg860,
                 reg859,
                 forvar858,
                 reg857,
                 forvar856,
                 reg855,
                 reg854,
                 reg853,
                 reg852,
                 reg851,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 forvar846,
                 reg845,
                 forvar844,
                 forvar843,
                 reg842,
                 reg841,
                 reg840,
                 forvar839,
                 reg838,
                 reg837,
                 reg836,
                 forvar835,
                 forvar834,
                 reg833,
                 forvar832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 reg827,
                 reg826,
                 reg825,
                 reg824,
                 reg823,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 reg818,
                 forvar817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 reg812,
                 reg811,
                 forvar810,
                 reg809,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 wire804,
                 wire803,
                 reg802,
                 reg801,
                 reg800,
                 reg799,
                 forvar798,
                 reg797,
                 reg796,
                 reg795,
                 reg794,
                 reg793,
                 reg792,
                 reg791,
                 reg790,
                 reg789,
                 wire788,
                 wire787,
                 reg786,
                 reg785,
                 reg784,
                 reg783,
                 forvar782,
                 forvar781,
                 reg780,
                 reg779,
                 reg778,
                 reg777,
                 forvar776,
                 reg775,
                 reg774,
                 forvar773,
                 reg772,
                 reg771,
                 forvar770,
                 reg769,
                 reg768,
                 reg767,
                 reg766,
                 reg765,
                 reg764,
                 wire763,
                 reg762,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg762 <= $signed(wire761);
    end
  assign wire763 = ($unsigned(((&(wire759 >>> wire759)) ?
                       "w46KH2KSk0wA8yGPAsMJm3" : ($signed(wire759) ?
                           (wire758 ?
                               wire760 : (8'hac)) : wire758))) << $signed($unsigned((-"es21MG2uDVDMOk8rnbm"))));
  always
    @(posedge clk) begin
      reg764 <= (reg762[(1'h0):(1'h0)] <= ((wire759[(4'ha):(2'h3)] ?
          (wire760[(2'h3):(1'h1)] ?
              wire761 : wire761[(4'ha):(1'h0)]) : (&wire758)) >> wire760[(3'h7):(3'h7)]));
      reg765 <= {(($signed((reg762 && (7'h4d))) ?
                  $unsigned(wire758) : {(~|wire759)}) ?
              wire758[(2'h3):(2'h2)] : ($signed((8'hae)) >= "UPve55lN"))};
      reg766 <= wire758;
      reg767 <= (-(^reg764[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg768 = ((wire761 ?
          $unsigned(wire763[(5'h14):(5'h14)]) : (~^reg762)) <<< (|(8'hb9)));
      reg769 <= (~&wire758);
      for (forvar770 = (1'h0); (forvar770 < (2'h2)); forvar770 = (forvar770 + (1'h1)))
        begin
          reg771 <= wire758;
          reg772 = $unsigned(((^$unsigned($signed(reg771))) ?
              {$unsigned(reg766[(4'hb):(1'h0)]),
                  reg768[(4'h8):(3'h6)]} : "VEk42V3O"));
        end
    end
  always
    @(posedge clk) begin
      for (forvar773 = (1'h0); (forvar773 < (1'h0)); forvar773 = (forvar773 + (1'h1)))
        begin
          reg774 = $unsigned($signed({"lRLClQQirbRXSpZJzzok1"}));
          reg775 = "QeiSEr";
          for (forvar776 = (1'h0); (forvar776 < (1'h1)); forvar776 = (forvar776 + (1'h1)))
            begin
              reg777 <= (($unsigned($unsigned({reg774})) ?
                  $unsigned((~&"0UlogsyH2WNoyw")) : $unsigned("")) <<< {reg767,
                  (~^$unsigned(wire759))});
              reg778 <= "HxETSEFabwzw8KnVkSyQ";
              reg779 = {($unsigned({reg768[(4'ha):(3'h7)]}) ?
                      "JqG6VCtWFGuOa5PRswa1W" : ((wire760[(5'h14):(5'h11)] ^ (forvar770 != reg767)) ?
                          (!$unsigned(wire759)) : ((~|(8'ha2)) || $signed(reg765)))),
                  (^~"912LokSKdNJNz20WdLYw0vBA")};
              reg780 = wire761[(4'ha):(4'h8)];
            end
          for (forvar781 = (1'h0); (forvar781 < (3'h5)); forvar781 = (forvar781 + (1'h1)))
            begin
              for (forvar782 = (1'h0); (forvar782 < (1'h1)); forvar782 = (forvar782 + (1'h1)))
                begin
                  reg783 = {(("7eY1TPyyH5snOORkx" ^~ (-$signed(reg768))) > wire759)};
                  reg784 <= ((~$signed((^$unsigned((8'ha5))))) ?
                      "aKZTuUL76O5v3N85YmDgpP" : ((forvar770 ?
                              $unsigned(reg769) : forvar770[(1'h0):(1'h0)]) ?
                          {(8'hb1)} : reg777[(5'h12):(4'h9)]));
                  reg785 <= $unsigned($signed($signed("OadR7AIMy")));
                end
            end
          reg786 <= (^$unsigned(reg768));
        end
    end
  assign wire787 = $signed(wire758[(4'h8):(1'h1)]);
  assign wire788 = (((~^{(reg777 ?
                           (8'hbf) : reg768)}) >= "SH6FK8Rd7ymey") - $unsigned((&{reg785[(1'h1):(1'h0)],
                       reg775[(4'h8):(1'h1)]})));
  always
    @(posedge clk) begin
      reg789 <= "RRCXZ3KTkcxbuhZaAArGOCqcX";
      reg790 <= (+$signed($unsigned((reg772 >> ((8'hba) ? reg774 : reg785)))));
      reg791 <= forvar782;
      if (("ep7XabnnlN" >= forvar781[(3'h7):(3'h5)]))
        begin
          reg792 = reg766[(3'h5):(2'h3)];
          reg793 <= $signed($unsigned(($unsigned(reg780[(2'h3):(2'h3)]) ?
              $signed({reg784, reg784}) : reg768[(4'hb):(4'ha)])));
        end
      else
        begin
          reg792 <= (|(|((forvar781[(4'he):(3'h5)] ?
                  (forvar781 ? reg791 : (8'ha8)) : reg765[(3'h4):(1'h0)]) ?
              (reg789[(3'h4):(2'h3)] ?
                  "mVmqstbLTAHT6nNNSLG" : reg791) : ((reg768 - reg774) ?
                  (forvar781 + reg775) : $signed(reg768)))));
          reg793 <= ($signed(reg772) <<< $signed((($signed(reg762) ?
              $unsigned(reg792) : (~^(7'h46))) != forvar773[(4'h9):(1'h1)])));
          reg794 <= ((((reg790[(5'h10):(3'h6)] >>> reg778[(1'h1):(1'h0)]) ?
              ({reg767} ?
                  $signed(reg786) : (reg789 & reg793)) : reg777) != ("9RimpQET" ?
              "lxFaZhqLnygOz3ncPDeSrUm" : reg774[(3'h7):(3'h5)])) > $signed($signed($unsigned($signed(wire758)))));
          reg795 <= (("GF0QlPPcw2Wtd" >= $unsigned({$signed(forvar773),
              ((8'hb9) << reg769)})) * $signed((+reg785[(3'h5):(3'h5)])));
          reg796 <= (!$unsigned($unsigned(($signed(reg794) && (forvar776 * reg767)))));
          reg797 = ((!(~&wire787)) * $signed(reg779));
        end
      for (forvar798 = (1'h0); (forvar798 < (1'h0)); forvar798 = (forvar798 + (1'h1)))
        begin
          reg799 <= ($signed(reg765[(4'he):(4'hc)]) ? wire761 : reg795);
          reg800 = $signed(reg785[(1'h1):(1'h0)]);
          reg801 <= "Mr71AYY";
          reg802 <= reg796;
        end
    end
  assign wire803 = forvar773[(1'h1):(1'h1)];
  assign wire804 = (|$unsigned((^~$unsigned(forvar776))));
  always
    @(posedge clk) begin
      reg805 = "w5He4V2Xu";
      reg806 <= "IHNn4YFV4T";
      reg807 <= $signed((|({$signed(reg801),
          reg793[(5'h10):(4'h8)]} >> "vha")));
      reg808 <= (^~$unsigned({(((8'hba) ? forvar781 : (7'h4c)) ?
              {reg795} : reg771[(1'h1):(1'h0)])}));
      reg809 <= $unsigned(reg778[(1'h0):(1'h0)]);
      for (forvar810 = (1'h0); (forvar810 < (3'h5)); forvar810 = (forvar810 + (1'h1)))
        begin
          reg811 = $signed(({(!(reg808 | wire759)),
              ({(7'h47)} & wire758)} > (^reg769[(2'h2):(1'h1)])));
          reg812 <= (&{reg768[(4'ha):(3'h6)],
              ("FKQXu8Sc" || ((reg807 < reg800) != (!reg786)))});
          reg813 <= reg772;
        end
    end
  always
    @(posedge clk) begin
      reg814 <= (+$signed((((reg783 & (7'h49)) ?
              forvar798 : ((8'hbc) ? reg777 : reg779)) ?
          {(reg789 ? wire763 : reg775),
              (forvar798 ? reg767 : reg802)} : ($signed(reg777) ?
              $signed(reg792) : $unsigned(reg792)))));
      reg815 <= $signed($signed($signed($unsigned($unsigned(reg783)))));
      reg816 <= $signed("eaPDbKnVxH0aM6D7I7QC");
      for (forvar817 = (1'h0); (forvar817 < (3'h4)); forvar817 = (forvar817 + (1'h1)))
        begin
          reg818 <= (reg766 ?
              $signed($signed((~|$unsigned(reg794)))) : (reg793[(3'h5):(3'h5)] ?
                  (+((|reg790) < "CY1MrJWBu6Bied")) : forvar773[(3'h4):(2'h2)]));
          reg819 <= $unsigned((^{$signed((^reg767))}));
          reg820 <= (reg807 <= (reg795[(3'h4):(3'h4)] ?
              $unsigned(reg772[(4'hb):(3'h5)]) : ""));
          reg821 = (8'hb6);
          reg822 = reg794;
          reg823 = $signed("7kggb9ldX64");
        end
      reg824 <= reg768[(2'h2):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg825 <= {reg820[(3'h5):(3'h5)], (!(-{"ZtQoWuRNKvrOTvcu1NSIpt"}))};
      reg826 <= reg790;
    end
  always
    @(posedge clk) begin
      reg827 <= reg762;
      reg828 <= reg821[(2'h2):(1'h0)];
      reg829 <= $unsigned(forvar810[(3'h5):(3'h5)]);
    end
  always
    @(posedge clk) begin
      reg830 <= (reg813[(3'h7):(3'h5)] >>> $signed($signed(("6WbOt2Q" && "cf"))));
      reg831 = ("h" ?
          (reg762[(1'h0):(1'h0)] ?
              ("LqUMcYV4qXOy" ?
                  $signed({reg799}) : {(^reg821),
                      {forvar798}}) : "6kAJ4M2z8O4DQshl") : (~^$unsigned(reg793)));
      for (forvar832 = (1'h0); (forvar832 < (3'h5)); forvar832 = (forvar832 + (1'h1)))
        begin
          reg833 <= (reg786 ?
              "XvkwoaWH" : $signed(($signed(reg821[(2'h3):(1'h0)]) ?
                  reg791 : reg826[(5'h11):(4'hb)])));
          for (forvar834 = (1'h0); (forvar834 < (1'h0)); forvar834 = (forvar834 + (1'h1)))
            begin
              for (forvar835 = (1'h0); (forvar835 < (1'h1)); forvar835 = (forvar835 + (1'h1)))
                begin
                  reg836 <= reg771[(2'h2):(1'h0)];
                  reg837 <= {"6pLVIWGVeA4dKUeDhSwM",
                      $unsigned(reg824[(3'h7):(3'h4)])};
                  reg838 <= {(!{$signed($signed(forvar773)), (~^(|wire761))})};
                end
              for (forvar839 = (1'h0); (forvar839 < (3'h5)); forvar839 = (forvar839 + (1'h1)))
                begin
                  reg840 <= $signed($signed($unsigned({reg830})));
                end
            end
        end
      reg841 <= (reg826 ?
          ($signed("OcCYpTf32AM06lbnBGM0") | (({reg827, reg783} ?
              "FlbTPUs92zAVVs3" : (reg807 ?
                  reg789 : forvar776)) + $signed(reg768))) : "");
    end
  always
    @(posedge clk) begin
      reg842 <= reg815;
      for (forvar843 = (1'h0); (forvar843 < (3'h5)); forvar843 = (forvar843 + (1'h1)))
        begin
          for (forvar844 = (1'h0); (forvar844 < (1'h1)); forvar844 = (forvar844 + (1'h1)))
            begin
              reg845 <= {($signed($signed((wire804 ?
                      reg837 : reg775))) > "mVz3LEKxN54skghEZk4Tz"),
                  ((8'hb3) ? (7'h4d) : $unsigned((^~(^reg809))))};
              for (forvar846 = (1'h0); (forvar846 < (2'h3)); forvar846 = (forvar846 + (1'h1)))
                begin
                  reg847 <= (-(((~^reg780) ?
                      {$unsigned(wire763),
                          (reg824 ?
                              forvar844 : (8'h9e))} : (7'h4b)) > reg831[(3'h7):(3'h6)]));
                  reg848 <= (reg822[(2'h2):(2'h2)] ?
                      (forvar782[(3'h5):(2'h2)] ?
                          ((~&"EAwPNdnAF0") ?
                              ((forvar839 ?
                                  reg845 : reg801) | $unsigned((8'hbc))) : $unsigned("NzWm51y")) : $unsigned(((~|reg836) <= $signed(reg829)))) : (+(~|((!(7'h4b)) + (reg768 == (8'hb2))))));
                  reg849 <= (reg784 * ((~$unsigned((~^reg789))) ?
                      ((((7'h46) - reg786) > $signed(forvar776)) >>> reg825) : {reg786}));
                  reg850 <= (reg795[(2'h3):(2'h2)] | ($signed(reg830[(1'h1):(1'h1)]) + $signed((&(forvar776 ?
                      reg802 : reg814)))));
                  reg851 <= $signed(($signed($unsigned((-reg807))) - {$unsigned($unsigned(reg838))}));
                end
              reg852 <= (+{$unsigned("gfYvBkZsY6WKceiiLmU5zuw1")});
              reg853 = $unsigned($signed(($unsigned((reg811 ?
                      reg820 : reg762)) ?
                  {$signed(reg845)} : "Q62arwcpC")));
            end
          reg854 <= (-wire758);
        end
      reg855 <= "PFo9";
      for (forvar856 = (1'h0); (forvar856 < (3'h4)); forvar856 = (forvar856 + (1'h1)))
        begin
          reg857 <= (({$unsigned((reg854 ? reg816 : (7'h42))),
                  $unsigned(forvar834)} ^~ ((~|reg850) <= ($signed(reg851) ~^ $unsigned(reg795)))) ?
              $unsigned((8'ha9)) : {$signed($unsigned((~reg764))),
                  reg820[(1'h0):(1'h0)]});
          for (forvar858 = (1'h0); (forvar858 < (1'h1)); forvar858 = (forvar858 + (1'h1)))
            begin
              reg859 <= (reg784 ? reg822 : forvar858[(1'h1):(1'h1)]);
              reg860 <= $unsigned("5vzZ6IUe6eJTZn");
            end
          reg861 <= "3RFRcV8FE1Fwyt";
          reg862 <= "l55iy7SCwWO";
        end
      reg863 <= $signed((~^(((reg825 - reg826) != {reg822}) ?
          $signed((forvar856 ? reg813 : wire763)) : ($signed(reg860) ?
              $signed((8'ha1)) : $unsigned((8'hbc))))));
      reg864 <= reg806;
    end
  always
    @(posedge clk) begin
      reg865 <= forvar843[(3'h4):(2'h3)];
      reg866 <= forvar858;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module690
#( parameter param753 = ({((~((7'h42) || (8'ha9))) ? (^~{(7'h43)}) : (((8'hba) ^ (8'h9d)) ? ((7'h42) ? (7'h4b) : (8'hae)) : ((7'h40) <<< (8'ha4))))} > (~^(+(((8'ha6) - (8'ha2)) ? ((8'ha2) ? (8'hbc) : (8'hb6)) : ((8'hbb) ? (8'hb2) : (8'h9d))))))
, parameter param754 = param753 )
(y, clk, wire694, wire693, wire692, wire691);
  output wire [(32'h343):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h16):(1'h0)] wire694;
  input wire signed [(3'h4):(1'h0)] wire693;
  input wire [(5'h18):(1'h0)] wire692;
  input wire signed [(5'h15):(1'h0)] wire691;
  reg [(2'h2):(1'h0)] reg752 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg751 = (1'h0);
  reg [(4'ha):(1'h0)] reg750 = (1'h0);
  reg [(5'h13):(1'h0)] reg749 = (1'h0);
  reg [(4'hd):(1'h0)] reg748 = (1'h0);
  reg [(4'ha):(1'h0)] reg747 = (1'h0);
  reg [(4'hf):(1'h0)] reg746 = (1'h0);
  reg [(3'h6):(1'h0)] reg745 = (1'h0);
  reg signed [(4'he):(1'h0)] reg744 = (1'h0);
  reg [(3'h5):(1'h0)] reg743 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire742;
  reg signed [(4'he):(1'h0)] reg741 = (1'h0);
  reg [(3'h5):(1'h0)] reg740 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg739 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg738 = (1'h0);
  reg [(4'h8):(1'h0)] forvar737 = (1'h0);
  reg [(5'h17):(1'h0)] reg736 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg735 = (1'h0);
  reg [(5'h14):(1'h0)] reg734 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg733 = (1'h0);
  reg [(5'h1a):(1'h0)] reg732 = (1'h0);
  reg [(5'h17):(1'h0)] forvar731 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg730 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg729 = (1'h0);
  reg [(4'hb):(1'h0)] reg728 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg727 = (1'h0);
  reg [(5'h1a):(1'h0)] reg726 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar725 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg724 = (1'h0);
  reg [(3'h5):(1'h0)] reg723 = (1'h0);
  reg [(5'h1a):(1'h0)] reg722 = (1'h0);
  reg [(3'h7):(1'h0)] reg721 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar720 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg719 = (1'h0);
  reg [(2'h3):(1'h0)] reg718 = (1'h0);
  reg [(5'h10):(1'h0)] forvar717 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire716;
  reg [(4'he):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg714 = (1'h0);
  reg [(5'h14):(1'h0)] reg713 = (1'h0);
  reg [(3'h4):(1'h0)] reg712 = (1'h0);
  reg [(3'h4):(1'h0)] reg711 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg710 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg709 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg708 = (1'h0);
  reg [(4'h9):(1'h0)] reg707 = (1'h0);
  reg [(5'h13):(1'h0)] reg706 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar705 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg704 = (1'h0);
  reg [(5'h15):(1'h0)] reg703 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg702 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg701 = (1'h0);
  reg [(5'h18):(1'h0)] reg700 = (1'h0);
  reg [(5'h18):(1'h0)] forvar699 = (1'h0);
  reg [(2'h3):(1'h0)] reg698 = (1'h0);
  reg [(3'h6):(1'h0)] reg697 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg696 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar695 = (1'h0);
  assign y = {reg752,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 reg747,
                 reg746,
                 reg745,
                 reg744,
                 reg743,
                 wire742,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 forvar737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 reg732,
                 forvar731,
                 reg730,
                 reg729,
                 reg728,
                 reg727,
                 reg726,
                 forvar725,
                 reg724,
                 reg723,
                 reg722,
                 reg721,
                 forvar720,
                 reg719,
                 reg718,
                 forvar717,
                 wire716,
                 reg715,
                 reg714,
                 reg713,
                 reg712,
                 reg711,
                 reg710,
                 reg709,
                 reg708,
                 reg707,
                 reg706,
                 forvar705,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 forvar699,
                 reg698,
                 reg697,
                 reg696,
                 forvar695,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar695 = (1'h0); (forvar695 < (3'h4)); forvar695 = (forvar695 + (1'h1)))
        begin
          reg696 <= wire693[(2'h2):(1'h1)];
          reg697 <= "qt7chkyBEzrKuLxm";
          reg698 <= "MAxT";
          for (forvar699 = (1'h0); (forvar699 < (3'h4)); forvar699 = (forvar699 + (1'h1)))
            begin
              reg700 <= $unsigned((~(^$signed($signed(forvar695)))));
            end
          reg701 <= $signed($signed((($signed((8'hb4)) >= {wire691}) == (~|forvar695[(3'h4):(2'h2)]))));
        end
      reg702 <= $unsigned("cXDEua");
      reg703 <= forvar699[(5'h17):(5'h16)];
      reg704 = ({("a9Y" == $unsigned((wire691 ?
              reg696 : wire692)))} || $signed("9NnE1m1dqX62d81Q78aq"));
      for (forvar705 = (1'h0); (forvar705 < (3'h5)); forvar705 = (forvar705 + (1'h1)))
        begin
          reg706 <= $unsigned(($signed($signed(forvar695)) ?
              $unsigned((reg704[(2'h3):(2'h3)] ?
                  (forvar695 ?
                      forvar695 : reg700) : (reg697 ~^ reg703))) : forvar705));
          reg707 = (8'hbf);
          reg708 = (reg697 < "JFLu6hIYJXAOxUJr");
          reg709 = reg704[(1'h0):(1'h0)];
        end
      reg710 <= "MW";
    end
  always
    @(posedge clk) begin
      reg711 <= $unsigned(wire693[(3'h4):(3'h4)]);
      reg712 = reg703;
      reg713 <= (~$unsigned(($signed((reg711 ?
          reg701 : forvar699)) >>> $signed($unsigned(reg711)))));
      reg714 = wire693[(3'h4):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg715 = "RcR3QotlSn5IcbGRDDYBH";
    end
  assign wire716 = ({forvar705[(4'h9):(3'h6)]} ?
                       "3kONbzwM0x61f15" : "L9s3Xo6ra8L7adt1fyvc");
  always
    @(posedge clk) begin
      for (forvar717 = (1'h0); (forvar717 < (2'h3)); forvar717 = (forvar717 + (1'h1)))
        begin
          reg718 = $unsigned((reg710[(2'h3):(1'h1)] ?
              {(^~$unsigned(reg712)),
                  reg702[(3'h5):(3'h5)]} : $signed(wire716[(3'h7):(3'h7)])));
          reg719 = forvar717[(4'h8):(3'h5)];
          for (forvar720 = (1'h0); (forvar720 < (3'h4)); forvar720 = (forvar720 + (1'h1)))
            begin
              reg721 = $signed(reg719[(4'hf):(4'hb)]);
              reg722 <= $signed((-{{$unsigned(reg706),
                      (wire716 << forvar699)}}));
              reg723 = $unsigned(({{(+reg721)},
                  "HLwS"} && ((~^forvar705) & "AQfQ4umfVhtf")));
              reg724 <= reg701[(1'h1):(1'h0)];
              for (forvar725 = (1'h0); (forvar725 < (1'h0)); forvar725 = (forvar725 + (1'h1)))
                begin
                  reg726 = {"eVufNS6YGaf", reg713};
                  reg727 <= reg702[(1'h1):(1'h1)];
                  reg728 <= forvar717;
                  reg729 <= $unsigned((~^(&((-(8'hb9)) ?
                      (+forvar720) : (reg701 ? forvar695 : (8'hab))))));
                  reg730 = ($signed((~&$signed((!reg697)))) ?
                      $unsigned(reg726) : ({reg729[(2'h2):(1'h0)], reg718} ?
                          ($signed(((8'hba) ? (7'h4c) : reg711)) ?
                              "VFC17dIXU0r9hpd" : {wire694,
                                  $signed(reg707)}) : ($signed($unsigned(reg707)) ?
                              $signed($unsigned(forvar717)) : {reg708[(3'h6):(3'h6)]})));
                end
            end
          for (forvar731 = (1'h0); (forvar731 < (1'h1)); forvar731 = (forvar731 + (1'h1)))
            begin
              reg732 <= $unsigned((|reg726[(4'hb):(2'h3)]));
              reg733 = ({({{(8'hbd)}} ?
                      reg718[(2'h3):(2'h2)] : (((7'h43) ?
                          (8'hb8) : reg708) * $unsigned((8'ha3)))),
                  ((wire694[(3'h4):(3'h4)] ?
                          reg700 : ((7'h4e) ? reg723 : wire693)) ?
                      {"7o204oGM8iabC3kS7lwozINL"} : reg700)} > ((~^(|reg713)) + (7'h44)));
              reg734 <= (~^{wire716[(2'h3):(1'h1)]});
              reg735 <= "JdcBVpKQi025";
              reg736 = reg700[(4'hb):(4'h8)];
              for (forvar737 = (1'h0); (forvar737 < (1'h1)); forvar737 = (forvar737 + (1'h1)))
                begin
                  reg738 = (reg724 ? reg696[(2'h2):(1'h1)] : reg708);
                end
            end
          reg739 <= {{($unsigned(forvar705[(4'h9):(1'h1)]) ?
                      {(forvar725 ?
                              forvar695 : reg729)} : ((reg724 >>> reg721) ?
                          reg702 : reg697))},
              $unsigned({(~&$unsigned(reg722)),
                  (&(forvar717 ? forvar699 : (8'hb5)))})};
          reg740 <= reg714;
        end
      reg741 <= {{(^reg702)}, forvar737[(3'h4):(1'h1)]};
    end
  assign wire742 = ("9V7krv" ?
                       ((!reg721) ?
                           reg701[(4'h8):(2'h2)] : $signed(((-reg734) ?
                               $unsigned(wire693) : (forvar737 ?
                                   wire716 : wire694)))) : reg712[(3'h4):(1'h0)]);
  always
    @(posedge clk) begin
      reg743 = $unsigned((reg719 ?
          $signed($unsigned(reg735)) : (-$unsigned((reg707 ?
              reg726 : forvar705)))));
      reg744 <= $unsigned($signed({$unsigned(reg740)}));
      reg745 = $signed($signed((^~((reg710 & reg726) < (wire716 ?
          reg701 : reg744)))));
      reg746 = ((|(reg728[(2'h3):(2'h3)] ?
              ((reg728 ? forvar717 : (7'h46)) ?
                  reg704[(4'he):(4'ha)] : reg729) : reg734)) ?
          {$unsigned({reg723[(3'h4):(2'h2)]}), "whAWTJYmgxzJA5"} : "koVph");
      reg747 <= {wire694[(4'hf):(4'hf)]};
      reg748 <= ($unsigned(($unsigned((forvar737 ? reg739 : reg704)) ?
              reg728[(3'h4):(1'h0)] : (~|((8'hb8) ? reg707 : reg747)))) ?
          reg723[(2'h3):(1'h1)] : $signed($signed((~&forvar725[(3'h5):(1'h1)]))));
    end
  always
    @(posedge clk) begin
      reg749 <= reg714;
      reg750 <= reg736;
      reg751 <= forvar717;
      reg752 <= $signed(((($signed(reg739) * (reg709 ?
          wire692 : wire691)) && (&(~^wire693))) | (($signed(reg734) && ((8'ha1) ?
          reg749 : reg711)) > $signed((reg730 >> reg744)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2707  (y, clk, wire2712, wire2711, wire2710, wire2709, wire2708);
  output wire [(32'h436):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire2712;
  input wire [(4'he):(1'h0)] wire2711;
  input wire [(5'h19):(1'h0)] wire2710;
  input wire signed [(5'h16):(1'h0)] wire2709;
  input wire [(5'h19):(1'h0)] wire2708;
  reg signed [(5'h19):(1'h0)] reg2793 = (1'h0);
  reg [(3'h7):(1'h0)] reg2792 = (1'h0);
  reg [(5'h12):(1'h0)] forvar2791 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2790 = (1'h0);
  reg [(2'h3):(1'h0)] reg2789 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2788 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar2787 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2786 = (1'h0);
  wire [(5'h12):(1'h0)] wire2785;
  wire signed [(3'h7):(1'h0)] wire2784;
  reg signed [(2'h2):(1'h0)] reg2783 = (1'h0);
  wire [(2'h2):(1'h0)] wire2782;
  reg signed [(5'h11):(1'h0)] reg2781 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2780 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2779 = (1'h0);
  reg [(5'h18):(1'h0)] forvar2778 = (1'h0);
  reg [(5'h14):(1'h0)] reg2777 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2776 = (1'h0);
  reg [(4'ha):(1'h0)] reg2775 = (1'h0);
  reg [(3'h4):(1'h0)] reg2774 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2773 = (1'h0);
  reg [(4'hc):(1'h0)] reg2772 = (1'h0);
  reg [(2'h2):(1'h0)] reg2771 = (1'h0);
  wire [(5'h13):(1'h0)] wire2770;
  reg [(4'hd):(1'h0)] reg2769 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2768 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2767 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2766 = (1'h0);
  reg [(5'h14):(1'h0)] reg2765 = (1'h0);
  reg [(5'h18):(1'h0)] reg2764 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2763 = (1'h0);
  reg [(3'h6):(1'h0)] reg2762 = (1'h0);
  reg [(3'h6):(1'h0)] reg2761 = (1'h0);
  reg [(3'h4):(1'h0)] reg2760 = (1'h0);
  reg [(5'h19):(1'h0)] reg2759 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2758 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2757 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2756 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2755 = (1'h0);
  reg [(3'h6):(1'h0)] reg2754 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2753 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2752 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2751 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2750 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2749 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2748 = (1'h0);
  reg [(4'ha):(1'h0)] reg2747 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire2746;
  wire signed [(5'h15):(1'h0)] wire2745;
  wire [(5'h17):(1'h0)] wire2744;
  wire signed [(4'h8):(1'h0)] wire2743;
  wire [(5'h16):(1'h0)] wire2742;
  wire [(5'h11):(1'h0)] wire2741;
  reg [(4'h8):(1'h0)] reg2740 = (1'h0);
  reg [(3'h5):(1'h0)] reg2739 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2738 = (1'h0);
  reg [(4'h9):(1'h0)] reg2737 = (1'h0);
  reg [(5'h12):(1'h0)] reg2736 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2735 = (1'h0);
  reg [(3'h6):(1'h0)] reg2734 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2733 = (1'h0);
  reg [(4'ha):(1'h0)] reg2732 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2731 = (1'h0);
  wire signed [(4'he):(1'h0)] wire2730;
  reg signed [(5'h11):(1'h0)] reg2729 = (1'h0);
  reg [(5'h18):(1'h0)] reg2728 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2727 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg2726 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2725 = (1'h0);
  reg [(5'h10):(1'h0)] reg2724 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2723 = (1'h0);
  wire [(5'h13):(1'h0)] wire2722;
  reg signed [(5'h1a):(1'h0)] reg2721 = (1'h0);
  reg [(5'h12):(1'h0)] reg2720 = (1'h0);
  reg [(4'hb):(1'h0)] reg2719 = (1'h0);
  reg [(3'h6):(1'h0)] reg2718 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2717 = (1'h0);
  wire [(4'hc):(1'h0)] wire2716;
  wire signed [(5'h19):(1'h0)] wire2715;
  wire [(2'h3):(1'h0)] wire2714;
  wire [(5'h13):(1'h0)] wire2713;
  assign y = {reg2793,
                 reg2792,
                 forvar2791,
                 reg2790,
                 reg2789,
                 reg2788,
                 forvar2787,
                 reg2786,
                 wire2785,
                 wire2784,
                 reg2783,
                 wire2782,
                 reg2781,
                 reg2780,
                 reg2779,
                 forvar2778,
                 reg2777,
                 forvar2776,
                 reg2775,
                 reg2774,
                 forvar2773,
                 reg2772,
                 reg2771,
                 wire2770,
                 reg2769,
                 reg2768,
                 reg2767,
                 reg2766,
                 reg2765,
                 reg2764,
                 reg2763,
                 reg2762,
                 reg2761,
                 reg2760,
                 reg2759,
                 reg2758,
                 forvar2757,
                 reg2756,
                 forvar2755,
                 reg2754,
                 reg2753,
                 reg2752,
                 reg2751,
                 reg2750,
                 reg2749,
                 reg2748,
                 reg2747,
                 wire2746,
                 wire2745,
                 wire2744,
                 wire2743,
                 wire2742,
                 wire2741,
                 reg2740,
                 reg2739,
                 reg2738,
                 reg2737,
                 reg2736,
                 forvar2735,
                 reg2734,
                 reg2733,
                 reg2732,
                 forvar2731,
                 wire2730,
                 reg2729,
                 reg2728,
                 reg2727,
                 reg2726,
                 reg2725,
                 reg2724,
                 forvar2723,
                 wire2722,
                 reg2721,
                 reg2720,
                 reg2719,
                 reg2718,
                 reg2717,
                 wire2716,
                 wire2715,
                 wire2714,
                 wire2713,
                 (1'h0)};
  assign wire2713 = (($unsigned($unsigned(wire2711)) ^~ wire2708[(5'h16):(4'hd)]) ?
                        (^{$unsigned("pIuwkCFLDXX31LD8")}) : $signed((8'hae)));
  assign wire2714 = ($signed($unsigned(((~^wire2712) ?
                        wire2713 : (^wire2709)))) ^ $signed(wire2711));
  assign wire2715 = ((wire2711[(4'hc):(4'ha)] ?
                            wire2714 : (((^wire2710) ?
                                $signed(wire2711) : (~^wire2712)) >>> ((wire2714 ?
                                wire2708 : wire2714) > wire2713[(2'h2):(1'h0)]))) ?
                        wire2711 : ($unsigned((wire2708 ?
                                (wire2710 + wire2714) : (7'h4b))) ?
                            $unsigned(wire2710) : ((|"gFvQCEHa8rhuSWeTe1") == ((8'hbc) || (wire2713 ?
                                wire2709 : wire2712)))));
  assign wire2716 = $signed(wire2711[(4'h9):(3'h5)]);
  always
    @(posedge clk) begin
      reg2717 = wire2709;
      reg2718 <= ("EXRRlolr4U00333ZEEAIevpW" >>> "wo5MaMKIk");
      reg2719 = {wire2714[(2'h3):(1'h1)]};
      reg2720 <= reg2718[(2'h2):(1'h0)];
      reg2721 <= wire2708[(5'h13):(5'h12)];
    end
  assign wire2722 = $signed("eycpu3XYFrxtsmJgtAwSSz");
  always
    @(posedge clk) begin
      for (forvar2723 = (1'h0); (forvar2723 < (1'h0)); forvar2723 = (forvar2723 + (1'h1)))
        begin
          reg2724 <= wire2712;
          reg2725 <= ($signed((forvar2723 << $signed(reg2718))) ?
              ((+wire2713) ^~ (($unsigned((8'hb5)) ?
                  $unsigned(reg2721) : "r2OQUmL1P3xFZGa42C") >>> $unsigned("tbseFJ5v0ag"))) : $unsigned(reg2717));
        end
      reg2726 <= $unsigned((!wire2710));
    end
  always
    @(posedge clk) begin
      reg2727 = $unsigned($unsigned("0JNz7VbD0r6"));
      reg2728 = $unsigned(($unsigned(((wire2713 < reg2725) ?
              (wire2713 ? reg2726 : reg2719) : wire2711[(4'hd):(4'hb)])) ?
          $unsigned($signed($signed(reg2727))) : $unsigned($unsigned($signed(wire2711)))));
      reg2729 <= reg2727[(2'h2):(2'h2)];
    end
  assign wire2730 = reg2719[(4'h8):(2'h3)];
  always
    @(posedge clk) begin
      for (forvar2731 = (1'h0); (forvar2731 < (3'h4)); forvar2731 = (forvar2731 + (1'h1)))
        begin
          reg2732 <= (wire2709[(4'he):(4'ha)] & $unsigned($signed(forvar2731)));
        end
      reg2733 <= $unsigned((7'h42));
      reg2734 <= {"PnfL5XJYB4JnsLVwIdm38", reg2727[(1'h0):(1'h0)]};
      for (forvar2735 = (1'h0); (forvar2735 < (2'h3)); forvar2735 = (forvar2735 + (1'h1)))
        begin
          reg2736 <= ((~(wire2711 ?
              $signed(((7'h4c) != reg2717)) : $signed($signed(wire2713)))) <= wire2711[(4'hb):(4'h8)]);
          reg2737 <= wire2710;
          reg2738 = (+(^(wire2714[(1'h0):(1'h0)] ?
              "Fw" : ($unsigned((8'hbc)) ?
                  (forvar2723 ? (8'hb2) : forvar2731) : $signed(wire2709)))));
        end
      reg2739 <= {(((reg2737 ? wire2709 : (wire2709 << reg2728)) << {(wire2730 ?
                      wire2709 : reg2737)}) ?
              {({reg2732, reg2734} ?
                      $signed(wire2722) : $unsigned(reg2733))} : wire2708)};
      reg2740 <= $signed((wire2712 ~^ (~^$signed((reg2724 ?
          wire2715 : reg2736)))));
    end
  assign wire2741 = $signed(reg2724[(4'ha):(4'h9)]);
  assign wire2742 = (reg2724 ? wire2716[(3'h5):(3'h5)] : forvar2735);
  assign wire2743 = $unsigned(wire2711[(4'hd):(1'h1)]);
  assign wire2744 = ("pCfzpTDL3V2O5" == wire2711);
  assign wire2745 = reg2738;
  assign wire2746 = {(($unsigned("VLzFXgelGXCEHK7EyfkBsKcrn") ?
                            ({reg2720,
                                (8'had)} <= reg2738[(1'h1):(1'h0)]) : {{reg2717,
                                    forvar2723},
                                reg2733[(4'hb):(4'ha)]}) > $signed({(wire2708 ?
                                (7'h48) : reg2720),
                            {reg2727}})),
                        $signed($signed("nyix2UfV7XFlVd"))};
  always
    @(posedge clk) begin
      reg2747 <= (~$signed(($unsigned("WXpa6myGtB0Ru") - ($signed(wire2730) ?
          $unsigned(reg2734) : (reg2726 >> reg2738)))));
      reg2748 <= wire2709;
      reg2749 <= reg2729;
      reg2750 <= forvar2731[(3'h5):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg2751 <= $unsigned((^reg2729[(3'h6):(2'h3)]));
      reg2752 = $signed($signed($unsigned(wire2708[(5'h12):(4'hd)])));
      reg2753 <= (~$signed($unsigned({$signed(reg2729)})));
      reg2754 <= ((reg2748 == $signed((wire2722 ?
          "8a7Pdl7CyJEB" : $signed(wire2716)))) | (((8'ha2) * (~^$unsigned(wire2716))) >> $unsigned({$signed(wire2715),
          (reg2728 > wire2715)})));
      for (forvar2755 = (1'h0); (forvar2755 < (2'h2)); forvar2755 = (forvar2755 + (1'h1)))
        begin
          reg2756 <= $signed("End67QbAKdX4qSL4t");
          for (forvar2757 = (1'h0); (forvar2757 < (1'h0)); forvar2757 = (forvar2757 + (1'h1)))
            begin
              reg2758 <= $unsigned(((wire2713[(4'hb):(1'h1)] ?
                      $unsigned("zb2v5YtK") : {wire2730}) ?
                  ($unsigned((wire2730 & (7'h49))) ?
                      wire2716 : "WGp0w") : wire2744));
              reg2759 <= "VpK";
              reg2760 = (+((reg2732[(4'ha):(2'h3)] & reg2737[(4'h8):(3'h7)]) ?
                  ("n8dHT" ?
                      (reg2737[(2'h2):(1'h1)] ~^ (reg2729 ?
                          wire2746 : reg2750)) : "C6kdMPWe7UbUwCfEJxmT68") : reg2756));
              reg2761 <= $unsigned(("MDqfepi5C" << $unsigned({$signed(reg2727),
                  "f"})));
              reg2762 <= ((reg2725 ? $signed(reg2720) : {"49DnJ"}) ?
                  "SgpS0xTOAxBfvSIyH2U" : $unsigned(wire2715));
            end
          reg2763 <= {"CiFDR4He", "DpT"};
        end
      reg2764 = ((~&"6gyWWe9Nf6qDQ2cpG") ? {reg2740[(1'h0):(1'h0)]} : (8'hb8));
    end
  always
    @(posedge clk) begin
      reg2765 <= reg2728;
      reg2766 <= "3USBHyddY0dQf";
    end
  always
    @(posedge clk) begin
      reg2767 <= $unsigned("XboDwZNpOFkmfTRUh");
      reg2768 = $signed(((reg2732[(1'h0):(1'h0)] ?
          reg2747 : $unsigned($unsigned(forvar2731))) >= $signed(reg2763[(2'h3):(2'h3)])));
      reg2769 <= reg2729;
    end
  assign wire2770 = {"Z1BpAd", (^(|"3ZPsJLDKh1ar4ds"))};
  always
    @(posedge clk) begin
      reg2771 <= ({reg2740[(1'h0):(1'h0)], forvar2757} > $unsigned(("Hvy6s" ?
          (reg2720[(4'hf):(3'h6)] | ((7'h41) ?
              reg2724 : (8'ha9))) : ((reg2729 >= wire2708) ?
              (reg2717 <<< forvar2755) : (wire2730 ? (8'h9d) : reg2734)))));
      reg2772 <= "yAX4173SfDr";
      for (forvar2773 = (1'h0); (forvar2773 < (3'h4)); forvar2773 = (forvar2773 + (1'h1)))
        begin
          reg2774 = wire2730[(4'ha):(3'h4)];
          reg2775 <= $unsigned(reg2768[(3'h6):(3'h6)]);
          for (forvar2776 = (1'h0); (forvar2776 < (1'h0)); forvar2776 = (forvar2776 + (1'h1)))
            begin
              reg2777 = (forvar2776 > $signed(reg2758));
            end
        end
      for (forvar2778 = (1'h0); (forvar2778 < (1'h1)); forvar2778 = (forvar2778 + (1'h1)))
        begin
          reg2779 <= reg2733;
          reg2780 = (~$unsigned(((~|reg2769) ?
              (^~$signed((8'hae))) : (((8'h9e) <= reg2750) ?
                  {wire2713, reg2733} : (7'h4b)))));
        end
      reg2781 <= (&(&("5mdlGikCg4FgsrPniqgJKbH9" ?
          $signed(reg2765[(5'h13):(4'ha)]) : (&reg2751[(4'hb):(1'h0)]))));
    end
  assign wire2782 = (reg2736[(4'hd):(3'h6)] ?
                        reg2765 : $unsigned({{((8'hb0) ? reg2768 : wire2741)},
                            reg2780}));
  always
    @(posedge clk) begin
      reg2783 <= (+(wire2745 ?
          reg2758[(4'hd):(4'hd)] : $unsigned((|wire2716))));
    end
  assign wire2784 = (($signed(forvar2776) >= (^~reg2780)) ?
                        "8zRaU49cuJDiPx5BRK36" : {(wire2745 >= "a1I1t6sEluDyu")});
  assign wire2785 = ($signed($unsigned(reg2740[(3'h6):(1'h1)])) + $signed((^~(wire2716[(1'h0):(1'h0)] ?
                        (reg2729 ? reg2719 : (8'hb6)) : $unsigned(reg2718)))));
  always
    @(posedge clk) begin
      reg2786 = reg2779[(4'hb):(1'h1)];
      for (forvar2787 = (1'h0); (forvar2787 < (3'h4)); forvar2787 = (forvar2787 + (1'h1)))
        begin
          reg2788 <= {(reg2728[(3'h7):(3'h5)] < (|("t64fD34Ep5fl1LpBWGGe5" ?
                  $signed(reg2760) : "QX77LUF"))),
              {"iFDspZw20wyUN", reg2759}};
          reg2789 <= (($signed(wire2743[(3'h6):(3'h4)]) ?
                  reg2761 : $signed(reg2780)) ?
              reg2726 : reg2786);
          reg2790 <= "wh1dpZQTqMm595Gabe";
          for (forvar2791 = (1'h0); (forvar2791 < (1'h1)); forvar2791 = (forvar2791 + (1'h1)))
            begin
              reg2792 <= "7fPBXxIAbrcStQCddf";
              reg2793 <= $unsigned($unsigned($unsigned(((&reg2736) ?
                  $signed(forvar2776) : (~&reg2732)))));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2691
#( parameter param2703 = ((8'hb8) ? ((-(~|(^(8'ha2)))) ? {(7'h46), (~&(8'hb3))} : {({(7'h49), (8'haf)} ? ((7'h43) ? (8'ha0) : (8'hab)) : ((8'hb3) >>> (8'hb6)))}) : (8'hb2))
, parameter param2704 = ((-(((param2703 ? param2703 : param2703) ? (~^param2703) : {param2703}) ? ((param2703 ? (8'ha1) : param2703) <<< (param2703 != param2703)) : {(param2703 >> param2703), (-param2703)})) ? (((~|(param2703 ? param2703 : (8'ha4))) ? ((8'hb8) * param2703) : param2703) ? (param2703 && ((-param2703) >> (^param2703))) : (param2703 << (~^(param2703 ? param2703 : (7'h46))))) : {(~(^~(param2703 ? param2703 : param2703)))}) )
(y, clk, wire2696, wire2695, wire2694, wire2693, wire2692);
  output wire [(32'h62):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire2696;
  input wire signed [(4'hf):(1'h0)] wire2695;
  input wire [(4'hd):(1'h0)] wire2694;
  input wire signed [(5'h12):(1'h0)] wire2693;
  input wire [(4'hc):(1'h0)] wire2692;
  reg signed [(5'h14):(1'h0)] reg2702 = (1'h0);
  reg [(3'h4):(1'h0)] reg2701 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2700 = (1'h0);
  wire [(4'h8):(1'h0)] wire2699;
  reg signed [(5'h1a):(1'h0)] reg2698 = (1'h0);
  wire [(5'h17):(1'h0)] wire2697;
  assign y = {reg2702, reg2701, reg2700, wire2699, reg2698, wire2697, (1'h0)};
  assign wire2697 = ("NoTJLqEBM" ?
                        $signed((~^wire2696[(3'h5):(1'h0)])) : (&(!((wire2696 <= wire2692) ?
                            {wire2692} : (wire2696 ? wire2692 : wire2693)))));
  always
    @(posedge clk) begin
      reg2698 <= (&("ShTQ" ^~ $unsigned((wire2695 < {wire2695, (8'hb9)}))));
    end
  assign wire2699 = reg2698;
  always
    @(posedge clk) begin
      reg2700 <= "Pbr2VqGX5tJfhVaQ";
      reg2701 <= (($unsigned((~&wire2697[(5'h17):(1'h0)])) ?
              $signed($unsigned(reg2698)) : ("n3TX6Lst" ?
                  ("HuAs8Edc4e1cCUJc00KYB" ?
                      {wire2699} : $signed(wire2694)) : $signed({reg2698,
                      wire2697}))) ?
          $unsigned(($signed({reg2698}) ?
              wire2694 : {reg2698[(4'hf):(4'h9)]})) : wire2696[(4'hc):(2'h2)]);
      reg2702 = reg2698[(4'hf):(4'hb)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2592
#( parameter param2688 = ((((((8'hb6) ? (7'h47) : (8'hbc)) < {(8'hb7)}) >= (^((8'hb9) ? (8'ha6) : (7'h49)))) ? ((8'hb8) * (~^((8'ha9) != (8'haa)))) : (~&(7'h4a))) ? ({{(~(8'ha9))}} ^~ ((((8'ha7) <<< (8'hb1)) >= ((8'hbd) ? (8'h9d) : (8'hb8))) ? ({(8'ha3), (8'hb9)} ? ((8'hab) ? (7'h4c) : (8'hbd)) : ((8'hb1) <<< (8'ha4))) : (|((8'h9f) + (7'h4c))))) : (8'hab)) )
(y, clk, wire2596, wire2595, wire2594, wire2593);
  output wire [(32'h559):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire2596;
  input wire signed [(5'h11):(1'h0)] wire2595;
  input wire [(5'h10):(1'h0)] wire2594;
  input wire signed [(2'h3):(1'h0)] wire2593;
  reg signed [(5'h19):(1'h0)] reg2687 = (1'h0);
  reg [(4'he):(1'h0)] reg2686 = (1'h0);
  reg [(4'hc):(1'h0)] reg2685 = (1'h0);
  reg [(5'h15):(1'h0)] reg2684 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2683 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2682 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2681 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2680 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2679 = (1'h0);
  reg [(5'h14):(1'h0)] forvar2678 = (1'h0);
  reg [(5'h12):(1'h0)] reg2677 = (1'h0);
  reg [(5'h11):(1'h0)] reg2676 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2675 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2674 = (1'h0);
  reg [(3'h7):(1'h0)] reg2673 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2672 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2671 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2670 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2669 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2668 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2667 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2666 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2665 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2664 = (1'h0);
  reg [(2'h2):(1'h0)] reg2663 = (1'h0);
  reg [(5'h15):(1'h0)] forvar2662 = (1'h0);
  reg [(4'hb):(1'h0)] reg2661 = (1'h0);
  reg [(3'h5):(1'h0)] reg2660 = (1'h0);
  reg [(5'h16):(1'h0)] reg2659 = (1'h0);
  reg [(3'h6):(1'h0)] reg2658 = (1'h0);
  reg [(3'h7):(1'h0)] reg2657 = (1'h0);
  reg [(5'h11):(1'h0)] reg2656 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2655 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2654 = (1'h0);
  reg [(4'he):(1'h0)] reg2653 = (1'h0);
  reg [(5'h17):(1'h0)] reg2652 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2651 = (1'h0);
  reg [(5'h11):(1'h0)] reg2650 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2649 = (1'h0);
  reg [(5'h12):(1'h0)] reg2648 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2647 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2646 = (1'h0);
  reg [(5'h10):(1'h0)] reg2645 = (1'h0);
  reg [(5'h17):(1'h0)] reg2644 = (1'h0);
  reg [(5'h18):(1'h0)] reg2643 = (1'h0);
  reg [(5'h14):(1'h0)] reg2642 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2641 = (1'h0);
  reg [(5'h12):(1'h0)] reg2640 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2639 = (1'h0);
  reg [(3'h6):(1'h0)] reg2638 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2637 = (1'h0);
  reg [(5'h11):(1'h0)] reg2636 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2635 = (1'h0);
  reg [(3'h6):(1'h0)] reg2634 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2633 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2632 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2631 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2630 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2629 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2628 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2627 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2626 = (1'h0);
  reg [(5'h18):(1'h0)] reg2625 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2624 = (1'h0);
  reg [(4'hb):(1'h0)] reg2623 = (1'h0);
  reg [(4'he):(1'h0)] reg2622 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2621 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2620 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2619 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar2618 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar2617 = (1'h0);
  reg [(3'h4):(1'h0)] reg2616 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2615 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2614 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2613 = (1'h0);
  wire signed [(5'h16):(1'h0)] wire2612;
  reg [(4'he):(1'h0)] reg2611 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2610 = (1'h0);
  reg [(5'h18):(1'h0)] reg2609 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2608 = (1'h0);
  reg [(2'h3):(1'h0)] reg2607 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2606 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar2605 = (1'h0);
  reg [(5'h18):(1'h0)] reg2604 = (1'h0);
  reg [(3'h4):(1'h0)] reg2603 = (1'h0);
  reg [(5'h18):(1'h0)] forvar2602 = (1'h0);
  reg [(4'he):(1'h0)] forvar2601 = (1'h0);
  reg [(4'h8):(1'h0)] reg2600 = (1'h0);
  reg [(5'h15):(1'h0)] reg2599 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2598 = (1'h0);
  reg [(3'h5):(1'h0)] reg2597 = (1'h0);
  assign y = {reg2687,
                 reg2686,
                 reg2685,
                 reg2684,
                 reg2683,
                 reg2682,
                 reg2681,
                 reg2680,
                 reg2679,
                 forvar2678,
                 reg2677,
                 reg2676,
                 forvar2675,
                 reg2674,
                 reg2673,
                 reg2672,
                 reg2671,
                 reg2670,
                 reg2669,
                 reg2668,
                 reg2667,
                 reg2666,
                 reg2665,
                 reg2664,
                 reg2663,
                 forvar2662,
                 reg2661,
                 reg2660,
                 reg2659,
                 reg2658,
                 reg2657,
                 reg2656,
                 reg2655,
                 forvar2654,
                 reg2653,
                 reg2652,
                 reg2651,
                 reg2650,
                 reg2649,
                 reg2648,
                 reg2647,
                 forvar2646,
                 reg2645,
                 reg2644,
                 reg2643,
                 reg2642,
                 forvar2641,
                 reg2640,
                 forvar2639,
                 reg2638,
                 forvar2637,
                 reg2636,
                 reg2635,
                 reg2634,
                 reg2633,
                 reg2632,
                 reg2631,
                 reg2630,
                 reg2629,
                 forvar2628,
                 reg2627,
                 forvar2626,
                 reg2625,
                 reg2624,
                 reg2623,
                 reg2622,
                 reg2621,
                 reg2620,
                 reg2619,
                 forvar2618,
                 forvar2617,
                 reg2616,
                 forvar2615,
                 reg2614,
                 reg2613,
                 wire2612,
                 reg2611,
                 reg2610,
                 reg2609,
                 reg2608,
                 reg2607,
                 reg2606,
                 forvar2605,
                 reg2604,
                 reg2603,
                 forvar2602,
                 forvar2601,
                 reg2600,
                 reg2599,
                 reg2598,
                 reg2597,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg2597 <= wire2596[(3'h6):(1'h1)];
      reg2598 = $signed($unsigned(wire2596[(1'h0):(1'h0)]));
      reg2599 <= ($unsigned($unsigned(((~|wire2593) && {reg2598}))) != $signed(reg2597));
      reg2600 <= "3v";
      for (forvar2601 = (1'h0); (forvar2601 < (2'h3)); forvar2601 = (forvar2601 + (1'h1)))
        begin
          for (forvar2602 = (1'h0); (forvar2602 < (2'h3)); forvar2602 = (forvar2602 + (1'h1)))
            begin
              reg2603 <= ($signed((wire2593 ?
                  $signed($signed(forvar2602)) : ($unsigned(wire2593) - (8'ha0)))) * "c69XJ0d");
              reg2604 <= {{wire2596[(2'h2):(1'h1)],
                      (~&($unsigned(reg2600) == (reg2598 ?
                          wire2596 : wire2594)))},
                  $signed($unsigned((8'hb3)))};
            end
          for (forvar2605 = (1'h0); (forvar2605 < (3'h4)); forvar2605 = (forvar2605 + (1'h1)))
            begin
              reg2606 <= $unsigned(reg2600[(2'h2):(1'h1)]);
              reg2607 <= ("dNgifDamc0FCKT4DIsO" ?
                  $unsigned("yOYhJydZDfF") : (((reg2603 + (forvar2601 ?
                          reg2606 : forvar2601)) == reg2599[(4'he):(3'h5)]) ?
                      $signed($signed(forvar2601[(3'h4):(3'h4)])) : (~&(^~$signed(reg2597)))));
              reg2608 <= $signed((8'hbc));
              reg2609 <= $signed((~|((8'ha9) ?
                  $signed({reg2599}) : $unsigned(reg2600[(2'h2):(1'h0)]))));
            end
          reg2610 <= $signed("gd8t95r2gBwo6E5yxuQ");
        end
      reg2611 = "UXScG2mUtzFd5l";
    end
  assign wire2612 = $signed((-(|$unsigned(((8'hb5) == wire2594)))));
  always
    @(posedge clk) begin
      reg2613 <= $unsigned((8'ha3));
      reg2614 = $signed((^~({(wire2596 ?
              wire2596 : (8'hb8))} ^~ $unsigned((reg2611 ?
          (7'h43) : reg2598)))));
      for (forvar2615 = (1'h0); (forvar2615 < (1'h0)); forvar2615 = (forvar2615 + (1'h1)))
        begin
          reg2616 <= reg2599[(4'hf):(4'ha)];
          for (forvar2617 = (1'h0); (forvar2617 < (1'h0)); forvar2617 = (forvar2617 + (1'h1)))
            begin
              for (forvar2618 = (1'h0); (forvar2618 < (2'h2)); forvar2618 = (forvar2618 + (1'h1)))
                begin
                  reg2619 <= ((~(wire2594 ?
                          (-$unsigned(wire2593)) : reg2598[(1'h1):(1'h1)])) ?
                      (+reg2606) : ((-"rpH6ahq9pkeihHs") ^ forvar2601));
                  reg2620 <= (forvar2615[(1'h0):(1'h0)] <= "bckBYarJ");
                  reg2621 <= (~{(8'ha0),
                      ((^~(wire2593 ? forvar2602 : (7'h47))) & ((^reg2606) ?
                          reg2613 : (8'hbd)))});
                  reg2622 <= $unsigned(reg2619[(2'h2):(1'h0)]);
                  reg2623 <= forvar2602;
                  reg2624 <= forvar2602[(3'h7):(3'h6)];
                end
            end
          reg2625 = ((~wire2593) * $unsigned("pWme0HPf1JhHMgQSBJ"));
          for (forvar2626 = (1'h0); (forvar2626 < (1'h0)); forvar2626 = (forvar2626 + (1'h1)))
            begin
              reg2627 = reg2610;
              for (forvar2628 = (1'h0); (forvar2628 < (2'h3)); forvar2628 = (forvar2628 + (1'h1)))
                begin
                  reg2629 <= $signed($unsigned(((&$signed((7'h49))) < ((^(7'h43)) > (&reg2603)))));
                  reg2630 <= reg2613[(5'h16):(4'h8)];
                  reg2631 <= ("hb8LXapvs996Jramy" <<< ({reg2624[(1'h0):(1'h0)],
                      (~|(^(8'ha0)))} ^~ (~|$signed((&reg2623)))));
                  reg2632 <= reg2621[(1'h0):(1'h0)];
                  reg2633 = $signed("B0cOJ3u");
                  reg2634 = (("JqwrT" ?
                      $signed(reg2608[(1'h1):(1'h1)]) : reg2620[(4'h8):(3'h5)]) || $unsigned((~|$signed(forvar2626[(3'h7):(3'h4)]))));
                end
              reg2635 <= (-forvar2615[(1'h1):(1'h1)]);
            end
          reg2636 <= (({reg2625[(3'h6):(1'h0)]} ?
              (((reg2634 ?
                  reg2598 : reg2599) ^~ reg2598) >>> "nLQ6rFzR") : $signed(((~|forvar2617) ?
                  "1W1mXf" : {(7'h43), reg2599}))) <<< $signed("Zl8qS8f"));
        end
      for (forvar2637 = (1'h0); (forvar2637 < (2'h2)); forvar2637 = (forvar2637 + (1'h1)))
        begin
          reg2638 <= ((reg2621 ?
                  $signed(forvar2626[(4'hd):(4'ha)]) : wire2612[(1'h0):(1'h0)]) ?
              (wire2595[(3'h7):(2'h3)] | {{(+reg2620)}}) : {$signed((^(&reg2633))),
                  ("Xm0qfivqKVRaz75d" <<< ((reg2633 ? wire2595 : reg2634) ?
                      (&reg2629) : $signed(wire2596)))});
          for (forvar2639 = (1'h0); (forvar2639 < (3'h5)); forvar2639 = (forvar2639 + (1'h1)))
            begin
              reg2640 <= ((+(reg2600 || (|reg2625))) ?
                  reg2638 : reg2638[(2'h3):(1'h1)]);
              for (forvar2641 = (1'h0); (forvar2641 < (3'h4)); forvar2641 = (forvar2641 + (1'h1)))
                begin
                  reg2642 <= "JI3";
                  reg2643 = reg2625[(5'h18):(4'h8)];
                  reg2644 = forvar2639[(3'h5):(2'h2)];
                  reg2645 = $unsigned($unsigned($signed((~&wire2596))));
                end
              for (forvar2646 = (1'h0); (forvar2646 < (2'h2)); forvar2646 = (forvar2646 + (1'h1)))
                begin
                  reg2647 <= (((~|{(reg2632 <= reg2627),
                          $unsigned(forvar2605)}) ?
                      reg2638 : ("NnE6ee3UPoS3v1" ?
                          ({reg2599} ?
                              (forvar2628 <<< reg2604) : (reg2623 ?
                                  reg2629 : (8'h9f))) : reg2644[(4'he):(4'ha)])) ~^ $unsigned(forvar2601));
                  reg2648 = forvar2605;
                  reg2649 <= (~|(7'h42));
                  reg2650 <= $unsigned(reg2644[(4'hb):(1'h1)]);
                  reg2651 <= ((~^$unsigned(($signed(reg2648) & {reg2631,
                          (8'hb5)}))) ?
                      reg2598 : (-forvar2615));
                  reg2652 <= reg2629;
                end
              reg2653 <= (~^(({"gelnWIpEGYlxFVExGLlGkd",
                      $unsigned(reg2614)} & $signed({(8'ha2)})) ?
                  (^~"wCG63zwEgV9C") : "4d9ufLUKGF0Ki"));
            end
          for (forvar2654 = (1'h0); (forvar2654 < (1'h0)); forvar2654 = (forvar2654 + (1'h1)))
            begin
              reg2655 <= (~reg2616);
              reg2656 <= forvar2618[(4'he):(2'h3)];
              reg2657 <= (forvar2618[(4'hb):(1'h0)] ?
                  $unsigned("2ElPG2OYi") : (reg2603[(3'h4):(1'h0)] <<< $unsigned((((7'h4c) >>> reg2620) || (~forvar2646)))));
              reg2658 <= reg2651[(1'h0):(1'h0)];
              reg2659 <= (|(($unsigned(reg2620) <= ((reg2638 || (8'ha4)) ?
                  reg2607 : {reg2635,
                      reg2643})) > (forvar2601 && (reg2619[(2'h3):(2'h3)] != reg2657[(3'h4):(1'h0)]))));
              reg2660 <= $signed("");
            end
          reg2661 <= wire2596[(1'h0):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar2662 = (1'h0); (forvar2662 < (1'h0)); forvar2662 = (forvar2662 + (1'h1)))
        begin
          reg2663 <= "i37XdIa6U2";
        end
      reg2664 <= (~^(&{({reg2638, reg2640} <= (forvar2601 ? reg2651 : reg2659)),
          reg2643}));
      if ((!reg2655[(5'h17):(4'ha)]))
        begin
          reg2665 <= {($unsigned($signed(wire2612[(5'h12):(4'ha)])) ?
                  $unsigned($signed($unsigned((7'h45)))) : forvar2615)};
        end
      else
        begin
          reg2665 <= ((reg2635[(2'h2):(1'h1)] * $signed((reg2640 ?
              (reg2606 ?
                  reg2633 : forvar2602) : $unsigned(forvar2641)))) <<< (($signed((forvar2605 ?
              reg2653 : forvar2605)) <= $signed((reg2657 ?
              wire2596 : reg2607))) & (8'hba)));
          reg2666 <= (&$signed("ZSvD"));
          reg2667 <= ($unsigned($signed("DZpgvL")) | ((reg2597[(1'h0):(1'h0)] ?
              $signed((reg2606 > (7'h49))) : (8'hbf)) ^~ (!$signed($signed((7'h42))))));
        end
      reg2668 <= $signed("qiKTlrrfxKX");
      reg2669 <= reg2606[(5'h10):(2'h3)];
      reg2670 <= "pstFEuH0";
    end
  always
    @(posedge clk) begin
      reg2671 <= ({$signed(reg2647)} > "wSbP7TouZm658p8");
      reg2672 <= {$signed("hdUWo60E5FsnJPrZ5nN")};
      reg2673 = $signed(($signed("D07Vo6yg") * reg2647[(2'h3):(2'h2)]));
      reg2674 <= $unsigned(($signed(reg2632[(4'hc):(3'h5)]) ?
          $unsigned($signed("Hoa6JT6alL0Z1d1")) : ((~^reg2649[(2'h2):(1'h1)]) ?
              {(wire2594 && (7'h41))} : $unsigned((~^(7'h46))))));
    end
  always
    @(posedge clk) begin
      for (forvar2675 = (1'h0); (forvar2675 < (1'h0)); forvar2675 = (forvar2675 + (1'h1)))
        begin
          reg2676 <= reg2664;
          reg2677 = ($unsigned(($unsigned((~&reg2642)) || "hRWFGw2rsnRDhOePzXmi")) <<< ($unsigned("UrS") ^ {(-"QifZmXNYQkGcIwU4ac7")}));
          for (forvar2678 = (1'h0); (forvar2678 < (2'h3)); forvar2678 = (forvar2678 + (1'h1)))
            begin
              reg2679 <= reg2609;
            end
          reg2680 <= (8'hb6);
          reg2681 <= (!"8K0SIFiOzNRhOF5lB");
        end
      reg2682 <= ((-($signed(reg2640) != ((!reg2627) ?
              {reg2629, reg2606} : ((7'h48) == forvar2618)))) ?
          (($unsigned((forvar2678 ? reg2616 : reg2666)) ?
                  ($unsigned(reg2676) <= (8'hb4)) : $signed((~^forvar2602))) ?
              ((8'ha4) ?
                  wire2612[(3'h4):(1'h0)] : reg2671) : ((~^reg2610) >> $signed((reg2630 ?
                  (7'h4b) : forvar2662)))) : wire2594);
      reg2683 = $signed("ce5sZfHMLKzS");
      reg2684 = ("HcHLR4" || {{reg2633[(4'h8):(4'h8)],
              $signed((reg2598 + reg2682))}});
    end
  always
    @(posedge clk) begin
      reg2685 <= {"v5y9cl", ("WSUhIx0XSBpdu8wyD" ^~ reg2682)};
      reg2686 <= $signed($unsigned((~|$signed(reg2657))));
      reg2687 <= reg2665;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2538
#( parameter param2588 = {((|(~^(~&(8'hb4)))) != ((8'hbe) ^ (8'hba)))}
, parameter param2589 = {(!({(~&param2588)} ? (~&(&param2588)) : ((^~param2588) ? (^~param2588) : (param2588 << param2588))))} )
(y, clk, wire2543, wire2542, wire2541, wire2540, wire2539);
  output wire [(32'h278):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h17):(1'h0)] wire2543;
  input wire [(5'h15):(1'h0)] wire2542;
  input wire signed [(3'h6):(1'h0)] wire2541;
  input wire signed [(4'hf):(1'h0)] wire2540;
  input wire signed [(5'h14):(1'h0)] wire2539;
  reg signed [(5'h14):(1'h0)] reg2587 = (1'h0);
  reg [(5'h12):(1'h0)] reg2586 = (1'h0);
  reg [(3'h6):(1'h0)] reg2585 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2584 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2583 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2582 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2581 = (1'h0);
  reg [(3'h5):(1'h0)] reg2580 = (1'h0);
  reg [(5'h10):(1'h0)] reg2579 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2578 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2577 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2576 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2575 = (1'h0);
  reg [(5'h11):(1'h0)] reg2574 = (1'h0);
  reg [(4'he):(1'h0)] reg2573 = (1'h0);
  reg [(3'h7):(1'h0)] reg2572 = (1'h0);
  reg [(4'ha):(1'h0)] reg2571 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2570 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2569 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2568 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2567 = (1'h0);
  wire [(4'hc):(1'h0)] wire2566;
  wire signed [(4'h9):(1'h0)] wire2565;
  wire [(4'hb):(1'h0)] wire2564;
  wire [(5'h10):(1'h0)] wire2563;
  wire signed [(5'h11):(1'h0)] wire2562;
  wire signed [(5'h18):(1'h0)] wire2561;
  reg [(4'hd):(1'h0)] reg2560 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2559 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2558 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2557 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2556 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2555 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2554 = (1'h0);
  reg [(3'h6):(1'h0)] reg2553 = (1'h0);
  reg [(5'h12):(1'h0)] reg2552 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2551 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2545 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2550 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2549 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2548 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2547 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2546 = (1'h0);
  reg [(4'hd):(1'h0)] reg2545 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2544 = (1'h0);
  assign y = {reg2587,
                 reg2586,
                 reg2585,
                 reg2584,
                 reg2583,
                 reg2582,
                 reg2581,
                 reg2580,
                 reg2579,
                 forvar2578,
                 reg2577,
                 reg2576,
                 reg2575,
                 reg2574,
                 reg2573,
                 reg2572,
                 reg2571,
                 reg2570,
                 forvar2569,
                 forvar2568,
                 forvar2567,
                 wire2566,
                 wire2565,
                 wire2564,
                 wire2563,
                 wire2562,
                 wire2561,
                 reg2560,
                 reg2559,
                 reg2558,
                 reg2557,
                 reg2556,
                 reg2555,
                 forvar2554,
                 reg2553,
                 reg2552,
                 reg2551,
                 forvar2545,
                 reg2550,
                 reg2549,
                 reg2548,
                 reg2547,
                 reg2546,
                 reg2545,
                 forvar2544,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar2544 = (1'h0); (forvar2544 < (3'h4)); forvar2544 = (forvar2544 + (1'h1)))
        begin
          if ({$unsigned((|$unsigned(wire2539))), (|(8'ha6))})
            begin
              reg2545 <= (wire2540 >> "g8gP");
              reg2546 <= (|$unsigned({$unsigned($signed(wire2542)), "5i"}));
              reg2547 <= $signed((+reg2545));
              reg2548 <= (8'hab);
              reg2549 <= reg2548;
              reg2550 <= $unsigned({(((&reg2548) ?
                          (wire2541 && reg2548) : ((8'hb4) ?
                              reg2549 : (8'ha7))) ?
                      (reg2549[(4'hc):(4'h8)] - (forvar2544 * wire2541)) : reg2546[(4'h8):(2'h2)]),
                  $signed(((~|(8'hbe)) ? "bsCSF0d9ZI5ALu9e" : (~&wire2543)))});
            end
          else
            begin
              for (forvar2545 = (1'h0); (forvar2545 < (3'h4)); forvar2545 = (forvar2545 + (1'h1)))
                begin
                  reg2546 <= (reg2545[(4'ha):(3'h6)] ?
                      (wire2541[(3'h4):(1'h1)] != $unsigned("RraIrZlSXG2rPuW0SN5rB")) : $signed({$unsigned((reg2546 ^~ reg2547)),
                          wire2539[(1'h1):(1'h1)]}));
                  reg2547 <= "sT9zamTbrxtkqqBC9fMZ";
                  reg2548 = (((((!reg2547) << forvar2545[(3'h7):(3'h6)]) <= $signed(((7'h4d) ^ reg2547))) ?
                      reg2550[(4'h8):(1'h1)] : {reg2546[(5'h16):(4'h8)]}) <<< "4DpdR2VSY");
                  reg2549 = ((reg2550 >> reg2546[(1'h1):(1'h1)]) ?
                      wire2541 : "Ju2Bgsa");
                  reg2550 <= (({((8'ha4) ?
                          $signed(wire2539) : (reg2547 >> wire2541)),
                      $unsigned(wire2540[(4'hb):(4'h9)])} >> "2iV5K7e1UE0") >= {reg2546[(5'h15):(3'h4)]});
                  reg2551 <= (reg2550[(4'ha):(3'h4)] & $signed(forvar2544));
                end
              reg2552 = ($unsigned($signed($unsigned((forvar2544 && reg2550)))) ?
                  $signed(((reg2550 ?
                      $signed(forvar2545) : wire2541) & wire2540[(3'h4):(3'h4)])) : "H1Yv");
              reg2553 <= reg2545[(3'h7):(1'h0)];
              for (forvar2554 = (1'h0); (forvar2554 < (2'h3)); forvar2554 = (forvar2554 + (1'h1)))
                begin
                  reg2555 = "dwsu5Mkz8";
                end
            end
          reg2556 <= ($unsigned(forvar2545) ?
              ((^~$unsigned((reg2550 ?
                  wire2540 : reg2549))) ~^ reg2553[(3'h5):(3'h4)]) : reg2547);
          reg2557 <= $unsigned(({reg2545, reg2551[(3'h5):(3'h4)]} ?
              $signed($unsigned(reg2555[(4'h8):(3'h4)])) : reg2545));
          reg2558 <= (~reg2548[(2'h2):(2'h2)]);
          reg2559 <= "qtlBB8fP3CWg6zJVBCs2EPeJ";
          reg2560 <= $unsigned((-(~|(+"U0LkAmc0C30H"))));
        end
    end
  assign wire2561 = ((~"nCYWzT1k30pmGMQK") << "CsYsK9o");
  assign wire2562 = $unsigned("gS");
  assign wire2563 = $signed($signed($unsigned("apvtDQAV")));
  assign wire2564 = reg2550[(5'h11):(2'h2)];
  assign wire2565 = $unsigned((^(~^wire2561)));
  assign wire2566 = "hw";
  always
    @(posedge clk) begin
      for (forvar2567 = (1'h0); (forvar2567 < (1'h0)); forvar2567 = (forvar2567 + (1'h1)))
        begin
          for (forvar2568 = (1'h0); (forvar2568 < (2'h3)); forvar2568 = (forvar2568 + (1'h1)))
            begin
              for (forvar2569 = (1'h0); (forvar2569 < (3'h4)); forvar2569 = (forvar2569 + (1'h1)))
                begin
                  reg2570 <= {wire2542,
                      ("VOlWsy1wUJWIdyYOo" ?
                          wire2542 : (&((reg2556 ? reg2548 : (8'hbb)) ?
                              (forvar2569 < (8'hb1)) : reg2559[(2'h3):(2'h3)])))};
                  reg2571 = wire2564;
                  reg2572 <= (~^("VCBP69gyK9" ?
                      forvar2568[(2'h3):(2'h3)] : wire2564[(1'h0):(1'h0)]));
                  reg2573 <= $signed("S53ML1");
                end
              reg2574 = (|reg2555);
              reg2575 <= ($signed(wire2539[(1'h0):(1'h0)]) && "Hpal2QE2f5CKIN3Fw");
              reg2576 <= reg2573[(1'h0):(1'h0)];
            end
          reg2577 <= {{reg2546, forvar2567[(4'h8):(3'h5)]}};
          for (forvar2578 = (1'h0); (forvar2578 < (2'h2)); forvar2578 = (forvar2578 + (1'h1)))
            begin
              reg2579 <= reg2571[(3'h4):(3'h4)];
              reg2580 <= wire2561;
              reg2581 <= $signed("3Lg3ChU");
              reg2582 <= $unsigned((~(~|reg2580)));
            end
        end
      reg2583 <= $signed($signed(({$unsigned(reg2575)} * forvar2568)));
      reg2584 <= {(~(((~reg2559) + (7'h4c)) ?
              (wire2543 == $unsigned(forvar2568)) : forvar2545[(5'h18):(5'h18)]))};
      reg2585 <= forvar2568;
      reg2586 <= (($unsigned(((forvar2568 > reg2553) ?
              $unsigned(reg2546) : {(7'h46)})) ~^ (+((8'ha2) & (|reg2576)))) ?
          $signed({"pp"}) : (((+(reg2545 ? wire2543 : reg2583)) ?
                  reg2549[(4'ha):(3'h7)] : wire2543) ?
              (((|(8'hb5)) ?
                  (reg2552 ? reg2583 : reg2581) : (forvar2545 ?
                      reg2575 : reg2581)) * ($unsigned((7'h4e)) && "MHzQPdfhoCCW2whThgaxkH")) : $signed("mPBkiQExXzT4E0H48qUOoXYD")));
      reg2587 <= "ioqg4Z9tU72BM4LakJV";
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2349  (y, clk, wire2353, wire2352, wire2351, wire2350);
  output wire [(32'h9ab):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire2353;
  input wire signed [(5'h10):(1'h0)] wire2352;
  input wire [(5'h19):(1'h0)] wire2351;
  input wire [(4'hf):(1'h0)] wire2350;
  reg signed [(3'h5):(1'h0)] reg2530 = (1'h0);
  reg [(4'hb):(1'h0)] reg2529 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2528 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2527 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2526 = (1'h0);
  reg [(5'h18):(1'h0)] reg2525 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar2524 = (1'h0);
  reg [(5'h12):(1'h0)] forvar2523 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2522 = (1'h0);
  reg [(4'ha):(1'h0)] reg2521 = (1'h0);
  reg [(3'h6):(1'h0)] reg2520 = (1'h0);
  reg [(5'h19):(1'h0)] reg2519 = (1'h0);
  reg [(5'h15):(1'h0)] reg2518 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2517 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2516 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2515 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2514 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2513 = (1'h0);
  reg [(3'h5):(1'h0)] reg2512 = (1'h0);
  reg [(4'hb):(1'h0)] reg2511 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2510 = (1'h0);
  reg [(5'h13):(1'h0)] reg2509 = (1'h0);
  reg [(4'h8):(1'h0)] reg2508 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2507 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2506 = (1'h0);
  reg [(5'h10):(1'h0)] reg2505 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2504 = (1'h0);
  reg [(5'h15):(1'h0)] reg2503 = (1'h0);
  reg [(5'h18):(1'h0)] reg2502 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2501 = (1'h0);
  reg [(3'h5):(1'h0)] reg2500 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2499 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2498 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2497 = (1'h0);
  wire [(5'h11):(1'h0)] wire2496;
  reg signed [(5'h14):(1'h0)] reg2495 = (1'h0);
  reg [(3'h6):(1'h0)] reg2494 = (1'h0);
  reg [(2'h3):(1'h0)] reg2493 = (1'h0);
  reg [(2'h3):(1'h0)] reg2492 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2491 = (1'h0);
  reg [(2'h3):(1'h0)] reg2490 = (1'h0);
  reg [(5'h11):(1'h0)] reg2489 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2488 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2487 = (1'h0);
  reg [(3'h6):(1'h0)] reg2486 = (1'h0);
  reg [(5'h15):(1'h0)] reg2485 = (1'h0);
  reg [(4'hc):(1'h0)] reg2484 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2483 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2482 = (1'h0);
  reg [(4'he):(1'h0)] reg2481 = (1'h0);
  reg [(4'hd):(1'h0)] reg2480 = (1'h0);
  reg [(2'h2):(1'h0)] reg2479 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2478 = (1'h0);
  reg [(5'h19):(1'h0)] reg2477 = (1'h0);
  reg [(5'h19):(1'h0)] reg2476 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2475 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2474 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2473 = (1'h0);
  reg [(5'h16):(1'h0)] reg2472 = (1'h0);
  reg [(5'h18):(1'h0)] reg2471 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2470 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2469 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2468 = (1'h0);
  reg [(5'h11):(1'h0)] reg2467 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2466 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2465 = (1'h0);
  reg [(5'h15):(1'h0)] reg2464 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2463 = (1'h0);
  reg [(5'h12):(1'h0)] reg2462 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2461 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2460 = (1'h0);
  reg [(4'hb):(1'h0)] reg2442 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2459 = (1'h0);
  reg [(5'h14):(1'h0)] reg2458 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2457 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar2456 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2455 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2454 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2453 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2452 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2451 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2450 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2449 = (1'h0);
  reg [(5'h11):(1'h0)] reg2448 = (1'h0);
  reg [(2'h3):(1'h0)] reg2447 = (1'h0);
  reg [(5'h17):(1'h0)] reg2446 = (1'h0);
  reg [(5'h17):(1'h0)] reg2445 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2444 = (1'h0);
  reg [(3'h7):(1'h0)] reg2443 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2442 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2441 = (1'h0);
  reg [(5'h12):(1'h0)] reg2440 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2439 = (1'h0);
  reg [(5'h17):(1'h0)] reg2438 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2437 = (1'h0);
  reg [(5'h15):(1'h0)] reg2436 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2435 = (1'h0);
  reg [(5'h16):(1'h0)] reg2434 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2433 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2432 = (1'h0);
  reg [(5'h18):(1'h0)] reg2431 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2430 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2429 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2428 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2427 = (1'h0);
  reg [(5'h11):(1'h0)] reg2426 = (1'h0);
  reg [(5'h13):(1'h0)] reg2425 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2424 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2423 = (1'h0);
  reg [(5'h16):(1'h0)] reg2422 = (1'h0);
  wire signed [(5'h16):(1'h0)] wire2421;
  wire signed [(5'h17):(1'h0)] wire2420;
  reg signed [(3'h6):(1'h0)] reg2419 = (1'h0);
  reg [(4'hb):(1'h0)] reg2418 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2417 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2416 = (1'h0);
  reg [(4'h8):(1'h0)] reg2415 = (1'h0);
  reg [(3'h5):(1'h0)] reg2414 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2413 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2412 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2411 = (1'h0);
  reg [(3'h4):(1'h0)] reg2410 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2409 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2408 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2407 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2406 = (1'h0);
  reg [(4'hc):(1'h0)] reg2405 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2404 = (1'h0);
  reg [(5'h11):(1'h0)] reg2403 = (1'h0);
  reg [(4'ha):(1'h0)] reg2402 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2401 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2400 = (1'h0);
  reg [(3'h6):(1'h0)] reg2399 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2398 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2397 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2396 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2395 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2394 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2393 = (1'h0);
  reg [(5'h17):(1'h0)] forvar2392 = (1'h0);
  reg [(4'he):(1'h0)] reg2391 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2390 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2389 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2388 = (1'h0);
  reg [(4'hb):(1'h0)] reg2387 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2386 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2385 = (1'h0);
  reg [(2'h3):(1'h0)] reg2384 = (1'h0);
  reg [(5'h15):(1'h0)] reg2383 = (1'h0);
  wire [(4'hc):(1'h0)] wire2382;
  reg signed [(2'h2):(1'h0)] reg2381 = (1'h0);
  reg [(3'h7):(1'h0)] reg2380 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2379 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar2378 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2377 = (1'h0);
  reg [(4'hc):(1'h0)] reg2376 = (1'h0);
  reg [(2'h3):(1'h0)] reg2375 = (1'h0);
  reg [(4'ha):(1'h0)] reg2374 = (1'h0);
  reg [(4'he):(1'h0)] forvar2373 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2372 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2371 = (1'h0);
  reg [(5'h16):(1'h0)] reg2370 = (1'h0);
  reg [(5'h12):(1'h0)] reg2369 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2368 = (1'h0);
  reg [(4'hf):(1'h0)] reg2367 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2366 = (1'h0);
  reg [(5'h18):(1'h0)] reg2365 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2364 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2363 = (1'h0);
  reg [(3'h5):(1'h0)] reg2362 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2361 = (1'h0);
  reg [(4'hb):(1'h0)] reg2360 = (1'h0);
  reg [(3'h5):(1'h0)] reg2359 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2358 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2357 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2356 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar2354 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2355 = (1'h0);
  reg [(5'h10):(1'h0)] reg2354 = (1'h0);
  assign y = {reg2530,
                 reg2529,
                 reg2528,
                 reg2527,
                 reg2526,
                 reg2525,
                 forvar2524,
                 forvar2523,
                 reg2522,
                 reg2521,
                 reg2520,
                 reg2519,
                 reg2518,
                 reg2517,
                 reg2516,
                 reg2515,
                 forvar2514,
                 reg2513,
                 reg2512,
                 reg2511,
                 forvar2510,
                 reg2509,
                 reg2508,
                 reg2507,
                 reg2506,
                 reg2505,
                 reg2504,
                 reg2503,
                 reg2502,
                 forvar2501,
                 reg2500,
                 forvar2499,
                 reg2498,
                 reg2497,
                 wire2496,
                 reg2495,
                 reg2494,
                 reg2493,
                 reg2492,
                 reg2491,
                 reg2490,
                 reg2489,
                 reg2488,
                 reg2487,
                 reg2486,
                 reg2485,
                 reg2484,
                 reg2483,
                 forvar2482,
                 reg2481,
                 reg2480,
                 reg2479,
                 reg2478,
                 reg2477,
                 reg2476,
                 reg2475,
                 forvar2474,
                 reg2473,
                 reg2472,
                 reg2471,
                 reg2470,
                 reg2469,
                 reg2468,
                 reg2467,
                 reg2466,
                 forvar2465,
                 reg2464,
                 reg2463,
                 reg2462,
                 reg2461,
                 forvar2460,
                 reg2442,
                 reg2459,
                 reg2458,
                 reg2457,
                 forvar2456,
                 reg2455,
                 reg2454,
                 reg2453,
                 reg2452,
                 forvar2451,
                 reg2450,
                 forvar2449,
                 reg2448,
                 reg2447,
                 reg2446,
                 reg2445,
                 reg2444,
                 reg2443,
                 forvar2442,
                 reg2441,
                 reg2440,
                 reg2439,
                 reg2438,
                 forvar2437,
                 reg2436,
                 reg2435,
                 reg2434,
                 reg2433,
                 forvar2432,
                 reg2431,
                 reg2430,
                 forvar2429,
                 reg2428,
                 reg2427,
                 reg2426,
                 reg2425,
                 forvar2424,
                 reg2423,
                 reg2422,
                 wire2421,
                 wire2420,
                 reg2419,
                 reg2418,
                 reg2417,
                 reg2416,
                 reg2415,
                 reg2414,
                 forvar2413,
                 reg2412,
                 reg2411,
                 reg2410,
                 reg2409,
                 reg2408,
                 reg2407,
                 forvar2406,
                 reg2405,
                 reg2404,
                 reg2403,
                 reg2402,
                 reg2401,
                 reg2400,
                 reg2399,
                 reg2398,
                 reg2397,
                 reg2396,
                 reg2395,
                 forvar2394,
                 reg2393,
                 forvar2392,
                 reg2391,
                 forvar2390,
                 reg2389,
                 forvar2388,
                 reg2387,
                 reg2386,
                 reg2385,
                 reg2384,
                 reg2383,
                 wire2382,
                 reg2381,
                 reg2380,
                 reg2379,
                 forvar2378,
                 reg2377,
                 reg2376,
                 reg2375,
                 reg2374,
                 forvar2373,
                 forvar2372,
                 reg2371,
                 reg2370,
                 reg2369,
                 reg2368,
                 reg2367,
                 forvar2366,
                 reg2365,
                 reg2364,
                 reg2363,
                 reg2362,
                 reg2361,
                 reg2360,
                 reg2359,
                 reg2358,
                 reg2357,
                 reg2356,
                 forvar2354,
                 reg2355,
                 reg2354,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($signed(wire2350[(2'h3):(2'h3)]))
        begin
          reg2354 <= "ZZHSwSO4kpzmel7zARNot";
          reg2355 <= $unsigned("dl7TyHQYeEZJtROnNuAQ4G3");
        end
      else
        begin
          for (forvar2354 = (1'h0); (forvar2354 < (2'h2)); forvar2354 = (forvar2354 + (1'h1)))
            begin
              reg2355 <= $signed($unsigned(((+$signed((8'hbf))) >= $signed((wire2352 <= wire2350)))));
              reg2356 = ("dygPd271CB6ot" <= {$signed($signed(wire2351[(5'h13):(3'h6)]))});
              reg2357 <= $signed("UUe");
              if ($signed(($signed(($unsigned(forvar2354) << (|reg2356))) ~^ reg2357[(5'h11):(4'ha)])))
                begin
                  reg2358 <= (~&$signed($signed(((^~reg2354) ?
                      (reg2354 + reg2355) : "pHNmmAlHVaaOaXZnvla7PYW"))));
                  reg2359 = $unsigned($signed(("1J3LRpsexrWDn9QR2ZzNo" ?
                      wire2350[(4'h8):(1'h1)] : (|{wire2353}))));
                  reg2360 = wire2351;
                  reg2361 = $signed($unsigned(wire2352[(4'ha):(2'h2)]));
                  reg2362 <= reg2355;
                  reg2363 <= reg2355[(3'h5):(3'h5)];
                end
              else
                begin
                  reg2358 <= "gnghzr3UmaWFsToB8UDf";
                  reg2359 = $unsigned(((($signed(reg2356) ?
                      reg2358 : (~^reg2360)) < (wire2353 ?
                      {reg2358,
                          reg2363} : (reg2358 < reg2355))) >= $unsigned($unsigned({wire2353}))));
                  reg2360 <= {((8'hbd) + $unsigned(($signed((7'h4c)) ?
                          reg2363 : reg2358)))};
                  reg2361 <= "nGYbfbx8dugFdvy4XR6zV";
                  reg2362 = reg2358;
                end
              reg2364 <= (reg2357[(2'h2):(2'h2)] < $signed($signed(reg2363)));
              reg2365 <= (($signed((reg2364[(3'h6):(2'h2)] ?
                      (reg2358 ? (8'h9f) : reg2355) : (wire2352 ?
                          reg2359 : wire2350))) || reg2357) ?
                  wire2353 : (^$signed(reg2354)));
            end
          for (forvar2366 = (1'h0); (forvar2366 < (2'h2)); forvar2366 = (forvar2366 + (1'h1)))
            begin
              reg2367 <= (((-((reg2354 << forvar2354) ?
                          reg2354 : $unsigned(wire2351))) ?
                      wire2351 : "23ZAMqH6R0b78GI") ?
                  ((reg2365 ?
                          $signed((^~wire2351)) : $signed((wire2351 ^ reg2357))) ?
                      $signed($signed(reg2363[(5'h17):(3'h6)])) : $signed(((reg2363 <<< reg2363) ^~ (wire2351 < wire2350)))) : wire2353);
              reg2368 <= $unsigned(reg2356[(3'h6):(1'h0)]);
              reg2369 <= $signed(($unsigned("S1SzefaRCl9uv7beu3") ?
                  (($unsigned(reg2362) * $unsigned(reg2365)) >= ((reg2360 | reg2362) ?
                      reg2355 : "hae")) : (~^$unsigned({reg2367, reg2358}))));
              reg2370 = $signed(($unsigned(reg2362[(2'h2):(2'h2)]) ?
                  $signed("") : ((8'had) - (wire2353 ?
                      $unsigned(reg2367) : reg2364[(3'h6):(3'h4)]))));
              reg2371 <= wire2351[(3'h7):(3'h7)];
            end
        end
      for (forvar2372 = (1'h0); (forvar2372 < (3'h4)); forvar2372 = (forvar2372 + (1'h1)))
        begin
          for (forvar2373 = (1'h0); (forvar2373 < (1'h0)); forvar2373 = (forvar2373 + (1'h1)))
            begin
              reg2374 = ((reg2370[(5'h15):(4'hf)] >= ($signed((~wire2350)) ?
                      $unsigned({(7'h44)}) : reg2371[(1'h1):(1'h0)])) ?
                  (|reg2370[(4'h8):(4'h8)]) : $signed(wire2353[(1'h0):(1'h0)]));
              reg2375 <= {$signed("8Ruw69yeJ6bcUPSmPTYt1G9")};
              reg2376 <= wire2353;
              reg2377 <= "uQi8ky4";
              for (forvar2378 = (1'h0); (forvar2378 < (1'h1)); forvar2378 = (forvar2378 + (1'h1)))
                begin
                  reg2379 = (({wire2352[(2'h2):(2'h2)]} || (({reg2374} ?
                      $unsigned(reg2376) : $signed(reg2360)) * ($signed(reg2365) - ""))) >> (-$unsigned((~((8'hb7) ?
                      (8'haf) : wire2351)))));
                end
            end
          reg2380 <= {forvar2378[(5'h11):(2'h3)],
              (~((((8'h9f) ? reg2361 : reg2375) | "ACU") == reg2368))};
          reg2381 = (8'haa);
        end
    end
  assign wire2382 = (8'h9c);
  always
    @(posedge clk) begin
      reg2383 <= reg2364;
      reg2384 <= (($unsigned("6r557KhNNBVEPdL7chM0RpK") ?
          $unsigned(((^reg2371) ~^ (^(7'h48)))) : {$signed((7'h48))}) < reg2370[(5'h15):(5'h12)]);
    end
  always
    @(posedge clk) begin
      reg2385 <= ($unsigned(("iSrOmPDrGO" == $unsigned("fbuYu88fK2pQhb"))) >= {"",
          (reg2362 << (reg2369 <<< $unsigned((8'ha2))))});
      reg2386 <= reg2370[(3'h6):(3'h6)];
      reg2387 = $signed(reg2356[(5'h10):(3'h5)]);
      for (forvar2388 = (1'h0); (forvar2388 < (2'h2)); forvar2388 = (forvar2388 + (1'h1)))
        begin
          reg2389 <= (~&reg2384[(2'h3):(1'h0)]);
          for (forvar2390 = (1'h0); (forvar2390 < (2'h3)); forvar2390 = (forvar2390 + (1'h1)))
            begin
              reg2391 <= (!(|reg2360));
            end
          for (forvar2392 = (1'h0); (forvar2392 < (1'h0)); forvar2392 = (forvar2392 + (1'h1)))
            begin
              reg2393 <= $signed({{reg2361[(3'h7):(1'h0)], reg2385}, ""});
              for (forvar2394 = (1'h0); (forvar2394 < (1'h0)); forvar2394 = (forvar2394 + (1'h1)))
                begin
                  reg2395 <= $unsigned($signed((8'hbb)));
                  reg2396 <= $signed(wire2351);
                  reg2397 <= {{("Aqanz3d" ? (+(|reg2363)) : "M1k6mS"),
                          "KywukGlGu9b6qMMEdKmA"}};
                  reg2398 <= ((reg2383[(5'h14):(4'ha)] ?
                          (~&"sy2dtzKCTJMqisL5ZltMK") : $unsigned(({(8'haf),
                                  reg2354} ?
                              ((8'hbb) ? wire2353 : reg2379) : {reg2355}))) ?
                      (-"QMBoqa2AA") : "gRi7MiHqku");
                end
              reg2399 = (|(~|forvar2354));
            end
          reg2400 <= "k7FWY5C";
          reg2401 <= (^(reg2380[(3'h5):(3'h4)] >= (!$signed((reg2355 ?
              reg2370 : reg2398)))));
        end
      reg2402 <= ($unsigned(reg2395[(4'h8):(1'h1)]) ?
          $unsigned((~^("rg5cILZ32J4C705JpIBPaZl2" ?
              $unsigned(wire2350) : (+forvar2392)))) : $signed((reg2363[(1'h1):(1'h0)] ?
              (~&$signed(reg2384)) : forvar2373[(2'h2):(1'h0)])));
      reg2403 <= ((~wire2350[(3'h5):(1'h1)]) ?
          $signed($unsigned("X6bx4qfAYNGOOowdQBG7")) : (reg2399 ?
              {reg2402[(3'h5):(2'h3)]} : wire2352[(1'h0):(1'h0)]));
    end
  always
    @(posedge clk) begin
      reg2404 = (forvar2373 >= (($unsigned(reg2391[(3'h7):(2'h2)]) ?
              $signed((reg2383 ? reg2389 : reg2389)) : (~(reg2398 & reg2361))) ?
          (reg2400 - "1Npqfocaa6PXg2AiYgXp") : ((reg2368[(3'h7):(1'h1)] < reg2357[(3'h4):(3'h4)]) ?
              reg2385[(4'ha):(3'h4)] : ($signed(reg2400) ~^ wire2353))));
      reg2405 <= ({$unsigned($signed(forvar2366[(3'h6):(2'h3)])),
          reg2362[(2'h2):(1'h1)]} == reg2397);
      for (forvar2406 = (1'h0); (forvar2406 < (3'h5)); forvar2406 = (forvar2406 + (1'h1)))
        begin
          reg2407 <= reg2385[(4'h8):(3'h5)];
          reg2408 <= (^~(wire2351[(5'h15):(4'hf)] - (8'ha4)));
          reg2409 = wire2352;
          reg2410 = {$signed((^~$unsigned((reg2397 ~^ forvar2392))))};
          reg2411 <= forvar2390[(3'h5):(3'h5)];
          reg2412 <= $unsigned(((~^($unsigned(reg2391) ?
              (reg2356 ?
                  reg2367 : reg2363) : $unsigned(reg2367))) & $unsigned(reg2385[(1'h1):(1'h0)])));
        end
      for (forvar2413 = (1'h0); (forvar2413 < (3'h5)); forvar2413 = (forvar2413 + (1'h1)))
        begin
          reg2414 <= reg2358;
          reg2415 <= reg2409[(2'h2):(1'h0)];
          reg2416 <= reg2375[(2'h2):(1'h0)];
          reg2417 <= ($signed({wire2352[(2'h3):(2'h2)]}) ? reg2414 : reg2360);
          reg2418 <= $unsigned(reg2379);
        end
      reg2419 = reg2395[(3'h7):(3'h5)];
    end
  assign wire2420 = reg2400[(4'h9):(1'h1)];
  assign wire2421 = ($signed($signed(("Bf1NEOhxSO" & $signed(reg2363)))) & $signed((~|("y7mpG06gnK1LY37Cp1Wy" ?
                        {wire2350} : "7mLLAlQmgdJhr9EOc6XC"))));
  always
    @(posedge clk) begin
      reg2422 = "sDHCKgDxnEgXyTKnxws7TnB";
    end
  always
    @(posedge clk) begin
      reg2423 <= reg2414;
      for (forvar2424 = (1'h0); (forvar2424 < (1'h1)); forvar2424 = (forvar2424 + (1'h1)))
        begin
          reg2425 <= (-(reg2417 ?
              ((+reg2384) ?
                  reg2402[(2'h3):(1'h1)] : $unsigned($signed(forvar2390))) : $unsigned((reg2368 ^~ $signed(reg2376)))));
          reg2426 <= reg2403;
          reg2427 = (^reg2400);
        end
      reg2428 <= "ZAE1K7bH5oe34";
      for (forvar2429 = (1'h0); (forvar2429 < (3'h5)); forvar2429 = (forvar2429 + (1'h1)))
        begin
          reg2430 <= $signed({$unsigned($unsigned((-reg2426))),
              {(-forvar2373[(4'ha):(3'h4)])}});
          reg2431 <= ((~|reg2402) ?
              (~&reg2408) : ((-reg2398) + $signed(reg2427)));
        end
    end
  always
    @(posedge clk) begin
      for (forvar2432 = (1'h0); (forvar2432 < (1'h1)); forvar2432 = (forvar2432 + (1'h1)))
        begin
          reg2433 <= "SF3l0bHRwwP98hHY5i1rBld";
          if ((reg2402 ^ ""))
            begin
              reg2434 <= (((~|wire2350[(4'hf):(4'ha)]) ?
                  (reg2391[(3'h6):(3'h5)] ?
                      "SwQgSox53nkpAysEmmWdH" : forvar2429) : {(&reg2417[(4'h8):(4'h8)]),
                      ((-(8'ha6)) ?
                          $signed(reg2401) : $signed(reg2371))}) | $signed(wire2421[(4'ha):(1'h0)]));
              reg2435 = ($unsigned((reg2384[(1'h1):(1'h0)] + (|$unsigned(reg2386)))) ?
                  ((^~(~|(!reg2387))) < (&$unsigned(reg2374))) : reg2417);
            end
          else
            begin
              reg2434 <= "KRwx";
              reg2435 <= forvar2378;
              reg2436 <= (reg2368 ?
                  (7'h42) : (reg2409 + ((forvar2406[(2'h3):(1'h0)] + "7w6oiZYSCdCVII8p3q6") ?
                      $signed({reg2422, (8'hbb)}) : "Wt")));
            end
          for (forvar2437 = (1'h0); (forvar2437 < (1'h0)); forvar2437 = (forvar2437 + (1'h1)))
            begin
              reg2438 <= $signed($signed((~((reg2361 >> reg2393) > (&reg2409)))));
              reg2439 <= (^(reg2414 ?
                  $unsigned(reg2375[(1'h1):(1'h1)]) : (("YYm2CPbt3UiYZlN9hOS" != (reg2403 ?
                      reg2385 : reg2397)) * ((~|reg2411) ?
                      {reg2399} : (-forvar2437)))));
              reg2440 = $unsigned((~reg2427[(2'h2):(1'h1)]));
              reg2441 = reg2415[(3'h7):(3'h4)];
            end
          if (wire2350[(4'hc):(3'h5)])
            begin
              for (forvar2442 = (1'h0); (forvar2442 < (2'h3)); forvar2442 = (forvar2442 + (1'h1)))
                begin
                  reg2443 <= "95Zkltmr";
                  reg2444 <= (((~|"YF6TTqezMZc") ?
                          "dBwm" : $unsigned(reg2423[(3'h4):(3'h4)])) ?
                      "vezYdX1" : (reg2418 <<< "R8PKZVBdu4rohZD0"));
                  reg2445 <= "KKd5QPM5gozqwEfsqqs8ytBX";
                  reg2446 <= $signed(reg2418[(3'h7):(3'h5)]);
                  reg2447 <= (!$signed($signed(({reg2433, reg2402} ?
                      (reg2425 ?
                          reg2443 : (7'h41)) : reg2401[(1'h0):(1'h0)]))));
                  reg2448 <= $signed($unsigned((~$signed(reg2441[(1'h0):(1'h0)]))));
                end
              for (forvar2449 = (1'h0); (forvar2449 < (1'h0)); forvar2449 = (forvar2449 + (1'h1)))
                begin
                  reg2450 <= $signed("QNquMQG9");
                end
              for (forvar2451 = (1'h0); (forvar2451 < (2'h2)); forvar2451 = (forvar2451 + (1'h1)))
                begin
                  reg2452 = reg2419[(3'h6):(1'h1)];
                  reg2453 <= $signed(reg2403);
                  reg2454 <= reg2370[(5'h11):(3'h6)];
                  reg2455 = "";
                end
              for (forvar2456 = (1'h0); (forvar2456 < (3'h5)); forvar2456 = (forvar2456 + (1'h1)))
                begin
                  reg2457 <= wire2382[(4'hc):(2'h3)];
                  reg2458 <= (($signed(reg2374) ?
                      reg2419 : wire2420) ^~ ($unsigned(reg2408[(4'h9):(2'h2)]) | ($signed({forvar2388,
                          reg2457}) ?
                      $signed($unsigned(reg2365)) : (((8'hb9) ?
                              (8'h9f) : reg2412) ?
                          reg2453 : "7OhVFVe9r"))));
                end
              reg2459 <= reg2450;
            end
          else
            begin
              reg2442 <= reg2410[(3'h4):(1'h1)];
              reg2443 <= "SF0JJSHTPZuddu3pEU1Z4dRIs";
              reg2444 <= (^$signed(((reg2380 ?
                  $unsigned(reg2450) : forvar2354[(2'h2):(2'h2)]) ^ $signed($signed(forvar2373)))));
              reg2445 <= forvar2373[(2'h2):(1'h1)];
              reg2446 <= (reg2427 ?
                  "zcCdaFMIC" : (forvar2394 + ($signed((reg2363 > forvar2449)) ?
                      $signed($unsigned(wire2350)) : "TUnbqT")));
              reg2447 <= (((forvar2424 ?
                      reg2415[(3'h5):(3'h4)] : (^~(reg2375 ?
                          reg2396 : reg2402))) == reg2389) ?
                  $unsigned((!(8'hb3))) : $signed($unsigned(reg2383[(4'hc):(1'h0)])));
            end
          for (forvar2460 = (1'h0); (forvar2460 < (1'h0)); forvar2460 = (forvar2460 + (1'h1)))
            begin
              reg2461 <= ((8'hbf) ?
                  "JuD7TpZiM2rpisUsdEBSrc0" : ((~&"iVkH8XgTgp9A8") ?
                      (reg2395 ?
                          reg2409[(1'h1):(1'h0)] : {(reg2400 ?
                                  (8'hac) : (8'ha7))}) : {"PCQPZkokD"}));
              reg2462 = (8'hb6);
            end
          if ((reg2419 ?
              {(($signed((8'h9c)) ? $signed(reg2417) : {reg2400}) ?
                      reg2427[(1'h0):(1'h0)] : (!{(8'h9c), (8'hac)})),
                  $signed($unsigned($unsigned(forvar2378)))} : (+(forvar2378[(4'hf):(3'h4)] ?
                  $unsigned({reg2436}) : ((reg2381 ?
                      wire2353 : reg2425) > ((7'h41) <<< reg2427))))))
            begin
              reg2463 <= reg2370[(4'hd):(1'h0)];
              reg2464 = (^reg2380);
              for (forvar2465 = (1'h0); (forvar2465 < (1'h1)); forvar2465 = (forvar2465 + (1'h1)))
                begin
                  reg2466 <= (~|$unsigned((+((reg2461 <<< reg2426) ?
                      (reg2367 * reg2369) : (~^(8'hb7))))));
                  reg2467 <= ((^(~^((reg2414 | reg2457) >> $signed(reg2401)))) ?
                      wire2382[(3'h5):(3'h4)] : ({reg2415[(4'h8):(3'h5)],
                          (~|reg2375[(1'h1):(1'h1)])} ^~ {$unsigned((+reg2357)),
                          "N8"}));
                  reg2468 <= (&(reg2423 ? $unsigned("") : $signed(reg2434)));
                end
              reg2469 <= forvar2378;
            end
          else
            begin
              reg2463 <= ({reg2391,
                  forvar2456[(3'h7):(2'h2)]} << $signed($unsigned((-(wire2420 ?
                  reg2409 : reg2459)))));
            end
        end
      reg2470 = reg2425;
      reg2471 <= $signed("nJHJrkYr0pRHYBB9JkQ");
      reg2472 <= (("09TyWCZcAuM2YIbJ0lSBa" | forvar2388) >= ((~$unsigned((~^forvar2442))) ?
          wire2421 : $unsigned($unsigned((reg2440 ? reg2411 : reg2419)))));
      reg2473 <= (((|((~^(8'ha2)) >> (-reg2399))) <= ("XRtaEwL" + (&(^(7'h40))))) || ($signed({(forvar2456 ?
              reg2358 : forvar2432)}) <= $unsigned((8'h9c))));
    end
  always
    @(posedge clk) begin
      for (forvar2474 = (1'h0); (forvar2474 < (2'h3)); forvar2474 = (forvar2474 + (1'h1)))
        begin
          reg2475 = reg2355[(2'h2):(1'h1)];
          reg2476 = reg2415[(1'h1):(1'h1)];
          reg2477 <= ("" ? reg2408[(4'hc):(3'h4)] : "");
        end
      reg2478 = $unsigned((~^$signed((7'h43))));
      reg2479 <= "6ewUOLb";
      reg2480 <= {$unsigned((&reg2402))};
      reg2481 = (^~((~|(^$signed(forvar2366))) * (($unsigned(reg2415) <= {reg2367,
              reg2455}) ?
          $signed(reg2385) : ((reg2410 << reg2412) <= (reg2466 ?
              reg2371 : reg2374)))));
    end
  always
    @(posedge clk) begin
      for (forvar2482 = (1'h0); (forvar2482 < (2'h2)); forvar2482 = (forvar2482 + (1'h1)))
        begin
          reg2483 = {$unsigned(reg2422[(1'h1):(1'h1)])};
          reg2484 <= (7'h4b);
          reg2485 <= (~|(((~((8'hac) && reg2379)) && reg2362) >>> (^~reg2427)));
        end
      reg2486 <= (reg2407[(3'h5):(3'h5)] ?
          $signed(reg2434) : wire2420[(5'h14):(5'h14)]);
      reg2487 <= (^(~^(~&(reg2462[(4'h9):(3'h7)] ~^ (forvar2429 != reg2393)))));
    end
  always
    @(posedge clk) begin
      reg2488 = reg2459[(2'h3):(1'h0)];
      reg2489 <= "Ja4SsY2C";
    end
  always
    @(posedge clk) begin
      reg2490 <= ("wBOckq92PuZyVsR" ?
          (+forvar2390[(3'h4):(2'h3)]) : {reg2405[(3'h4):(1'h1)],
              ((wire2353[(3'h5):(2'h3)] ^ (reg2463 * reg2376)) != $signed(reg2455))});
      reg2491 <= reg2398[(4'he):(4'ha)];
      reg2492 = reg2369;
      reg2493 <= "DAfM57Q1N8U3L";
      reg2494 <= (reg2401 ?
          (!((-forvar2372) ?
              $signed(reg2463) : reg2443[(3'h4):(3'h4)])) : $unsigned(reg2447));
      reg2495 <= ((8'h9f) ?
          ("rx0FB77qQxAmB8svnKTWnB" ?
              $unsigned(forvar2429[(2'h2):(1'h0)]) : "Z") : ("x99Ku6neSrCTe" < (&(~(~reg2400)))));
    end
  assign wire2496 = (~&reg2371[(2'h2):(1'h1)]);
  always
    @(posedge clk) begin
      reg2497 <= $signed({(reg2371[(2'h3):(1'h1)] ?
              reg2387[(4'ha):(3'h7)] : (reg2446[(3'h6):(3'h4)] ?
                  ((8'hbf) ^ reg2354) : "S")),
          reg2399});
    end
  always
    @(posedge clk) begin
      reg2498 <= ($unsigned($signed(("h" + reg2430[(3'h4):(1'h1)]))) ?
          $signed((|$signed((reg2457 ?
              reg2479 : reg2374)))) : ($signed(("JPTufdUq7LMlF7sc0HTEywh8h" ?
              reg2375 : reg2383[(4'ha):(1'h1)])) - (reg2360 || ($signed(reg2389) ?
              ((7'h41) >>> reg2472) : reg2381))));
      for (forvar2499 = (1'h0); (forvar2499 < (3'h4)); forvar2499 = (forvar2499 + (1'h1)))
        begin
          reg2500 <= (~^reg2414);
          for (forvar2501 = (1'h0); (forvar2501 < (3'h5)); forvar2501 = (forvar2501 + (1'h1)))
            begin
              if (($unsigned("cLuWbUIWhalfXWLpTXgOW4") ?
                  $unsigned((8'ha2)) : ($unsigned((+(forvar2424 ?
                      reg2452 : (8'haf)))) ~^ forvar2474)))
                begin
                  reg2502 <= (|"TWriu3UKZ");
                  reg2503 <= reg2377[(2'h2):(1'h0)];
                end
              else
                begin
                  reg2502 <= (reg2453 ? reg2468[(2'h2):(1'h1)] : forvar2373);
                  reg2503 <= {($signed((^~$unsigned(reg2461))) ?
                          "FKiDFVu" : (("qn2e4gsSkx" ?
                              (~|reg2462) : $unsigned(reg2398)) ^~ "aq8n"))};
                  reg2504 <= "J7JGw0TpnpbQD";
                  reg2505 <= (^~$signed("bzp"));
                  reg2506 <= "6YSI243KF3aLbPtqaRU";
                  reg2507 = reg2438[(5'h12):(1'h1)];
                end
            end
          reg2508 = $unsigned(forvar2460[(3'h6):(3'h4)]);
          reg2509 = $signed($signed({(-$unsigned(reg2386)),
              (^~(reg2466 ? (8'hbd) : reg2409))}));
          for (forvar2510 = (1'h0); (forvar2510 < (2'h3)); forvar2510 = (forvar2510 + (1'h1)))
            begin
              reg2511 = {{{((reg2495 ? (7'h4d) : forvar2501) ?
                              (^~reg2498) : "KuXEaT5MaNO2Bf")}}};
              reg2512 <= $unsigned(reg2356[(5'h11):(4'h8)]);
              reg2513 <= $unsigned("i");
              for (forvar2514 = (1'h0); (forvar2514 < (2'h3)); forvar2514 = (forvar2514 + (1'h1)))
                begin
                  reg2515 <= $unsigned($signed($signed($unsigned($signed(reg2439)))));
                  reg2516 <= ($unsigned(("bdqcBx" ?
                      forvar2406 : ($signed(forvar2372) ?
                          $signed(reg2397) : (reg2458 ?
                              forvar2390 : forvar2392)))) ^~ reg2358);
                  reg2517 = reg2452;
                  reg2518 <= $unsigned(forvar2451);
                  reg2519 <= (|((reg2439[(4'hb):(4'h8)] * ($signed((8'hbb)) ?
                          reg2355[(4'hd):(4'hd)] : (reg2491 ?
                              forvar2437 : wire2352))) ?
                      "DpCru9BhF7edBVTuqBo2" : $signed(reg2397[(3'h5):(3'h4)])));
                  reg2520 <= (({"xJ0bOANmM1fZb4",
                          $signed((reg2412 <= reg2399))} * reg2507[(2'h2):(2'h2)]) ?
                      $signed($unsigned(("URKwMwsKw" ?
                          (-reg2493) : (8'hb6)))) : (((^$signed(reg2485)) ?
                              (reg2384[(2'h2):(1'h1)] ?
                                  (|reg2422) : $signed(reg2389)) : (8'hb0)) ?
                          (($signed((8'ha5)) ?
                              ((8'haa) ?
                                  forvar2392 : reg2511) : $unsigned(reg2517)) && $signed(forvar2482)) : reg2507[(4'hc):(4'h8)]));
                end
            end
        end
      reg2521 <= (reg2473 ~^ $signed((("SySC7" << reg2488) ?
          "t7ycV8" : (reg2511[(3'h6):(3'h6)] ?
              {(8'ha3)} : {reg2385, reg2515}))));
      reg2522 <= reg2391;
      for (forvar2523 = (1'h0); (forvar2523 < (1'h0)); forvar2523 = (forvar2523 + (1'h1)))
        begin
          for (forvar2524 = (1'h0); (forvar2524 < (3'h4)); forvar2524 = (forvar2524 + (1'h1)))
            begin
              reg2525 = (reg2385[(3'h7):(2'h2)] ?
                  (&($unsigned($signed(reg2466)) << reg2491[(4'h9):(1'h1)])) : reg2393);
              reg2526 <= $unsigned("zZDt27KRYdAKvQBUYFtx");
              reg2527 <= reg2486;
              reg2528 <= "y2uSml1Exg2ewQJZhhMODqS";
            end
          reg2529 <= ("zzGoMbSMFUv4Cf4xwizkmy" ?
              reg2443 : $unsigned((("uXr" ?
                  $signed(reg2517) : (~&forvar2372)) == $unsigned(reg2407[(3'h4):(2'h2)]))));
          reg2530 = reg2433;
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2298  (y, clk, wire2302, wire2301, wire2300, wire2299);
  output wire [(32'h277):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire2302;
  input wire [(3'h4):(1'h0)] wire2301;
  input wire [(5'h13):(1'h0)] wire2300;
  input wire signed [(5'h18):(1'h0)] wire2299;
  wire [(2'h3):(1'h0)] wire2346;
  reg [(4'ha):(1'h0)] reg2345 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2344 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2343 = (1'h0);
  reg [(3'h5):(1'h0)] reg2342 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2341 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2340 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2339 = (1'h0);
  reg [(5'h14):(1'h0)] reg2338 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2337 = (1'h0);
  reg [(4'he):(1'h0)] reg2336 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2335 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2334 = (1'h0);
  reg [(5'h11):(1'h0)] reg2333 = (1'h0);
  reg [(4'h9):(1'h0)] reg2332 = (1'h0);
  reg [(4'he):(1'h0)] reg2331 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2328 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2330 = (1'h0);
  reg [(3'h6):(1'h0)] reg2329 = (1'h0);
  reg [(4'hf):(1'h0)] reg2328 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2327 = (1'h0);
  reg [(4'hc):(1'h0)] reg2326 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2325 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2324 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2323 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2322 = (1'h0);
  reg [(3'h4):(1'h0)] reg2321 = (1'h0);
  reg [(5'h17):(1'h0)] reg2320 = (1'h0);
  reg [(3'h4):(1'h0)] reg2319 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2318 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar2317 = (1'h0);
  wire [(5'h19):(1'h0)] wire2316;
  reg signed [(5'h1a):(1'h0)] reg2315 = (1'h0);
  reg [(4'hb):(1'h0)] reg2314 = (1'h0);
  reg [(4'h8):(1'h0)] reg2313 = (1'h0);
  wire [(4'hc):(1'h0)] wire2312;
  reg [(2'h2):(1'h0)] reg2311 = (1'h0);
  reg [(5'h10):(1'h0)] reg2310 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2309 = (1'h0);
  reg [(5'h17):(1'h0)] reg2308 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2307 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2306 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2305 = (1'h0);
  reg [(3'h7):(1'h0)] reg2304 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2303 = (1'h0);
  assign y = {wire2346,
                 reg2345,
                 reg2344,
                 reg2343,
                 reg2342,
                 forvar2341,
                 reg2340,
                 reg2339,
                 reg2338,
                 reg2337,
                 reg2336,
                 reg2335,
                 forvar2334,
                 reg2333,
                 reg2332,
                 reg2331,
                 forvar2328,
                 reg2330,
                 reg2329,
                 reg2328,
                 reg2327,
                 reg2326,
                 reg2325,
                 reg2324,
                 reg2323,
                 reg2322,
                 reg2321,
                 reg2320,
                 reg2319,
                 forvar2318,
                 forvar2317,
                 wire2316,
                 reg2315,
                 reg2314,
                 reg2313,
                 wire2312,
                 reg2311,
                 reg2310,
                 reg2309,
                 reg2308,
                 reg2307,
                 reg2306,
                 reg2305,
                 reg2304,
                 forvar2303,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar2303 = (1'h0); (forvar2303 < (2'h3)); forvar2303 = (forvar2303 + (1'h1)))
        begin
          reg2304 <= (!("vdAAmooAIndL0W9pzLb" ?
              forvar2303 : (((8'ha5) * (~|wire2299)) ?
                  $unsigned($signed(wire2299)) : (!"IJTGpzlyWaP8o"))));
          reg2305 <= ($unsigned((&((wire2302 ? wire2301 : forvar2303) ?
              reg2304 : $signed(wire2299)))) < ($signed(((wire2302 ?
              wire2302 : wire2300) | wire2301)) | wire2299[(5'h16):(1'h1)]));
          reg2306 <= (~(8'hb9));
          reg2307 <= (~(!"YkJNrRZ9lw46GDGnthQd"));
          reg2308 <= (^reg2304);
        end
      reg2309 = ({reg2308} != reg2307[(1'h1):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg2310 <= "tTLz1ybV6a9vhm";
      reg2311 = forvar2303;
    end
  assign wire2312 = "9tW9cxrU3";
  always
    @(posedge clk) begin
      reg2313 = (^($signed($unsigned(wire2312[(4'ha):(4'ha)])) ?
          (~|"D1CRkxJZOhCg3uFe9") : (("YEFR3eXyLuJ" ?
                  (wire2312 ? wire2302 : wire2300) : $signed(reg2311)) ?
              (~(wire2300 ?
                  wire2300 : reg2310)) : $unsigned($signed((7'h46))))));
      reg2314 <= reg2313[(2'h3):(1'h1)];
      reg2315 = (reg2305[(2'h3):(2'h2)] ?
          $signed($signed($signed("wVZrynN8g80NfpolJpTTLGNf"))) : wire2299);
    end
  assign wire2316 = {"JIZhwKsm6m7JlAos", "oHU"};
  always
    @(posedge clk) begin
      for (forvar2317 = (1'h0); (forvar2317 < (2'h3)); forvar2317 = (forvar2317 + (1'h1)))
        begin
          for (forvar2318 = (1'h0); (forvar2318 < (1'h0)); forvar2318 = (forvar2318 + (1'h1)))
            begin
              reg2319 <= $signed({({wire2302, $signed(forvar2317)} ?
                      "y8zSC9zry7N5Q9yC6k" : (&{reg2313, wire2312})),
                  $unsigned($unsigned((|(8'ha8))))});
              reg2320 = (reg2305 ?
                  $unsigned((|(+$unsigned((8'ha2))))) : $signed((-($signed(wire2299) - "kCmOrRq8DGKcAPMXsElIcWcE"))));
              reg2321 <= reg2308;
              reg2322 <= "WpazwnkRl";
              reg2323 <= $signed(wire2301);
            end
          reg2324 <= reg2319[(1'h0):(1'h0)];
        end
      if (reg2307[(3'h4):(2'h2)])
        begin
          reg2325 = wire2302[(4'ha):(2'h3)];
          reg2326 <= "Bq";
          reg2327 <= ((+(~&$unsigned($signed(reg2324)))) ?
              $unsigned("OqpwKUcqBuT") : reg2310[(4'he):(1'h0)]);
          reg2328 = $unsigned(("TS7mO7694" == $signed($signed(reg2322[(2'h2):(2'h2)]))));
          reg2329 <= $signed({{wire2299}, $signed(wire2312[(4'hb):(2'h2)])});
          reg2330 <= $unsigned("gN");
        end
      else
        begin
          reg2325 <= reg2327[(5'h19):(4'hb)];
          reg2326 <= ({($signed("kUV2") ?
                      ("WgqmV" ?
                          (forvar2303 ?
                              reg2307 : forvar2318) : "NlWyNHB") : $unsigned((wire2299 ?
                          reg2323 : wire2316)))} ?
              (reg2325[(5'h10):(4'hb)] ~^ ({"lPAHxqNUHAERBtecAt8Wvuhrw",
                      reg2307} ?
                  "6pU2q0ue4FQ" : (~^(~&reg2309)))) : $signed({$signed("GLdlVOZYWWMhIBlHBd"),
                  "sfDlnr08iXbYFw"}));
          reg2327 <= $signed((&"Fw1Rwi5O2qmHIIB9OL6fV"));
          for (forvar2328 = (1'h0); (forvar2328 < (2'h2)); forvar2328 = (forvar2328 + (1'h1)))
            begin
              reg2329 <= wire2316[(1'h0):(1'h0)];
              reg2330 <= {reg2321[(1'h1):(1'h1)],
                  $unsigned(((~^$unsigned(reg2323)) >> ((reg2307 ?
                      reg2305 : wire2300) ^ "14q0uIJB4c")))};
              reg2331 <= wire2316;
            end
          reg2332 <= reg2304[(1'h1):(1'h1)];
        end
      reg2333 <= ($unsigned($unsigned("4oe0lORhlXHxysf")) ?
          "qrvIDMKbxbO5B1C08NF8gEXe" : {"Tw1Al",
              (&{reg2329[(2'h3):(2'h2)], (7'h48)})});
    end
  always
    @(posedge clk) begin
      for (forvar2334 = (1'h0); (forvar2334 < (3'h4)); forvar2334 = (forvar2334 + (1'h1)))
        begin
          reg2335 = "HFuJo0";
          reg2336 = $signed(forvar2317[(4'hb):(3'h4)]);
        end
      reg2337 = $signed(wire2301[(1'h0):(1'h0)]);
      reg2338 <= (-($unsigned($unsigned(reg2331[(4'hb):(2'h3)])) ?
          {((reg2308 ? reg2329 : reg2309) * forvar2334),
              reg2331[(2'h3):(1'h0)]} : reg2323));
    end
  always
    @(posedge clk) begin
      reg2339 = $signed("eYLfQcEsOS");
      reg2340 <= ($unsigned($unsigned($unsigned("GS436YO5"))) >>> (8'haf));
      for (forvar2341 = (1'h0); (forvar2341 < (1'h0)); forvar2341 = (forvar2341 + (1'h1)))
        begin
          reg2342 <= (reg2321[(1'h1):(1'h1)] ?
              "cgkUC" : (forvar2303 ? {"mXUcG", reg2330} : reg2326));
        end
    end
  always
    @(posedge clk) begin
      reg2343 = $unsigned($unsigned($signed(reg2310)));
      reg2344 = $unsigned(reg2332[(3'h4):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg2345 <= ("yaRz50SYIDS" ?
          $signed((~$signed($unsigned((8'hac))))) : "4h6AeyL0XyoZ");
    end
  assign wire2346 = (~"sUJbs9");
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2227
#( parameter param2278 = (!(~&((((8'ha2) << (7'h41)) - ((8'hb8) <= (8'ha6))) << {{(8'h9f)}, ((8'hba) >= (7'h42))})))
, parameter param2279 = (^param2278) )
(y, clk, wire2231, wire2230, wire2229, wire2228);
  output wire [(32'h291):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire2231;
  input wire signed [(3'h4):(1'h0)] wire2230;
  input wire [(4'hc):(1'h0)] wire2229;
  input wire signed [(3'h6):(1'h0)] wire2228;
  wire [(5'h17):(1'h0)] wire2277;
  reg signed [(5'h11):(1'h0)] reg2276 = (1'h0);
  reg [(4'he):(1'h0)] reg2275 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2274 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2273 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2272 = (1'h0);
  reg [(4'h8):(1'h0)] reg2271 = (1'h0);
  reg [(4'hc):(1'h0)] reg2270 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2269 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2268 = (1'h0);
  reg [(5'h12):(1'h0)] forvar2267 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2266 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2265 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2264 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2263 = (1'h0);
  reg [(3'h5):(1'h0)] reg2262 = (1'h0);
  reg [(2'h2):(1'h0)] reg2261 = (1'h0);
  reg [(5'h17):(1'h0)] reg2260 = (1'h0);
  reg [(4'h8):(1'h0)] reg2259 = (1'h0);
  reg [(5'h14):(1'h0)] reg2258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2257 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2256 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2255 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2254 = (1'h0);
  reg [(4'hd):(1'h0)] reg2253 = (1'h0);
  reg [(4'ha):(1'h0)] reg2252 = (1'h0);
  reg [(2'h3):(1'h0)] reg2251 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2250 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2249 = (1'h0);
  reg [(5'h11):(1'h0)] reg2248 = (1'h0);
  reg [(4'hb):(1'h0)] reg2247 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2246 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2245 = (1'h0);
  reg [(3'h7):(1'h0)] reg2244 = (1'h0);
  reg [(5'h10):(1'h0)] reg2243 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2240 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2238 = (1'h0);
  reg [(5'h15):(1'h0)] reg2242 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2241 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2240 = (1'h0);
  reg [(5'h14):(1'h0)] reg2239 = (1'h0);
  reg [(5'h15):(1'h0)] reg2238 = (1'h0);
  reg [(3'h4):(1'h0)] reg2237 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2236 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2235 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2234 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2233 = (1'h0);
  wire [(5'h13):(1'h0)] wire2232;
  assign y = {wire2277,
                 reg2276,
                 reg2275,
                 reg2274,
                 forvar2273,
                 reg2272,
                 reg2271,
                 reg2270,
                 reg2269,
                 reg2268,
                 forvar2267,
                 forvar2266,
                 reg2265,
                 forvar2264,
                 reg2263,
                 reg2262,
                 reg2261,
                 reg2260,
                 reg2259,
                 reg2258,
                 reg2257,
                 reg2256,
                 reg2255,
                 reg2254,
                 reg2253,
                 reg2252,
                 reg2251,
                 reg2250,
                 reg2249,
                 reg2248,
                 reg2247,
                 reg2246,
                 forvar2245,
                 reg2244,
                 reg2243,
                 reg2240,
                 forvar2238,
                 reg2242,
                 reg2241,
                 forvar2240,
                 reg2239,
                 reg2238,
                 reg2237,
                 reg2236,
                 forvar2235,
                 reg2234,
                 reg2233,
                 wire2232,
                 (1'h0)};
  assign wire2232 = $signed(($unsigned("lO4mJDZGaCB") ^ $signed("PAWu6")));
  always
    @(posedge clk) begin
      reg2233 <= $signed($signed($unsigned(((wire2228 ? (8'hb2) : (8'ha4)) ?
          (8'had) : (wire2231 > wire2231)))));
      reg2234 = $unsigned("B9r0BP4zQVV5ltN");
      for (forvar2235 = (1'h0); (forvar2235 < (2'h3)); forvar2235 = (forvar2235 + (1'h1)))
        begin
          if ({"Ge8O8kzJaqDyuySqPfPLgHfS2"})
            begin
              reg2236 <= (("wi" ?
                  forvar2235 : wire2230) << (reg2233[(5'h16):(4'hb)] ?
                  reg2234[(3'h5):(3'h4)] : wire2228));
              reg2237 = {(~^wire2231[(4'hb):(3'h4)])};
              reg2238 = ((wire2230 || wire2232) | reg2234);
              reg2239 = wire2229;
              for (forvar2240 = (1'h0); (forvar2240 < (3'h5)); forvar2240 = (forvar2240 + (1'h1)))
                begin
                  reg2241 <= "oK8q4u94v83Pq";
                  reg2242 <= $signed(((reg2236 ~^ ("p5HNw" ?
                      $signed(wire2230) : (reg2237 ?
                          wire2231 : reg2234))) == forvar2235[(1'h1):(1'h1)]));
                end
            end
          else
            begin
              reg2236 = (forvar2240 ? reg2237 : (-(&"eprcgdPSwKXg")));
              reg2237 <= reg2236[(2'h2):(2'h2)];
              for (forvar2238 = (1'h0); (forvar2238 < (3'h4)); forvar2238 = (forvar2238 + (1'h1)))
                begin
                  reg2239 <= "eSZIOeZPXVKEtlyYr7b7NOp";
                  reg2240 <= $signed(reg2238[(4'h9):(1'h0)]);
                  reg2241 <= wire2228[(2'h2):(2'h2)];
                  reg2242 <= (~{reg2241[(4'h8):(2'h2)], forvar2238});
                  reg2243 <= (wire2229[(1'h1):(1'h0)] ?
                      "Fvx4dvrq7" : {forvar2238, forvar2235[(2'h2):(1'h1)]});
                  reg2244 = (^~($signed(wire2232[(5'h11):(2'h3)]) ~^ forvar2240[(1'h1):(1'h1)]));
                end
              for (forvar2245 = (1'h0); (forvar2245 < (2'h2)); forvar2245 = (forvar2245 + (1'h1)))
                begin
                  reg2246 <= forvar2240;
                  reg2247 <= $signed(((reg2242 >= "3ZstIeEdRUUOuVT7bPaRE") < reg2236));
                  reg2248 <= $signed((^(~|$signed("zEP5"))));
                  reg2249 <= forvar2245[(1'h0):(1'h0)];
                  reg2250 <= {"v"};
                end
              if ((~(($unsigned((~|wire2231)) || (~reg2241)) ?
                  (7'h47) : ((^forvar2235) || reg2246))))
                begin
                  reg2251 <= reg2248;
                  reg2252 <= $unsigned((~&"eHgcGsVNMS5x"));
                end
              else
                begin
                  reg2251 <= (({$signed((reg2243 * forvar2240)),
                          $signed($signed((7'h49)))} && $unsigned((8'h9e))) ?
                      reg2247[(4'hb):(1'h1)] : $signed(wire2230[(1'h0):(1'h0)]));
                end
            end
          reg2253 = "2LczL8IZGb9oPM3Ori0";
        end
      reg2254 <= $signed($signed(reg2236[(5'h18):(4'h9)]));
      reg2255 <= reg2254[(4'h9):(4'h9)];
      reg2256 <= reg2233;
    end
  always
    @(posedge clk) begin
      reg2257 <= $signed("7APoJlwUVs");
      reg2258 <= (8'haa);
      reg2259 = {wire2232};
      reg2260 <= (reg2252 & reg2254);
      reg2261 <= $unsigned($signed(reg2255[(4'hb):(4'h8)]));
    end
  always
    @(posedge clk) begin
      reg2262 <= "cMIhFavu5vvnYqMQiPgVr4mf";
      reg2263 = (7'h49);
      for (forvar2264 = (1'h0); (forvar2264 < (1'h0)); forvar2264 = (forvar2264 + (1'h1)))
        begin
          reg2265 <= (reg2258[(5'h14):(4'ha)] * $signed($signed(reg2263[(4'hf):(3'h4)])));
        end
      for (forvar2266 = (1'h0); (forvar2266 < (2'h2)); forvar2266 = (forvar2266 + (1'h1)))
        begin
          for (forvar2267 = (1'h0); (forvar2267 < (3'h5)); forvar2267 = (forvar2267 + (1'h1)))
            begin
              reg2268 <= (("5ZgPDAvT1rNNmDIF86g" >= (($signed((8'haf)) + "eyF") ^ $signed({reg2262,
                  (8'hb6)}))) ^ wire2229);
              reg2269 = ("wRGHlw" ?
                  reg2250[(3'h5):(1'h1)] : $unsigned((+wire2232[(5'h10):(4'hb)])));
              reg2270 <= ($signed($signed(forvar2266[(3'h5):(1'h1)])) >> $unsigned((^$unsigned($unsigned((8'hab))))));
              reg2271 <= (~^reg2250[(1'h0):(1'h0)]);
              reg2272 <= wire2230[(2'h2):(1'h0)];
            end
        end
      for (forvar2273 = (1'h0); (forvar2273 < (2'h2)); forvar2273 = (forvar2273 + (1'h1)))
        begin
          reg2274 <= forvar2238[(3'h4):(1'h1)];
          reg2275 <= "bMIkQedDq";
        end
    end
  always
    @(posedge clk) begin
      reg2276 <= ($signed((~|forvar2238[(1'h0):(1'h0)])) ?
          {"OI10fM4zWrKfip35L8h",
              (^~$unsigned({reg2256}))} : reg2236[(1'h0):(1'h0)]);
    end
  assign wire2277 = ("JHLXHumRFgShqm7xuFUvBbeuo" <= reg2261);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2112
#( parameter param2224 = {(^({((7'h44) > (8'hb2)), ((8'hbf) ? (7'h46) : (8'ha6))} ? (8'hb7) : {(~|(8'hb5))})), ((^(((8'ha8) ? (8'hab) : (8'hb7)) ? ((7'h4e) ? (8'hb4) : (7'h43)) : (~(7'h40)))) >>> {((&(8'hb3)) ? {(8'haf)} : (~|(8'haf)))})} )
(y, clk, wire2116, wire2115, wire2114, wire2113);
  output wire [(32'h5ae):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire2116;
  input wire [(5'h14):(1'h0)] wire2115;
  input wire signed [(2'h2):(1'h0)] wire2114;
  input wire signed [(4'hf):(1'h0)] wire2113;
  reg signed [(4'hb):(1'h0)] reg2223 = (1'h0);
  reg [(5'h10):(1'h0)] reg2222 = (1'h0);
  reg [(2'h2):(1'h0)] reg2221 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2220 = (1'h0);
  reg [(5'h11):(1'h0)] forvar2219 = (1'h0);
  reg [(3'h5):(1'h0)] reg2218 = (1'h0);
  reg [(5'h1a):(1'h0)] reg2217 = (1'h0);
  reg [(5'h15):(1'h0)] reg2216 = (1'h0);
  reg [(5'h15):(1'h0)] reg2215 = (1'h0);
  reg [(4'he):(1'h0)] reg2214 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2213 = (1'h0);
  reg [(4'he):(1'h0)] forvar2212 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar2211 = (1'h0);
  reg [(5'h11):(1'h0)] reg2210 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2209 = (1'h0);
  reg [(4'h8):(1'h0)] reg2208 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire2207;
  wire signed [(4'hc):(1'h0)] wire2206;
  wire [(5'h13):(1'h0)] wire2205;
  reg signed [(3'h4):(1'h0)] reg2204 = (1'h0);
  reg [(4'hf):(1'h0)] reg2203 = (1'h0);
  reg [(5'h16):(1'h0)] reg2202 = (1'h0);
  reg [(4'ha):(1'h0)] reg2201 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2200 = (1'h0);
  reg [(3'h5):(1'h0)] reg2199 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2198 = (1'h0);
  reg [(5'h11):(1'h0)] reg2197 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire2196;
  wire [(3'h4):(1'h0)] wire2195;
  wire [(4'h9):(1'h0)] wire2194;
  reg [(4'hb):(1'h0)] reg2193 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2192 = (1'h0);
  reg [(4'hf):(1'h0)] reg2191 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2190 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2189 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2188 = (1'h0);
  reg [(3'h4):(1'h0)] reg2187 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2186 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2185 = (1'h0);
  reg [(4'h9):(1'h0)] reg2184 = (1'h0);
  reg [(2'h2):(1'h0)] reg2183 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2182 = (1'h0);
  reg [(5'h12):(1'h0)] reg2181 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2180 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2179 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg2178 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire2177;
  reg [(5'h19):(1'h0)] reg2176 = (1'h0);
  reg [(5'h10):(1'h0)] reg2175 = (1'h0);
  reg [(3'h7):(1'h0)] reg2174 = (1'h0);
  reg [(5'h19):(1'h0)] reg2173 = (1'h0);
  wire signed [(5'h17):(1'h0)] wire2172;
  reg [(4'h9):(1'h0)] reg2171 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar2170 = (1'h0);
  reg [(3'h6):(1'h0)] reg2169 = (1'h0);
  reg [(5'h14):(1'h0)] reg2168 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2167 = (1'h0);
  reg [(3'h7):(1'h0)] reg2166 = (1'h0);
  reg [(4'hd):(1'h0)] reg2165 = (1'h0);
  reg [(3'h7):(1'h0)] reg2164 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2163 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2162 = (1'h0);
  reg [(5'h13):(1'h0)] reg2161 = (1'h0);
  reg [(4'h9):(1'h0)] reg2160 = (1'h0);
  reg [(5'h11):(1'h0)] reg2159 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2158 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2157 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2156 = (1'h0);
  wire [(4'hc):(1'h0)] wire2155;
  reg signed [(5'h11):(1'h0)] reg2154 = (1'h0);
  reg [(5'h14):(1'h0)] reg2153 = (1'h0);
  reg [(2'h2):(1'h0)] reg2152 = (1'h0);
  reg [(5'h19):(1'h0)] reg2151 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2150 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2149 = (1'h0);
  reg [(5'h15):(1'h0)] reg2148 = (1'h0);
  reg [(4'hc):(1'h0)] reg2147 = (1'h0);
  reg [(4'hb):(1'h0)] reg2146 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2145 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2144 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2143 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2142 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2141 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2140 = (1'h0);
  reg [(5'h15):(1'h0)] reg2139 = (1'h0);
  reg [(4'hb):(1'h0)] reg2138 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2137 = (1'h0);
  reg [(5'h14):(1'h0)] reg2136 = (1'h0);
  reg [(4'he):(1'h0)] forvar2135 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2134 = (1'h0);
  reg [(5'h11):(1'h0)] reg2133 = (1'h0);
  reg [(2'h2):(1'h0)] reg2132 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2131 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2130 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2129 = (1'h0);
  reg [(2'h2):(1'h0)] reg2128 = (1'h0);
  reg [(5'h13):(1'h0)] reg2127 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2126 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2125 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2124 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2123 = (1'h0);
  reg [(5'h18):(1'h0)] reg2122 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2121 = (1'h0);
  reg [(5'h11):(1'h0)] reg2120 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2119 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar2118 = (1'h0);
  reg [(4'he):(1'h0)] forvar2117 = (1'h0);
  assign y = {reg2223,
                 reg2222,
                 reg2221,
                 forvar2220,
                 forvar2219,
                 reg2218,
                 reg2217,
                 reg2216,
                 reg2215,
                 reg2214,
                 reg2213,
                 forvar2212,
                 forvar2211,
                 reg2210,
                 forvar2209,
                 reg2208,
                 wire2207,
                 wire2206,
                 wire2205,
                 reg2204,
                 reg2203,
                 reg2202,
                 reg2201,
                 reg2200,
                 reg2199,
                 reg2198,
                 reg2197,
                 wire2196,
                 wire2195,
                 wire2194,
                 reg2193,
                 reg2192,
                 reg2191,
                 reg2190,
                 forvar2189,
                 reg2188,
                 reg2187,
                 reg2186,
                 forvar2185,
                 reg2184,
                 reg2183,
                 reg2182,
                 reg2181,
                 reg2180,
                 reg2179,
                 reg2178,
                 wire2177,
                 reg2176,
                 reg2175,
                 reg2174,
                 reg2173,
                 wire2172,
                 reg2171,
                 forvar2170,
                 reg2169,
                 reg2168,
                 reg2167,
                 reg2166,
                 reg2165,
                 reg2164,
                 reg2163,
                 reg2162,
                 reg2161,
                 reg2160,
                 reg2159,
                 reg2158,
                 reg2157,
                 reg2156,
                 wire2155,
                 reg2154,
                 reg2153,
                 reg2152,
                 reg2151,
                 reg2150,
                 reg2149,
                 reg2148,
                 reg2147,
                 reg2146,
                 reg2145,
                 forvar2144,
                 reg2143,
                 reg2142,
                 forvar2141,
                 reg2140,
                 reg2139,
                 reg2138,
                 reg2137,
                 reg2136,
                 forvar2135,
                 forvar2134,
                 reg2133,
                 reg2132,
                 forvar2131,
                 reg2130,
                 reg2129,
                 reg2128,
                 reg2127,
                 reg2126,
                 reg2125,
                 reg2124,
                 reg2123,
                 reg2122,
                 reg2121,
                 reg2120,
                 reg2119,
                 forvar2118,
                 forvar2117,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar2117 = (1'h0); (forvar2117 < (1'h1)); forvar2117 = (forvar2117 + (1'h1)))
        begin
          for (forvar2118 = (1'h0); (forvar2118 < (1'h1)); forvar2118 = (forvar2118 + (1'h1)))
            begin
              reg2119 <= wire2115[(3'h6):(1'h1)];
              reg2120 <= "Yw";
              reg2121 = (8'hb0);
              reg2122 <= (forvar2117[(2'h3):(1'h0)] <= (-forvar2117[(4'ha):(4'h8)]));
              reg2123 <= (+"J6AuDu1n7aysTopLGZF48ei7b");
              if ($signed(($signed(reg2122[(1'h0):(1'h0)]) ?
                  (({reg2123, wire2116} ?
                      "Aa19fxfFQxM" : {forvar2117}) >> "m0zxHui") : reg2122[(4'h9):(3'h7)])))
                begin
                  reg2124 = "H";
                  reg2125 <= ((^~"ot") ?
                      (^~$signed(reg2121[(3'h7):(2'h2)])) : $signed("l93BQznVL"));
                  reg2126 <= (&(~(+forvar2117)));
                  reg2127 <= reg2122[(4'hb):(4'ha)];
                end
              else
                begin
                  reg2124 <= ({(((&reg2125) && (wire2114 ?
                          wire2114 : wire2114)) || (((7'h4d) ?
                              forvar2118 : forvar2118) ?
                          $unsigned(wire2115) : "4"))} >= (&"cqlACGmui4o4OfOvnohI"));
                  reg2125 <= forvar2117[(3'h6):(2'h2)];
                  reg2126 <= wire2114[(2'h2):(1'h0)];
                  reg2127 <= {wire2116,
                      (forvar2118 ?
                          reg2122[(2'h3):(2'h3)] : (+$unsigned(reg2126[(3'h5):(1'h0)])))};
                end
            end
        end
      reg2128 <= "QcZCfo4s";
      reg2129 <= "qaKLFk";
    end
  always
    @(posedge clk) begin
      reg2130 <= reg2122[(5'h10):(4'hf)];
      for (forvar2131 = (1'h0); (forvar2131 < (3'h4)); forvar2131 = (forvar2131 + (1'h1)))
        begin
          reg2132 <= ($unsigned({"vcrdXqdbMSDY8J"}) ?
              $signed($unsigned({reg2128})) : reg2126);
          reg2133 <= (8'ha6);
          for (forvar2134 = (1'h0); (forvar2134 < (3'h4)); forvar2134 = (forvar2134 + (1'h1)))
            begin
              for (forvar2135 = (1'h0); (forvar2135 < (1'h0)); forvar2135 = (forvar2135 + (1'h1)))
                begin
                  reg2136 <= (reg2124[(3'h4):(1'h1)] ?
                      ((($signed((8'ha1)) | "lORYVM") && {$unsigned((8'ha4)),
                              $unsigned(reg2125)}) ?
                          reg2123[(2'h3):(1'h0)] : ($signed(wire2113[(4'h8):(4'h8)]) ~^ $unsigned($unsigned((8'ha4))))) : "yGWIR7rCNlhwWPE7FPc6");
                  reg2137 = ($unsigned("YMd") <= $signed(reg2126));
                  reg2138 <= "uTr24OnJTF";
                end
              reg2139 <= reg2137[(3'h4):(3'h4)];
              reg2140 = reg2138;
            end
        end
      for (forvar2141 = (1'h0); (forvar2141 < (3'h4)); forvar2141 = (forvar2141 + (1'h1)))
        begin
          reg2142 <= $unsigned(($unsigned(({reg2124, reg2123} & (7'h4e))) ?
              reg2121[(1'h1):(1'h0)] : {("HqC" ?
                      $unsigned(reg2121) : (reg2122 ? reg2125 : reg2119))}));
        end
      reg2143 <= $unsigned($signed($signed("9FYrlf3PgH5pED")));
      for (forvar2144 = (1'h0); (forvar2144 < (3'h5)); forvar2144 = (forvar2144 + (1'h1)))
        begin
          reg2145 <= (~^(forvar2117[(4'hb):(4'h9)] ^~ reg2120[(1'h1):(1'h1)]));
          reg2146 <= forvar2131[(1'h0):(1'h0)];
          reg2147 = (8'ha8);
          reg2148 = forvar2117;
          reg2149 <= ($signed($unsigned(reg2124)) ?
              (($unsigned($unsigned(wire2113)) & reg2120) == (|reg2143[(4'h8):(2'h3)])) : (^(^reg2126)));
        end
      reg2150 = (((((reg2127 ? (8'hb8) : reg2126) ?
              reg2137 : reg2124) >> {(reg2145 <<< (8'ha0))}) ?
          forvar2144[(4'hf):(4'hb)] : {(7'h48)}) != (forvar2134[(3'h6):(2'h2)] ?
          $unsigned(reg2143) : ($signed((reg2143 & wire2115)) << (^$signed(forvar2117)))));
    end
  always
    @(posedge clk) begin
      reg2151 <= ({(forvar2141 <= $unsigned((-reg2149))),
              (&({(8'hbb)} != (-forvar2134)))} ?
          $unsigned((wire2115[(5'h11):(1'h0)] - (7'h46))) : (reg2136 ?
              ((^~(~reg2125)) ^ wire2116) : ("" < (reg2145 ~^ {forvar2135,
                  reg2143}))));
    end
  always
    @(posedge clk) begin
      reg2152 <= ($signed((~^reg2124[(2'h3):(2'h3)])) ?
          (+($unsigned(reg2124) & ($unsigned(reg2151) ?
              $unsigned(reg2129) : $signed(reg2150)))) : ($signed($unsigned($signed(wire2114))) >= $signed($unsigned((reg2126 ?
              (8'hbe) : (7'h47))))));
      reg2153 = reg2147[(1'h0):(1'h0)];
      reg2154 = $signed({"fs3k"});
    end
  assign wire2155 = $unsigned((^"0vfR1gX5Ve2Hbuxd8p"));
  always
    @(posedge clk) begin
      reg2156 <= forvar2118;
    end
  always
    @(posedge clk) begin
      reg2157 <= $signed($signed(reg2148[(4'h8):(1'h1)]));
      reg2158 = $unsigned((-{reg2125, $signed(reg2133)}));
      reg2159 <= $unsigned({{($signed(wire2115) || (reg2151 ?
                  reg2151 : (8'hbf)))},
          $unsigned(($unsigned(wire2116) && $unsigned(reg2140)))});
      reg2160 <= reg2146;
      reg2161 <= (8'hbb);
    end
  always
    @(posedge clk) begin
      reg2162 = (reg2129[(4'hd):(3'h5)] ? wire2155[(2'h3):(2'h3)] : reg2127);
      reg2163 <= (^~(+(^~reg2153[(5'h11):(5'h10)])));
      reg2164 = $signed(reg2129);
    end
  always
    @(posedge clk) begin
      reg2165 <= reg2137;
      reg2166 <= (reg2157[(3'h5):(2'h3)] >>> "7g");
      reg2167 <= reg2121;
      reg2168 <= (!"JMuToxNzVdTARPyeEvZ5k");
      reg2169 <= $signed(((^reg2157[(4'ha):(2'h2)]) ?
          (!(reg2138 ? wire2115 : (~^reg2156))) : (reg2151[(4'ha):(1'h0)] ?
              ({reg2160} << $unsigned((7'h4e))) : ("Z87BMnOoqfLqH9zDxPHs9J" ?
                  {forvar2118, reg2145} : $signed(reg2159)))));
      for (forvar2170 = (1'h0); (forvar2170 < (2'h2)); forvar2170 = (forvar2170 + (1'h1)))
        begin
          reg2171 <= ("JhGFSw" ?
              "s2NBnHaM35EYPFHp742f" : $signed((+$unsigned($unsigned(reg2160)))));
        end
    end
  assign wire2172 = (^reg2164[(2'h3):(2'h3)]);
  always
    @(posedge clk) begin
      reg2173 = reg2161;
      reg2174 <= forvar2118;
      reg2175 <= $signed(({((~&(8'hab)) ? wire2172[(4'h9):(3'h6)] : wire2114),
              (~^(reg2161 == (8'hbc)))} ?
          (({(8'hae)} ?
              $unsigned(reg2147) : (wire2155 <<< reg2120)) | (reg2140[(1'h1):(1'h0)] ?
              (reg2166 >> reg2121) : $unsigned(reg2124))) : reg2128));
      reg2176 <= "S1IFhC6zW90sp";
    end
  assign wire2177 = forvar2131[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg2178 = "5V";
      reg2179 <= reg2156;
    end
  always
    @(posedge clk) begin
      reg2180 <= "vioTuSr4DTfvSJZdF2XRnvAFO";
      reg2181 <= (("v1Gob8ZsRvIlFN7UeWJ" != (("m6DQNDWuwIbyfP8GTk" < "GIEUzUy5yKcoASRfGlMtkvkHT") <= ($unsigned(reg2137) ?
              (reg2152 ? reg2139 : reg2120) : $signed(reg2133)))) ?
          $signed({(reg2143 ? "X9lgrQD2ITy0" : $signed(reg2138)),
              $unsigned($unsigned(reg2129))}) : reg2142);
      reg2182 = $unsigned((^~"svKBg2i"));
      reg2183 <= reg2162;
      reg2184 <= (reg2180 ?
          reg2159[(3'h5):(3'h4)] : (|$signed($unsigned($unsigned(reg2142)))));
    end
  always
    @(posedge clk) begin
      for (forvar2185 = (1'h0); (forvar2185 < (1'h1)); forvar2185 = (forvar2185 + (1'h1)))
        begin
          reg2186 <= (^~$unsigned({$signed((reg2182 - reg2156))}));
          reg2187 = (|{{"eDSFAq6vgqa9BYLPt", {reg2122}},
              reg2175[(3'h6):(3'h4)]});
          reg2188 <= "ht3FYu7M";
          for (forvar2189 = (1'h0); (forvar2189 < (1'h0)); forvar2189 = (forvar2189 + (1'h1)))
            begin
              reg2190 <= $signed($signed((&reg2179[(2'h3):(1'h0)])));
            end
        end
      reg2191 <= (({($signed(forvar2185) ?
                      reg2120[(4'he):(4'hc)] : forvar2170[(2'h3):(1'h1)])} ?
              reg2147 : $signed((reg2182[(4'hc):(4'h8)] ?
                  (8'h9d) : (reg2156 ? reg2175 : reg2139)))) ?
          {reg2119[(3'h4):(1'h0)]} : "4cX");
      reg2192 <= (("tEMmIS3AzSAdW6Kbk" == forvar2117[(4'h8):(2'h2)]) ^ (reg2161[(4'hf):(3'h5)] <= reg2139[(3'h7):(3'h6)]));
    end
  always
    @(posedge clk) begin
      reg2193 <= ((!("7tU6Ptm2ez1MHgE15xG" || $unsigned("vqHET9z1FNqmYp"))) ?
          $signed($unsigned((((8'hb9) ^ reg2168) <<< (reg2162 ^~ reg2188)))) : reg2154[(4'hf):(3'h4)]);
    end
  assign wire2194 = ((~&$unsigned($signed("uIv5yo"))) ?
                        forvar2189 : (^(($unsigned(reg2184) ?
                                $unsigned(reg2156) : reg2164[(2'h3):(1'h1)]) ?
                            ($unsigned((7'h48)) >> $signed(reg2124)) : (&{(8'hb2),
                                reg2140}))));
  assign wire2195 = reg2174[(3'h5):(1'h1)];
  assign wire2196 = $unsigned($signed($unsigned((reg2167[(3'h6):(1'h1)] ?
                        "lVuAcSMSTzIK" : (8'hb8)))));
  always
    @(posedge clk) begin
      reg2197 <= reg2173;
      reg2198 <= (7'h4e);
    end
  always
    @(posedge clk) begin
      reg2199 = (reg2150[(3'h6):(2'h2)] != (^(({(7'h4a)} ?
          ((8'hbf) & (8'hb6)) : (^reg2138)) >>> "72cNDSLJR4yaSqNKQ9R")));
      reg2200 <= "rAq9RUgvhMsfzZepnO5ttCuQ2";
      reg2201 <= $unsigned(reg2171);
      reg2202 <= (8'haa);
      reg2203 <= "bnUPoLeTIqwYQ";
      reg2204 = ($unsigned((!$signed((reg2169 > reg2128)))) ?
          (reg2161 ?
              $signed($signed((reg2174 != wire2116))) : ("UkB8Runf" ?
                  reg2192 : (reg2183[(2'h2):(1'h1)] ^~ (forvar2117 > reg2130)))) : reg2202);
    end
  assign wire2205 = reg2162;
  assign wire2206 = $unsigned($unsigned(((8'hbf) >> (~reg2139))));
  assign wire2207 = $unsigned(("BvMa" ?
                        (reg2198[(1'h0):(1'h0)] >> (|{reg2171})) : (reg2201[(3'h4):(3'h4)] < $signed((reg2167 * wire2155)))));
  always
    @(posedge clk) begin
      reg2208 <= (reg2121[(1'h1):(1'h0)] >= (((-{reg2161, reg2149}) ?
          $unsigned((^~wire2207)) : reg2179) == "CECRfIuT4f5nb"));
      for (forvar2209 = (1'h0); (forvar2209 < (2'h3)); forvar2209 = (forvar2209 + (1'h1)))
        begin
          reg2210 <= {forvar2135[(4'h8):(3'h6)],
              ("7PgE" ?
                  {reg2180[(2'h2):(2'h2)],
                      $signed("5U19yzOmZvrh")} : $unsigned((((8'h9f) & reg2127) ?
                      (reg2181 ?
                          wire2172 : reg2123) : wire2207[(2'h2):(2'h2)])))};
          for (forvar2211 = (1'h0); (forvar2211 < (3'h5)); forvar2211 = (forvar2211 + (1'h1)))
            begin
              for (forvar2212 = (1'h0); (forvar2212 < (3'h4)); forvar2212 = (forvar2212 + (1'h1)))
                begin
                  reg2213 <= "Q2mSw";
                  reg2214 <= (($unsigned({reg2150[(4'h8):(3'h5)]}) >>> "hRHBU") ?
                      (!reg2192) : "20YhUMy5cdxWBtR6HyuDsHY");
                end
              reg2215 <= reg2164[(3'h4):(3'h4)];
            end
          reg2216 <= reg2192[(1'h0):(1'h0)];
          reg2217 <= (~&$unsigned($unsigned((reg2123[(1'h1):(1'h0)] ?
              $signed(reg2193) : reg2159[(4'hb):(4'h9)]))));
          reg2218 <= forvar2134;
        end
      for (forvar2219 = (1'h0); (forvar2219 < (1'h1)); forvar2219 = (forvar2219 + (1'h1)))
        begin
          for (forvar2220 = (1'h0); (forvar2220 < (3'h4)); forvar2220 = (forvar2220 + (1'h1)))
            begin
              reg2221 <= "YEJG5pnJYagwBghlOnRyGN";
            end
          reg2222 <= (-$unsigned(reg2130[(1'h1):(1'h1)]));
          reg2223 <= reg2129[(4'hc):(3'h4)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2028  (y, clk, wire2032, wire2031, wire2030, wire2029);
  output wire [(32'h3df):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire2032;
  input wire [(4'h9):(1'h0)] wire2031;
  input wire signed [(5'h15):(1'h0)] wire2030;
  input wire signed [(5'h15):(1'h0)] wire2029;
  reg [(4'h8):(1'h0)] reg2100 = (1'h0);
  reg [(5'h19):(1'h0)] reg2099 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2098 = (1'h0);
  reg [(4'h9):(1'h0)] reg2097 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2096 = (1'h0);
  reg [(5'h15):(1'h0)] reg2095 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2094 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2093 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2092 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2091 = (1'h0);
  reg [(2'h3):(1'h0)] reg2090 = (1'h0);
  reg [(5'h18):(1'h0)] reg2089 = (1'h0);
  reg [(5'h17):(1'h0)] reg2088 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2087 = (1'h0);
  reg [(4'hc):(1'h0)] reg2086 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2085 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2084 = (1'h0);
  reg [(5'h13):(1'h0)] reg2083 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg2082 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2081 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg2080 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2079 = (1'h0);
  reg [(5'h15):(1'h0)] reg2078 = (1'h0);
  reg [(3'h4):(1'h0)] reg2077 = (1'h0);
  reg [(4'hc):(1'h0)] reg2076 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2075 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar2074 = (1'h0);
  reg [(5'h11):(1'h0)] reg2073 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2072 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2071 = (1'h0);
  reg [(4'hc):(1'h0)] reg2070 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2069 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg2068 = (1'h0);
  reg [(5'h10):(1'h0)] reg2067 = (1'h0);
  reg [(5'h13):(1'h0)] reg2066 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2065 = (1'h0);
  reg [(5'h11):(1'h0)] reg2064 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar2063 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2062 = (1'h0);
  reg [(3'h5):(1'h0)] reg2061 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2060 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg2059 = (1'h0);
  reg [(4'hc):(1'h0)] reg2058 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2057 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2056 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2055 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2054 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2053 = (1'h0);
  reg [(4'he):(1'h0)] reg2052 = (1'h0);
  reg [(5'h11):(1'h0)] reg2051 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2050 = (1'h0);
  reg [(5'h12):(1'h0)] reg2049 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg2048 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2047 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2046 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg2045 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2044 = (1'h0);
  reg [(5'h16):(1'h0)] reg2043 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg2042 = (1'h0);
  reg [(3'h5):(1'h0)] reg2041 = (1'h0);
  reg [(5'h10):(1'h0)] reg2040 = (1'h0);
  reg [(5'h14):(1'h0)] reg2039 = (1'h0);
  reg [(5'h19):(1'h0)] reg2038 = (1'h0);
  reg [(5'h12):(1'h0)] reg2037 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2036 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2035 = (1'h0);
  reg [(5'h18):(1'h0)] forvar2034 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire2033;
  assign y = {reg2100,
                 reg2099,
                 reg2098,
                 reg2097,
                 reg2096,
                 reg2095,
                 reg2094,
                 reg2093,
                 reg2092,
                 reg2091,
                 reg2090,
                 reg2089,
                 reg2088,
                 forvar2087,
                 reg2086,
                 reg2085,
                 reg2084,
                 reg2083,
                 reg2082,
                 reg2081,
                 reg2080,
                 forvar2079,
                 reg2078,
                 reg2077,
                 reg2076,
                 forvar2075,
                 forvar2074,
                 reg2073,
                 forvar2072,
                 reg2071,
                 reg2070,
                 forvar2069,
                 reg2068,
                 reg2067,
                 reg2066,
                 reg2065,
                 reg2064,
                 forvar2063,
                 reg2062,
                 reg2061,
                 reg2060,
                 reg2059,
                 reg2058,
                 reg2057,
                 reg2056,
                 reg2055,
                 forvar2054,
                 reg2053,
                 reg2052,
                 reg2051,
                 forvar2050,
                 reg2049,
                 reg2048,
                 reg2047,
                 reg2046,
                 reg2045,
                 reg2044,
                 reg2043,
                 reg2042,
                 reg2041,
                 reg2040,
                 reg2039,
                 reg2038,
                 reg2037,
                 reg2036,
                 reg2035,
                 forvar2034,
                 wire2033,
                 (1'h0)};
  assign wire2033 = wire2030[(3'h5):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar2034 = (1'h0); (forvar2034 < (3'h4)); forvar2034 = (forvar2034 + (1'h1)))
        begin
          reg2035 <= wire2030;
          reg2036 <= (~|"w6mpqhc1zCtMShMbK80T8");
          reg2037 <= "FkALoRHnZw4";
          reg2038 <= $unsigned($signed(($unsigned("uyC7TDQe5BTumaWROkf3fT") ?
              ($signed((8'hb9)) ?
                  (7'h47) : (wire2033 ?
                      wire2033 : wire2032)) : (+reg2035[(1'h1):(1'h1)]))));
          reg2039 <= "";
          reg2040 <= ($unsigned("d") ?
              {(!(~^$unsigned(reg2036))),
                  reg2037} : (((&wire2029[(3'h7):(1'h1)]) ?
                      {(-reg2036),
                          (wire2029 < (7'h4e))} : (!reg2039[(1'h0):(1'h0)])) ?
                  "L5VETRpYeP2toREddY9Ols" : wire2030));
        end
      reg2041 <= (7'h45);
      reg2042 <= "6KdSA0KmF4x1M97UxE";
    end
  always
    @(posedge clk) begin
      reg2043 = "k6P8Usd6L3qMIpd9qF";
      reg2044 <= $unsigned(reg2041[(3'h4):(1'h0)]);
      reg2045 <= reg2039[(1'h1):(1'h0)];
      reg2046 = reg2038;
      reg2047 = ($unsigned((~|((reg2046 - wire2029) ?
          $unsigned(wire2033) : "O7biGKAUq"))) && $unsigned((($unsigned(wire2031) ?
          (|reg2046) : ((8'hb3) ? (8'hbe) : reg2043)) < (8'had))));
      reg2048 = {"rqt2L4C5zZMkTGzY2kAoR"};
    end
  always
    @(posedge clk) begin
      reg2049 <= $unsigned((wire2032[(2'h3):(1'h0)] >> reg2045[(3'h7):(3'h4)]));
      for (forvar2050 = (1'h0); (forvar2050 < (1'h0)); forvar2050 = (forvar2050 + (1'h1)))
        begin
          reg2051 = $unsigned({(|reg2035),
              $signed($signed((wire2029 ? reg2036 : wire2030)))});
          reg2052 <= wire2030[(4'hc):(2'h2)];
          reg2053 <= reg2042;
          for (forvar2054 = (1'h0); (forvar2054 < (3'h5)); forvar2054 = (forvar2054 + (1'h1)))
            begin
              reg2055 = reg2041[(2'h2):(2'h2)];
              reg2056 = reg2046;
              if (reg2039[(5'h10):(1'h0)])
                begin
                  reg2057 <= $unsigned(((&{forvar2050, (reg2046 ~^ wire2029)}) ?
                      (~^"4mJlu6N") : (&(|"70NQhaOuICIOUiH"))));
                  reg2058 <= $unsigned(wire2030);
                  reg2059 <= (^($unsigned("3Z7qEvKc9vEBJ6pSCf") * ((|reg2052[(1'h1):(1'h0)]) ?
                      (7'h48) : reg2052)));
                  reg2060 <= reg2053[(3'h5):(3'h4)];
                end
              else
                begin
                  reg2057 = ($unsigned("YAMb68l2") ?
                      ($signed((-reg2041[(3'h5):(3'h4)])) >= ($signed($unsigned(forvar2050)) ?
                          $unsigned("90dsU6Gbo1") : ("q6ItpoNQP" ?
                              (~|reg2044) : (wire2030 ?
                                  reg2038 : (8'h9e))))) : ($signed(reg2051[(3'h4):(1'h1)]) ?
                          reg2056 : (|reg2056)));
                  reg2058 = $signed(forvar2050[(3'h6):(1'h0)]);
                  reg2059 = reg2051;
                  reg2060 <= ($unsigned($signed((~|{reg2059,
                      forvar2050}))) >>> $unsigned($signed(((&reg2042) == (&reg2038)))));
                  reg2061 <= (!(&forvar2050[(1'h0):(1'h0)]));
                end
              reg2062 <= (~(+reg2056));
              for (forvar2063 = (1'h0); (forvar2063 < (2'h3)); forvar2063 = (forvar2063 + (1'h1)))
                begin
                  reg2064 = $unsigned((8'ha5));
                  reg2065 <= wire2031;
                  reg2066 = ((|(!(((8'ha7) << (8'hb4)) ?
                          reg2060[(3'h6):(2'h3)] : (reg2049 ?
                              (8'ha2) : (7'h4d))))) ?
                      $unsigned(reg2045) : ((($unsigned(reg2065) >> (&wire2030)) ?
                          "PJPG" : ((&reg2056) - wire2030)) >> $signed($unsigned($signed(wire2030)))));
                  reg2067 <= (^~((("5s5hTuTnymxgI1rYvCBdpG" ~^ ((7'h47) | wire2032)) ?
                          reg2058 : ($signed(reg2039) ?
                              $unsigned((7'h4a)) : (+reg2040))) ?
                      "sLWTA" : $signed($signed("6ZFmHwdGXpNLWcOqISrAL"))));
                end
              reg2068 = {reg2055};
            end
          for (forvar2069 = (1'h0); (forvar2069 < (2'h3)); forvar2069 = (forvar2069 + (1'h1)))
            begin
              reg2070 = reg2052;
            end
        end
      reg2071 = reg2060;
      for (forvar2072 = (1'h0); (forvar2072 < (1'h0)); forvar2072 = (forvar2072 + (1'h1)))
        begin
          reg2073 <= ("39lVD" ?
              (~^(~&$signed($unsigned(wire2033)))) : reg2066[(4'h9):(2'h3)]);
          for (forvar2074 = (1'h0); (forvar2074 < (1'h0)); forvar2074 = (forvar2074 + (1'h1)))
            begin
              for (forvar2075 = (1'h0); (forvar2075 < (1'h1)); forvar2075 = (forvar2075 + (1'h1)))
                begin
                  reg2076 = (!$signed({(reg2068 | forvar2069[(1'h0):(1'h0)])}));
                  reg2077 <= (~^{reg2055});
                end
              reg2078 <= (forvar2069[(1'h0):(1'h0)] ?
                  $signed(((!$unsigned((8'had))) ?
                      (reg2040 ?
                          {reg2067, reg2077} : (reg2055 ?
                              (8'ha5) : reg2070)) : reg2037)) : (($unsigned((&wire2032)) == reg2036) == ((~^$unsigned((8'ha0))) > $signed((reg2070 * reg2053)))));
              for (forvar2079 = (1'h0); (forvar2079 < (3'h4)); forvar2079 = (forvar2079 + (1'h1)))
                begin
                  reg2080 <= forvar2069;
                  reg2081 <= (8'hb6);
                  reg2082 = "cKR";
                  reg2083 <= (~"StlSUVQh1NQy9oIygp");
                  reg2084 <= $signed($signed((-$signed($unsigned(reg2041)))));
                end
              reg2085 <= $signed((-reg2053[(3'h4):(2'h2)]));
              reg2086 = wire2030;
              for (forvar2087 = (1'h0); (forvar2087 < (1'h0)); forvar2087 = (forvar2087 + (1'h1)))
                begin
                  reg2088 <= $signed("P0foUpiG7TAFEbPN4Gw7");
                  reg2089 <= reg2066[(2'h3):(1'h0)];
                  reg2090 <= {(($unsigned($unsigned((8'hb2))) ?
                          $signed(reg2056) : {(^~forvar2034),
                              $unsigned((7'h47))}) * ((!reg2070) ?
                          reg2084 : $signed($signed(forvar2072)))),
                      wire2033};
                  reg2091 = forvar2069[(2'h2):(1'h0)];
                  reg2092 <= ($signed(forvar2087[(1'h0):(1'h0)]) ^~ ($signed("XD0DbsgW") ?
                      "pHmiTym9EVlKU" : (reg2085 == {$signed(forvar2054)})));
                  reg2093 = $unsigned(("" ?
                      (|{"nma4d63", "8uBSYWEeSFU8PeoAhVG"}) : $signed("4R")));
                end
            end
        end
      reg2094 <= (~|(~&reg2071[(3'h5):(3'h5)]));
      reg2095 <= (~|(^$unsigned($unsigned(reg2051))));
    end
  always
    @(posedge clk) begin
      reg2096 <= {reg2085[(1'h1):(1'h1)]};
    end
  always
    @(posedge clk) begin
      reg2097 <= $signed((~^(!(((7'h49) + reg2095) ?
          $unsigned((8'ha2)) : $unsigned(reg2056)))));
      reg2098 <= reg2091[(4'h8):(3'h7)];
      reg2099 = {($unsigned("kk4GF5YVbJCb3EB8sBT") ?
              $unsigned((reg2091 ^~ (~|(8'ha7)))) : $signed(($signed(forvar2075) ^~ reg2060[(3'h5):(3'h5)]))),
          (8'had)};
      reg2100 <= {$unsigned($unsigned(reg2089[(5'h15):(1'h1)]))};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1953
#( parameter param2005 = ((((|((8'hb4) ? (7'h49) : (8'hb5))) ? (((7'h4d) ? (8'hac) : (8'ha1)) == (~^(8'ha5))) : ((8'hab) ? ((8'hb9) ? (8'ha7) : (8'ha9)) : {(8'hb6), (8'h9d)})) ? (~|(+((7'h4b) && (8'hae)))) : (({(8'ha9)} > ((8'hae) ? (8'hac) : (8'ha3))) ? {((8'ha0) ? (7'h48) : (7'h41))} : {(~^(7'h4b))})) ? ((({(8'hb4), (8'hb1)} ^ {(8'hbe)}) | ((~(8'hb7)) ? ((7'h4d) ? (7'h4c) : (8'hbe)) : (+(8'ha7)))) ? ((((7'h46) >>> (8'h9d)) && (|(7'h42))) ? ({(8'ha6)} ~^ (|(8'ha4))) : {(^~(8'ha6)), ((8'hbf) ? (8'hbf) : (7'h4a))}) : ((&{(7'h47), (8'h9f)}) <<< ((8'hbe) ? ((8'h9c) << (8'ha6)) : ((7'h45) << (8'hb2))))) : ((({(7'h4a)} ? ((8'h9f) ^~ (7'h43)) : ((8'hb0) ? (7'h49) : (7'h43))) ? ({(7'h40), (8'hbb)} >> ((8'hbd) ? (8'hb0) : (8'haf))) : (((8'h9f) != (7'h43)) ? ((7'h48) ? (7'h44) : (8'hbb)) : ((8'hab) ? (8'ha6) : (7'h49)))) >> ((~{(7'h48)}) ? (((8'hbe) >> (8'hb0)) ? ((7'h49) > (8'hb6)) : {(8'h9c), (8'hbe)}) : (((8'haa) ? (8'hb2) : (8'hb0)) ? ((7'h41) ? (8'h9e) : (8'hae)) : ((7'h43) <= (8'hbc)))))) )
(y, clk, wire1958, wire1957, wire1956, wire1955, wire1954);
  output wire [(32'h26f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire1958;
  input wire signed [(4'hc):(1'h0)] wire1957;
  input wire [(5'h12):(1'h0)] wire1956;
  input wire [(5'h15):(1'h0)] wire1955;
  input wire [(3'h7):(1'h0)] wire1954;
  wire [(5'h14):(1'h0)] wire2004;
  reg signed [(4'hf):(1'h0)] reg2003 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2002 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg2001 = (1'h0);
  reg [(4'h9):(1'h0)] reg2000 = (1'h0);
  reg [(4'he):(1'h0)] reg1999 = (1'h0);
  reg [(4'hd):(1'h0)] reg1998 = (1'h0);
  reg [(5'h18):(1'h0)] reg1997 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1996 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1995 = (1'h0);
  reg [(3'h4):(1'h0)] reg1994 = (1'h0);
  reg [(4'hd):(1'h0)] reg1993 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1992 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1991 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1990 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1989 = (1'h0);
  reg [(5'h19):(1'h0)] reg1988 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1986 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1987 = (1'h0);
  reg [(3'h6):(1'h0)] reg1986 = (1'h0);
  reg [(4'hf):(1'h0)] reg1985 = (1'h0);
  reg [(4'hb):(1'h0)] reg1984 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1983 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1982 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire1981;
  reg [(5'h14):(1'h0)] reg1980 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1979 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1978 = (1'h0);
  reg [(3'h5):(1'h0)] reg1977 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1976 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1975 = (1'h0);
  reg [(5'h11):(1'h0)] reg1974 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1973 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1972 = (1'h0);
  reg [(5'h11):(1'h0)] reg1971 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1970 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire1969;
  reg signed [(5'h14):(1'h0)] reg1968 = (1'h0);
  reg [(5'h19):(1'h0)] reg1967 = (1'h0);
  reg [(3'h7):(1'h0)] reg1966 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1965 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1964 = (1'h0);
  reg [(4'hd):(1'h0)] reg1963 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1962 = (1'h0);
  reg [(4'h8):(1'h0)] reg1961 = (1'h0);
  reg [(5'h12):(1'h0)] reg1960 = (1'h0);
  reg [(5'h12):(1'h0)] reg1959 = (1'h0);
  assign y = {wire2004,
                 reg2003,
                 reg2002,
                 reg2001,
                 reg2000,
                 reg1999,
                 reg1998,
                 reg1997,
                 reg1996,
                 reg1995,
                 reg1994,
                 reg1993,
                 forvar1992,
                 reg1991,
                 reg1990,
                 forvar1989,
                 reg1988,
                 forvar1986,
                 reg1987,
                 reg1986,
                 reg1985,
                 reg1984,
                 forvar1983,
                 reg1982,
                 wire1981,
                 reg1980,
                 reg1979,
                 reg1978,
                 reg1977,
                 forvar1976,
                 reg1975,
                 reg1974,
                 reg1973,
                 reg1972,
                 reg1971,
                 reg1970,
                 wire1969,
                 reg1968,
                 reg1967,
                 reg1966,
                 reg1965,
                 forvar1964,
                 reg1963,
                 forvar1962,
                 reg1961,
                 reg1960,
                 reg1959,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1959 <= wire1958[(2'h2):(2'h2)];
      reg1960 <= "1f1r71nJJRx8WooKIKB";
      reg1961 <= ((^~"Oz07aq8K5uHzG1Xv") ?
          ($signed($unsigned("ADOxqdaxB")) ?
              (((reg1959 ? (7'h40) : wire1955) ?
                  "Z5id9X" : (wire1954 ?
                      (8'h9e) : wire1957)) || {"lcGeE4YY5R61o0QSvIkMQ",
                  (wire1957 ?
                      wire1957 : wire1954)}) : wire1956) : ((~&$signed(((8'ha7) ?
                  wire1958 : wire1955))) ?
              {(^~"BorsXpno3BflBxvNOZzv8"), reg1959} : (!(^~(8'hbd)))));
      for (forvar1962 = (1'h0); (forvar1962 < (1'h0)); forvar1962 = (forvar1962 + (1'h1)))
        begin
          reg1963 <= wire1958[(2'h3):(2'h2)];
          for (forvar1964 = (1'h0); (forvar1964 < (2'h2)); forvar1964 = (forvar1964 + (1'h1)))
            begin
              reg1965 <= ({"ShGXX9TrO", wire1958} ?
                  "2QCPcSRQa3fGEVaG" : (forvar1964[(1'h1):(1'h1)] ~^ (((|(8'hbe)) | ((7'h49) ?
                      (8'ha8) : wire1957)) <= $unsigned((forvar1964 > (7'h4d))))));
              reg1966 <= reg1963[(4'h8):(3'h5)];
              reg1967 <= reg1960[(4'hf):(4'hb)];
            end
        end
      reg1968 <= $unsigned((wire1958[(3'h6):(3'h5)] ^~ forvar1962[(1'h0):(1'h0)]));
    end
  assign wire1969 = (8'h9c);
  always
    @(posedge clk) begin
      reg1970 <= $unsigned((~|wire1957[(3'h6):(3'h5)]));
      reg1971 = (~^$unsigned(($signed((reg1968 ? reg1959 : reg1967)) ?
          reg1968[(4'hb):(4'h9)] : reg1960[(4'he):(4'he)])));
      reg1972 <= (7'h40);
      reg1973 <= (|$unsigned($signed(wire1954[(1'h0):(1'h0)])));
      reg1974 <= $unsigned((|(($signed(wire1958) ^~ (reg1968 ?
          (8'hb7) : wire1955)) <= forvar1964[(1'h0):(1'h0)])));
    end
  always
    @(posedge clk) begin
      reg1975 <= ($signed({(wire1954[(2'h2):(2'h2)] == $signed(wire1955))}) && reg1971);
      for (forvar1976 = (1'h0); (forvar1976 < (2'h2)); forvar1976 = (forvar1976 + (1'h1)))
        begin
          reg1977 <= (!reg1973[(2'h3):(1'h0)]);
          reg1978 = "g8vA2sXet8WtIUFObKCuF";
          reg1979 = "dWm1de7BYUJQZXnRwQW";
        end
      reg1980 <= (~^$signed($signed({reg1970[(2'h2):(1'h1)]})));
    end
  assign wire1981 = $signed($unsigned(reg1967[(5'h10):(4'hb)]));
  always
    @(posedge clk) begin
      reg1982 <= $signed(reg1977);
      for (forvar1983 = (1'h0); (forvar1983 < (3'h4)); forvar1983 = (forvar1983 + (1'h1)))
        begin
          reg1984 <= wire1969[(2'h3):(2'h3)];
          if (((~&(~^(&(8'ha5)))) + $signed("axKwCyaswbrspkks")))
            begin
              reg1985 <= reg1978;
              reg1986 <= (~^reg1965[(3'h4):(1'h1)]);
              reg1987 <= "B129NEW009";
            end
          else
            begin
              reg1985 <= (~&reg1987[(1'h0):(1'h0)]);
              for (forvar1986 = (1'h0); (forvar1986 < (3'h5)); forvar1986 = (forvar1986 + (1'h1)))
                begin
                  reg1987 <= "V3";
                end
              reg1988 <= (($signed($signed(((8'haf) ^ reg1978))) ?
                  $signed((8'hbd)) : ((reg1966[(3'h4):(2'h2)] ?
                      {reg1966} : reg1970) && ({reg1966,
                      reg1963} && reg1961[(1'h1):(1'h1)]))) == (reg1974[(3'h5):(2'h3)] >>> ((-((7'h48) ?
                      wire1954 : wire1969)) ?
                  (+"2qANQih") : (~|"dx2m"))));
            end
          for (forvar1989 = (1'h0); (forvar1989 < (1'h0)); forvar1989 = (forvar1989 + (1'h1)))
            begin
              reg1990 <= reg1968[(5'h11):(4'hd)];
              reg1991 = (($signed((~|"ACbFX")) ?
                      forvar1983[(5'h15):(5'h11)] : (reg1984 & ($unsigned(forvar1976) == (reg1974 ?
                          reg1972 : reg1987)))) ?
                  "QoqD61Xio" : forvar1976);
              for (forvar1992 = (1'h0); (forvar1992 < (2'h3)); forvar1992 = (forvar1992 + (1'h1)))
                begin
                  reg1993 <= (^~reg1973[(2'h2):(2'h2)]);
                  reg1994 <= ({reg1965[(3'h4):(1'h1)]} | $unsigned((-"vH1tiKJFTpcpRU4qx")));
                  reg1995 <= (~reg1979);
                  reg1996 <= (wire1954[(2'h2):(2'h2)] << ($unsigned((wire1956 + (+forvar1992))) <= wire1958[(3'h5):(3'h5)]));
                  reg1997 = ("Hi6oce5V56tvKCR" > (($signed(reg1984[(4'hb):(1'h1)]) ?
                      $signed($unsigned((8'hbc))) : "UK0Seu") > forvar1976[(3'h7):(3'h4)]));
                  reg1998 <= reg1994;
                end
              reg1999 = $signed((~$signed(($unsigned(reg1975) * "tdXlkn"))));
              reg2000 <= forvar1964;
            end
          reg2001 <= $unsigned((7'h42));
        end
      reg2002 <= (^~({$unsigned((reg1970 ? reg1978 : reg1966))} ?
          (!(&$unsigned(reg1967))) : "OGmYgqhPhtFXW"));
      reg2003 <= "KZqWnEbiGx9eXYY61eYv";
    end
  assign wire2004 = {wire1954[(2'h3):(2'h2)], reg1975};
endmodule